`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17840)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCahs3fiyq/876fXZqyDwf+7PkhJpVv6VH4oTQGygL5Uv//sG6xEAcS9t
kDo+KloLrOgMhNR5L3CYwsHxaG9AbH4njT9wgB/3JQQEg6s7PIYDE3gBV9yk0uw7lfHn3lwq5YK3
I4Y/71qYBDAOKBaRZmulmJ7U7b7awKHQ15gdRWNLEI79CKizmbTKGlw846blXnqUKAviCDkRaB+I
NGpfpmKALav6iIc4hFA6re7Ob3MGTFhfFLEMpdPROfh3oyLv4yXwyLIRrpIygkUjK7knGEnuw/W6
Wr56V7o0/Kzl0Uwpxcf6T1maEjXAmah0KsBSl0t2qJOVNyivkqBYVjhRXPwLzSvwiqZPvwQGyLdE
Sd0WeftpzzaTHLvvWEL8gnnojw5I92kBdZjes58cIgrFRV7KBbOD7gzMX2sAHGiUGhIQywD/lz6S
U2Ppr20b7JgGrJe+U/+OwpZ+mSAuZDJozFZFHmCjOUrslYTdEgfQ5vtaTussENvoyqI+2CyYXPYx
cDuUl+ExTWte/GRSM1+yILuC2Aba+sxfEApYQa3fsf0lzftOJ38KK3UFnztW/VEAYsfqBpHworUb
uTnRGQs6FZRfjWgwZxENpRnOD2V7MQN4xIMF30R2Z0cSlImrm3ZMfNJCTgCglHQwG/OBmfmfMmOU
yXSH5yoHydNszITANIjRCqfjNnos7NMB22EhxhYX3UgK2wVHOg/Tl/8Ga06JLjYi8xGEyg32i3C4
TIGaIhPoxryD+8vNaVmDRMdS4m6qZAYf9imfeLWfmNPKp89Lq3u8qy/A0/sFSZbA7WUUkzhTRts9
UZ0LiRtNqpt9BkdayRdJbQknEiyo88URCPeGA0IO/mx7OtrKjcfDvfRvZxG0CmpWfNtJ+DO9f7Lb
Lt6U8y6qpkhfBSor7z1vCXwKlespRSdnJ+0Htk5ExBri2Gx1uIPtS/EHR1Sqy6lyPH8zVT0ip/yE
DlKuCMz3dBoPOQhhTfTZxXKUdsJ+yBKDIDMBtDUEDcDGGAm7VdbQsM+6pDZJw603vTyStCVmdiIx
cbeB3Eh/tD3WlTyuxBg3I/uo4eM+CeqqHTe/Ewq/Bi6w02xPz/wWcuyHL/a3GloQ/+gzJLoIygp+
mYAt/j6AVDa3Q1FHX6eftVJNYs1AHwoQuWypy7ApQGWWk1iui3kFO44Y2DZbNrQzbIILPxMZbvMN
9t4bFJ1jZa6xatUEooHmItmLHbOSIwDryjAPCOJv6q/lw5FXTiyhVhq7phAlBVd95PITyvStK13z
pc9oyeYqxrnRy95IFqwkl8smbtOpkpieEs5Zuk6FzXn6P+K0sg7kgSuy4Qxm4XXvJGL+KZLOtOu+
jii8WlikKmJR4vOs4+QI52O6nMWgP3ZG/NlPB3SNS0zy82rlCP+5jimWn+K1yvt3Y5uV522SCr9v
S5HClj2o0a+PcstH0n+B/78BykQ594O1aUMC6yZahLk3v8l7GwL3e39KjL8HCm59AMoWvVy5qJAk
/KEsqUf4UHY5rq++GXnKGYqulWM84YwrOva14aPZg/XkWx0Q5lKpg8RtIr5W0hFIVlsklwGnKiXB
Xfz1chp97lc4vGm+jys/26sb2S/YtwxdW1jhmSO5/ZHuBJIyBumi14EiFeG6kVt1nbKkqB+TXXlT
TK0SPwSMRsQI7oCpexw/Ruokza5ItUDLgoYqpNhpmnieJM2TIuRfjc9pKA0ipGguqwT1GbEvjXBR
SDw9IJd0CaPWH89jJwAnRNuPAlCdxyEs8Bia1OGWL25euSjiVmWVhayM39hl84JyxCmOYXQvSZpw
HMXI9kuI5KXh6FO96sHUJ4Z6ktCIwmuhzVF8zCIolisKeVEEjHyZSQVkn/upxXur0spegFsaC3+m
o8MhoCaO7iu7Ey9W4+VfzLJ6C4r1y0t8PuO10ciScVA5R1iBOFmXLGcVQZbYPtZGXaQlLgnfyHS2
KZVN3vQhJqGesIgmlbJ/P/OauZhrCK4+qSdz54Yt/t2HAhMD8kYv3o7rbMsMCve7PW/iADcsGT+K
xujYMFujT6VFn5JmjUMMk3azhgFuNSaYv99ZjucJ2B0+pKF4cspQXzV85qKQlHJfqjd0M/ps6RZC
/UjkW6eaN44j1RuqRwejDYierNQJ+N33g3NXuRVdesKiopdgW14qR5VEUUfRR3g2ejFNFZeVR4Yd
ErgCJDrjOkOhRFqd8M4BVzLokupnxic3lgQDgAuyuvpM5R9UdrDmUoOBga8uJP1qkxUFdungvsj1
o8QiFvfZ4OSjW6/X4T6VHUbc6hjb6k118I2hHRmu77moApzbnAa0gkMo/kflitsTfGZnJ0KvGgkW
nG3HSPa4Rk/dX4Z0Zj8TUjB+VqhIB0HhNHggZTBNbK8RAwk2oX+cVmg2HrwvyUnD9caTENXf+zwt
IRR0xZ05Jmc3WTNz5FOOzQU73cAc6jiQrdsL293N/5Kd27Inb2dc12adDYP3Rrt9T9O9GGhqXmbN
Aoy4/tuOdWdVXnHF0DtLJKn+z5p3BgB/QPPjK/kgZFfMeJPugijU33zM0xPODihvasr9eoaFT6Y+
AIyfwfC+rqvrlTmDnbtwbz9iNfk5mD4wVfNOU8GxbwXUtp13/13xIBo8UMJsDMFOGTGciuywH3wc
jaosu8ZKupsqwEwPP4LWzwKBQsrNlS0J7nNIv0msJhyScEuwtXc+utLUZlo+9GO3wRLZIuKQ8dH+
NtNSYswSbld1f6Jp8s1Wb7Pw3loEexgn528gY1Ws6cWPMghk4y8qQfuj88wItr0MsVB5U801ibPm
R88ZsnHA8vQycxIgWrYyxrhNpsGHpW7NaedQSVBc7MgWNGlwKRU8jsOZu95wYl31oSfGYew1HScs
NJld/PeVUeKcba4serKQRHa5NXCCN9dGJD74dx4zjQCc5xTz+jF3oCaNtFtCMHbkoumts506cG/o
Z/Z6fUV0NLmAV9JN7mQi8J1injVTDZ7wzjH22EYtFkM+vEy7gCCDk8nwZsBZikuPcKy55YNT3jet
pzRHeB36yM83VGHTDfJftExsrm+VXGFAn8mDZ2DHWPQ9cikApsvfvU78MYdMt9X9WYFMTA5c7O2S
D8iLhdvWtCurOzJmsRqzmcB/FJBVjBhKXgXZ5yRwyuS1SOJT0PlB8Pk1btYEVx7B1Q09aj9+1jbZ
8txVF6oWpSiiP0sCY14ItjFKVKgi4tooLk+Y1dOu4GrcLWh7Zf4HbMklluELlQfIMRaaH48EsgKl
rRFd/e3efUtodewfsCnkdU6lTONRYLFS3VJlxVW9HQtU4FJ5aIRs0J6FIqFUXqKvb+qrlthUD+qt
IysjLH1K9YCQkN421i3/MGW818JPa3vsP5ZsD10+8LvxDJojDDsTO7t4JQ3cTLC5fS88T6Ur5tRX
cK/mF3dJULxtAc0y1MEFeXnKo9uFU6lwENT5TcCiUbF45kWnNNnJV99IHhE6zK6sbmWajsnig86N
k2RFwt8B3/KlPzt2Dz0lxfK297hZHXb1yjc31kuPat93U8x6Vh7r4NAYJhdTTgeKX1alHQZagaKC
SU6OzoMJ1GaPSdSPJ+3MhvoMeLrn4HYnA2RYbG4G+eoGHWE8mUWBbCntT+lWHRMaUAqxvLEFeMof
uKOJh63ukbN4i3cY4kHM5ImLe/+wRXDvKjQFCbQbEg9Mw3LMr6dbXskqhB2ayG7vXp9UK6E6XlyL
FAf/3WJce+0t+hpAH5JbIpUz3B7rAQ5gQRfUrETtLIoaTPqQg5aY0QNW2DFtCkIorbUKVhsRo4Yb
cKTe4EKB+Q/qjeVLSJYUh6N6/Ymhoqqd2EPHIhINi3lwRXruT902YjRmfOlbpfM27XfvDSncs7Cv
9YQ926mbdNLxmGz0bXWzvb+mQVyohPMF+10B0CVoZXpTdAx3io3pPkRiRr95xanqJRO6+5l6yUjT
quofSeQ+2EOXlp8VvNvedMHG4uAQs/mBzXkyynp2G6SF2XxKCY2s/fxbjO1I+Jtu7qeMjuLNzIYR
6ygblF3mBNy8E31moV1Ua6K+noeMnx79ba5kQIWpjkWwtO5Ec7MhBvNoCsKiZwiuv5GiGFt2Vgk6
sF40LGWcoDPvYTyOtDBVoJV+3toRDZHbiYM+Qnm83IdZYvubMaXgB2KFyQMqA+n14QYgTAKSamb/
s8mT8OEadKPYSRrVC+evNDCzqJvBy4LAJguf+A5UWCflMbMkT3rPdLv9dXpBgWVr1I6s8etHVm5o
Vj2rJeJQF7zfrvdyk9ImyqA4VjdvX+wSW50ztrYn34xr2Xm6IeirVGIVExqyLD1tiVrTWtum4KR/
y6Zs0fnXYtZ+gpJT9YEHc8GEgcNOlXP83F35+USFjX2HQMDQvsOSLxNtKlTZtdRPQvFLU/IthRRW
dsSo41J8nGd9TUuvrlCFDaomh748hix7wqGAwiR/4MHI1e9F0rvoOlhGHM8r93rxLgAl8eewYGIR
fgdsWFW7S+L2ddPl3DppCYwhVpstFfuhaiab2ip4LI9vVonFw15XYNZx7PvZx3UQOg4zc7Z2uj2Y
id/PvpHEhGE+BHKwIw/X4zro2dbLk/9XtZpjNefRaeLpKglbPpFKLdpgwcNFtBfqlfTT0ZVpAwRj
zyGxN0spmN/qNkOzNrT4Fthr9LhXxiVOOGrpWZ7xKPeyYNPhQFh93DMouj32aL2XsWnCAj3AvYXk
1AtD+OFFbDVUnA+rwtaGtrZ0EpAz0liS8SmmJ9AmBYwGrwNB2G7uHj+h6OjCNsNhfA9pbaDbvFoQ
cfvsrId4SOA6Ki7GxhGOTCDJVzp0CJtfXAbLY4aI9NBYiZBbEfAzppVWL9y0ecqg/qAj9ifGJcVZ
mhH8LlgTlnJUF8bFy4y8DlSbfJRNsc65giydaTPBxD/BwRz//06uujgLT314V2Y59Tt8pguipHnN
EN1osyA32u7CN+fBE/TXGsX2D3uHgskSgAVOxYHnNQ9a3jTzKc9rOPiYO0TS32lcaGkvLJjCLDAu
c6qnnEW4Ysnn2Z3ZNhDVseU0JpXkyDRDynRdGBtu2qmTGRYro+2idAqiKoz95bOE/INg9XbdA18C
Aww5OggVmGONj8uYrTk2Fd7KyuseU4kue27aNo9P8I6nWGyD7fZHqCp7uwaWqhwCWnGvw91GIkxg
rMXSJaiySruPqzxcYry7aeZnLVmuXEnsju6KDmILPHnP4fJ/bUnXCdN9rYGP+RusemFgN+uX4i37
1kWIPLFIgEjHyzdtAZMEQBo1cdoiVYc5v44j/8UxZzuw/TILjwx2HFqt7wJvrwOmiFPjGEZRM4WF
QTx17q6ww9AV6bShQe1Smz3hUf8pmYGp0wqduCOjvQZheF+76mUgHJZEB8GCtP9UYPl3QnkckpoC
wJBuLHV7mW1JBATAMrTXX13sVU/uQ4NIo0C/KgL4pthiCJIzqQzizaBcQAS9Tq4R5444z4PJVHnm
6wnRdWhTurgsI3L2IB+2RTmYgn1Ym3fE2gaEISTR5tzN8NVeDHk7cgti5fx+9vBFqQJOu5jZ1IlB
U6HBZcooNWAvJJXYEl6+CLLIr3DK89pEWN5cG5b/agWoA1ZtV3qvDKHJ/NhEGIkGqNniADIlzIZP
8hAqwPA/8q4W1IvLCixEZnW6eEutujTdmOekzN7oKGOdTOlwXe+mzVzGcDvkSL0D1wGi57cKbnOR
yjs80FRTFKMwRrFNICKZvcBiGWj42eRMXFnNuTLFjNPB3lMCHKyaJ046u66lPd+HxjZekgdpGpOu
nJxRDzCxrjWOo+2ADzlKvas9GobhybcJY5usN1nVFFumEnEH3qi7njWWc38IeMTVfrqcvKusXhN4
2uqUgRi0FfjUxKAB6MFc9ZI6v2WQRZ1VDixO4wdKOdpbc44f1qbfkQXcR484iSRQgMZKznVBWoif
uxLOQIf9+LdvYr9UyJejv5V1FUK9s1rHpz4uu4nPgVsyVYv6pcMDMbv5fhyOihFMSrilEwFMSk03
0gOFJSeYNtYgVCxbG5bJKZfPYav/zGN9j079kKMWlWiPHgfg6wd0hVo5p4gQgVFn5o+AZmFCOXaM
e3aNYNALv9N9xasFc4rqfxKAr51hp+kPlZQjf2PEYdXXNKNNxQG3yEa/mi270C0E3Rn3abT9FTTh
+dvC79Cwxk0WNWWGsoeyGd55l6biqArEfGRjxTNx58AFwlufgWK4SWUxk/6uClFPofV7J+h1rzMd
CYFQQtvTX5BI0MwR7RpWnOfM/F59gjl5owjx9w47Ltp8aKRxN4WQTZm9oLYeULZ+/A2Y4kJzYn/E
Yck+awEo/QSiFCxR0I/OxM1wSj7ECmfISj2uLIKmbxuyylQkAtuVSkHtDElY+sKIzoILt4RK/Vk1
hPDTEetJedEauPsFjq1jtuuPyWVnYj57eFL20TLM9quz3OeC6XSUWRNFi42haY+J6WWFyyb+1S6g
rEBJUXwDBIdfe6tLozFjPG77x252lG+SFxlVvQfYs6Hu5adIf5rYIaUqb+Vy+gy6qXsDgWPwOEuD
KGFiUkRPMC+5eJfg0T3GIR59uaOWdeS3onX3imNFqSNzW+lyYhDpGC2bsyYywDZCbReZcvn7OPMA
Mbu3MOL9Rbr555gUZSPmi2MeWOVC79L9sbf9S+qJX4FvaxfIv3/VsZ71NfzNbbLicOIgQYCbn6gI
mREsQn07tTd3e+AoxS3YsQvqzpawFmIDbJgZcyL0vkn3L8ga+WKeKZN6nPNXrBj9OHIe3WdFrOvA
e+X98gH7zTx3hLlA5KQ9TKhNW6UfFChkQIYV9W4fpYnfiwZQAlxB2Pj+Ubssrohbkyb41JgLaPFT
IZFkCcqhTBnEIyO339dSkD2hPqLHk4p40HOT86tsxpvHkHDuWEo2sCzHV7c8FT4IA7q/DOb5PivP
luHFfuSU+T58S63P+lyJpQel9/mZJKkcsZs9lA8o1qJ7qdg8tr7dnzGYbz0vDFUepMEqf7s+A4ln
qP6D+YtqVaYvYJO7KASQoqsBWFbViPfFprssFmrR/5I61KO9YOnmP4o+g0ZipjCbdPk/+SESVyL4
jxF/QsEKGE3fKDcIvuRwdBg8CL275nEUI5fSI7/F6R2c5Z1OzlTLoqPGxOTr/NlTYW/Y8Ix6CA5y
36GFj89+MHeRbY7iklV0hD4I8BcR15pYi54BYPTmSLYCjeU3FwCi/9GX21SQeYSNXXlDJLhTPM8F
E8jWjbuj4zRMZEmwlo9FHhKQFcL8RFls1pspxNiz96kGRgO0zGzI3DvdghI1yLrcVZ4wrOFZCC7r
juaacER2BIbKw9zfUQnHt7YktNe49or0lF/IPcFQANrU8O/0pK2VRFDP7Yiw/0VxU57CBGw4x5Y6
WhtuIGIdN+icANyjeYCQYJEPIUBkpz5qYVz3O5FQUJhH5ibQgVv9IcgMx5BdDDomBFs9fWcCSpte
AaEgciAxxB1nmagy/rfzwRtnGU1aV2vV6ijgJCIEcnq4MP9xpnQhy2F6SEhsF1Mty0cVeD892h/s
nO2tPbVl0ARq6OaR3L2vYhkjH5y+tbHKgVr877+Z+GkweUT3ThzPqoCTCb46QdrfKtP4n1KYZEOc
1ENmlL0EJzZatSA6hI9iAAU1MYUw0e/CoCTXnvtQcHQmWcJlZCo8zXyRtayyE703QACB462g1fgu
Jnw3BVfKzrec9/kT2FJk+DKtxP3B685dIlmXDXiy+KSIGIWgL1bY1aUnF+GzLmpWd5YnK4ULHieG
W4miseOc4qtJq3yYDkPNh/JLCS3QoLkNk6nYZIqNsRv7DSjbUdcaior/gKCuKnQ7znazhtKkdVZH
EKk9DLA5lvRlt3XMC1KoH0OgU8m84TuaLiT8Urq7VOt8/4uN8UjUsbgnplk3IyPu0U3QnG8IZ2F9
aGYJXzDGM0xlWZfRD1IG7MWoLJzqlybi8sf2Eg3+z9YXrc56/pTFNgONTXFf3gRymmLO8kaN5uwW
ERPQzlmkBtWNLC8cWWacKaQCQQaTeawyRG3aaf9L7V+Muk4Z99xzlCev/C40qnu2BoRLNJzc6A4N
0u6G+60DgRgPhOeT7O1K0sCve0mT7W8rPLvDDNNDJqBKmi9faYd9bPzh2Y0vo9ClHP3CXrN7QyoV
av9s15NdvKkb/nbC82ysCMhs48Fz8Z0zJ5JaN8m48yEepw/gOmC62+bMaRc02OsrSmHqUN4XhafJ
x+LSt2r0AhhC0O9wR6YSgBOUUX4+BPOvaWA/Wa0fKhB74ragrGpvpfJJSMBatYiS6+M1S5YoRHKF
FzFqGS9f1DzeAgSSDcntkWSjQSyJKVU4RzviXpB/jKnh25KXrOtIEu/oIfo8jmP9KKff3Ey1j21U
bnHx4C+s/VMTXo7vCnCzurviFd4QNXSuUbrS3f2IzdizWfW9oguHKOWxSZgVnVU6yiHjofzJYz9C
CClPlme46N6pd24RUwuHHcvVcHVDEo71cBKwzjQiVtajqqe1i4EokR7kpuACFsSQDk0jREWdpqtu
w74Hx12ZLQL4jqa/z0bcMbp74BTE/2YVoB0JcO1IDpvg3ZmMUgKxhmz31Xz2SDaCWEhe9po4CmPa
5+fEQ4cVioruRUHt75YuFNjI2og5VdOjJ75OrDgDf4snOgbZ0peS/AoOvNjW3+YF6dzSNFijcycp
1DEyirN4w/EQf/P0RFu1FnJ9w9a1KwIIqy1/HKrUmSxaZaioQSM+PEnMHNqXVg8Pf++H4baHwOA7
Z8aOlHOp27Rw52CsPQNws4FEf5HUa7gA73c/JuwDEhJw4NhnXqA7ud9rW71hRiGGL0iAMOTeS627
AP+TEF/uUMEkFBFg4RXWv7r8puA6RnrkcdRmEuT3jqYPEfid6teEmSHIN6ZKh6snUbXPdoxQTSuD
i6kr150fc32ZhOAvbDwmRn7K/jq3LZYk/LaR+sV2MQN45AuReszI4Bu9jjqCsaWDpYmc5jsIuQ3u
/mlzwk+N7nQqDbrPqei4MfTrHvBJG61rqbFB+tZTSxIqJ+0eKdKRRWgKe4f29tsXHNX54B9EnY6G
8sytjrOEWbJZek0+yFX8WeBbNR7RVq/4m/mU3rzEp8tLb78sWtyrZorSW0BJB78Stg5qSAZLEDrw
ykJawHUwJrlkK6H5b9TePauVI4sTooj6TjG9b8/4MZA1k/9lIfxe9BJIGPYM92w7AhhwZ1a9rN2r
5xfvUNkhBypXS7Ypj8wYvcQ0FOxBbPJ/uexi5+/jcAxujE++KItYKa0Ra7PvEO7mLhH0EzDNaIVN
mRbqfGDTVfwcyfCDX8Am3RrcD+0q3iUyraecnO+B8NJM6MubJIE8QRRd7AbQiPC4w4oZIJ53y0jF
BdHltCc97/ynu7l6RrBISym64B0q1Yb67Z1xqk/F1JlrPPRYJGCgjchf2bckqYZCQbn0k8m1IRMK
6Q58TnIy8fCMdDD8IqsywhNaAyTimt2P3pnbLVDo2dqD99xZoz+yPLSI4dFWFSXXZ110Z5Y4Teu9
aSKm7Kd2Uc/FTieAZzxpLkq++lClViN2v2d9BHpKuhTGoURBPB/qhXCTMHibUmr0fkALEHEucR/K
Qd1qK+t0f1T9HubOZ0IZUBkdTyDasXl8jGt+0TU24MwDBu4WBTU/O1Nf+CCWCaKoGdZT+WbBXMRD
/12cMsAYo5Lx9Jwm2diUhzW6FSv8yR7zWoTGWBQc+4Tu8rXISPi/+3EH3uy/39SnkA9AKVydphkF
dcwK4s9uJFFkTvJqNJqPxDAcZYszfTyceVMhbB4B4ke5S6tUxnn4LYwErI8kFy51xUXJqda4j51m
n/rrziea10ZQ1eOMBCX3KOFcJltx7+Blil0FeRFlwEy2N9eq4M6IYGUWlD/8oENjxLIl70JWlV1x
b+PNUDCuYLOcuV1WdBoUOrI39RoCLbcEK3IBtXt/s6pyF2WmIuxjdVc+ed5SI+j7+bCxGRy6Oxao
XaLo3qqlCCAU0CUzKm+t8mvRm5XIV6O1kBpcp+aqGKVuxRvmftI6QaxYQ4c+Ivrx2Ihu6nrfGJEH
1gzjkYlDBVEdbss1Hr7LvI/jLAuQuOgbGEP0VlMrriqVI4ttDnhqBmQrN51dNegE1mMJst+Y4mXX
xOh/feZBfYjuedKK19bElIZyV8Qu89WCE9hSnqKuVR+x3v1S96jRuHWMtL/iDOFM+cW5+S3NB479
tnDa18olCsWJiYVCvaJq6TAFHRB/8mbyfiqbQqKH91FlULiMz/CJIXg+pVNikYXGJq8ZWuJeUa7Q
oOFbhTlH5RR2cj9moPk9s0yjlcmdDyzf7005wxfEu2jsFUmuzVXU3VL4osq8FVh2o+h46XDEaRfc
ayIqX1TdxaB31/3YikwBJY9W0A+Ye5gfI111Ae6lKIaDVt6rLWYxgDc5j9008AQs5jsbzPaQedC0
TcEQYnpPWEhV/Vsbba0cdI1gzpGKpcWsWzu3Vu55ZerCflqQdtROn+epUeETRbLxMxYIv3l52Qie
PyLs0RJW8+597tWHQTlljF9D+Hfh0XRgBxA9cQ/azOsr7joVJmxqTBMyTAX4eE+CYHEhwmG7zt5V
045YueQ3YxX+LvuwYwCoWXKV/jmM6UR5vw+4DFRJViZS5avxq995tmSxfaFfwzdT9A6aqwF0p7UD
Jhf1gM0l9/thoP2IlaUFRSia4tT+g1o1ivosxvVWjFp1mB9kC2HEdgK6UGAsywVSAADggr0qGkxA
azQ4/jzAZQYYY5wb+jhXpui3vE1p9K7dAE0NP6PvAxGu+8lgxTFFiCuqcGGapMJssH1zNdqqENve
eyRPyrHNIvnBO6UQZSiEDk9eJRREAShDdYfj7AKFctIAiucPpdu+dBsfCKUk7IJnaPlsO014Oa8t
81OtGd6X5yhFySM4tWSEuh8UHCDqt09zNNSjChEPysMKP0XC47nD7IBuTVT/R9Xlsiukyp1AaIl8
qVQsScantb2TOB3OJ6E5myts9LQEixaucZEyNmAfIyIu22qK/4e+UUiCCXDg8r7GEIwoBqgI+Eiz
kR8LlkI6LNnHP93hrLh88w6o3ZNCE4VpgFH+YB7FZK0FkKRkH7vhf+CnyuRa7pD6r4Cep7WpwoJW
kqs68bam5U68Jgtgpf55I4gS9OSZlgR+qEe88JKMt3AjeyBfLF/gMKgzaNrMXFYtgfORshwAKp4t
LOTzqYekibjqYfZhkClWiaWIivcdrNEDTgwrpG9udwjWxtZ1PeMReWGNu2LiVzj47QbMRwEWmdzq
3AA05OfzrCM50VPRL8ZNCraqgZx8n5HmQXH1JZlCJVkfREYm3dMNuMRY0a/McMY1migJto6els0c
aEDPLdd+ZHpHEV2+PZ1Fcy8IODuERJMNzyQ/4kMiVDKUk+Nh8gOOcVNSKLE8r23j8cFWjHsNcOXe
qPjTyXilsi4ubs6/CTyN9bhCEhdqP0GwMYkscdJLtFn6RXaoI4zkOIDC4Wbssvky83HZbi7mIkBl
yK8AQexqWu6abD+gN0wfYrew/0gEiWiUkGfaBLMJyR087AWiVE+lVqJfIaS4QQvpV357p/gJfIu2
CaGVoz10Z83utQnmvwK/c3GJQ6aHRSV94nTHZGHzj+ngvCZEf0C04V+oRRs+6ueqc2lwFq6LYaIa
K+NsXPIHQA5qK4gYm970Rwvoe/cC4ng3QHLn28ustWo18fBj9pzhfQBkdq+HbxOn4fRM3xYqkux5
DHjf8SyyBaeDaCCiOhIrdaXpiCEwsEQHWR3IiO865u28xZtfWgZ38n+VfSokyd3h4Dl2SGWRPZcR
tg76TV0ylR4cFyXspm+x8+f2T8WuENfzfoIkWaLSwEm1U+agip4Q/7cWvjdr/5shVQJhP60TJAok
ETlbOOup/GTZYoIlyEQy9cWd+zdohHgy8PiKjTVzB4feoK0n7Zp1wo8odhCw5phAJK38BIDaJRmZ
+JTOSwT/9VQQyUOdy1JWtiyKGEK7fitQU5EImp2XJRylHVede6fbOseViI6/59jK4KzcWGVpLWaF
G9UXLge161qB9rmXapWbz0FxYBP14VMzaAz+SpqZRc9P7OcywBjt9WAZSzS192hqSz+I/B5MgL2C
O+C1zzrY7thcNBV5g21dC1jSWmSSB/IQsmiTrVFtjh3bJEX2Ie3i45ZYL8n7xur2yXjEFzP2oigU
sSGyr+CxonHYVLEYqlJSInP4/Do8aBSs0Y8XCQmeD6ZWkGlEROP+C+1y/13+/3PLHEsm95LUPPmP
7TTQgJHwBNlmRXNy3OU4s/LuWCA8Ga3pws5FWqZsPLnVHZlV60wz174xxhORVoXEJLNbszolpz00
rxJ3Ll8LsCgRtYzQ0VS6Qtyn5jMq4CAlgczmtKwODjhz7ciTC/UFGFDm/DaH8EBI1wpmIWniiRRU
t3zQ8u5sp+h+yvEvIcYhjsOY1EZ66fuu4lDMTbQV2/g4PsZktwjlWkxNCQ/QmCBcJfc3yYem/3L2
aX5ivpmPpAH0e3T59vwAgrG3IZkL7NYsCECF5nD89Q9JEGtGrHbXmNCbhKZ01rAlYGWwUIGhyBRa
C5uwiBZ0vZxnKZCzlqLucV8jENfUAs98eeBYN2vi0ZSE/iNTtMBTNw3uDBeAsqdOUnMkbANFiDeH
Jb5dj/3WMJiLDxSgkK/BrnGNRiOW3rb9+DV+s7vbRY+IW2tfxx4BSc9sIgursm+zWBfXgyCPRuaJ
Kof66UsjYbeLKpDiMJx4XldU4up7gZ+GhnerMMbPEYPosTLvrRM5mD0LCABWcZAVRS4oxkxkm4iW
UDKC55IErbtA8ifwpFi3D/f3ydBRMzFKONuiA1K1kJpOUVXSKSy82QzUbSwxv9TagoLNUj8mIMFM
kPy/g6so6fAWJm6J9LBxufzmysHIzqSSoN1dn0LoPddQN+wNYpooGAF//+ObZaBsop0AIHRPByTA
+YIlaJTIs7sn9RyQQH13HGOp7wwjBE3ubF995K3sy3jiF/FmGz2tfy6AvuLcIlfLYxUykvWyitry
5V4sv+wQ9+8C0eJsfTUKrnm3Ic9qvM5eZyqD+gX8GbWibjeGNABZYLpdpz+EiiMQNN62TxXrdTUd
tKXGRb/bqvW3jglzEnN/mPizx4D76GmSJMOf0M0eIa7SHxa5VVBRKXyxjZOz6yzblL2CeQphCEqU
FTDyeUvtyAQ2fpzN6i7ZBpKBq6jrq0TXe8+T8TF+Pl+LwmQune21lAja3Hzc9tDbwSYdlIvPtVec
EMAB2cjA7dgKA1o1CvGi16IDH27OvfxPirVbBUWau0GR8sLj0aUBOdHExN/a1Dhnx33ErtdPxHTn
N+GPCksEtbumygKk3HpFTh/0KrOohebYCz1Qxy44NfSPefQuxgYEUcVhv8VqPNOhqWxR7wAFwJVP
Ej9JGNXzfw7daOf/7YpDYltV7tMeF+u8QI66ZVjIrDCS493v97dLA+7QsfxtIrgw83InD24Y65IF
eblP0lSGMueteg5SyFFDhzJkoh03miU3OskuJ4ZCUKTB45/wQkZkh1Ce0vE6/NsblukmisysBCPW
TH0onJnSrTyaGL6noEpk/mFI9dZs8asbsmIJURuIO2LwRzNY03Ng4+o0+KaUevcF8D84SfU2Yp5e
23U51bQmRP0OSKLTSaZdOUKhXqIQELovo4dZ6TkronoHwkO2RauYjaAPABLnx6wdmxKWwSAtjVJ6
iO9kBSnhiLLdH1V08WF9ZSV4lq5SH6scwZTXh/kHDwbyds702YkQ4Dm9Tc1Z3R6BBtutp3Hxca6o
PWApe5fMv1gUqvMDb+g90cKgTpJw9Pop0iMBqgGkAr5SoAoFStb5mXjVpkeyFNuQvxMRmtlTEh5x
oYVLxVPfhWl8yjCxw/J8e2eMd2LeEHf+ySpOf8puMM/EGTVi8fh2NJjeg7+gqYWiV7LDlqiU5En5
G4s0nJW6IrYRMuXyKC/orXemIy4FqFWQsheXg1G38KMdTVNLtjgVqJD1tXUJB+LMYJHvnOpnym54
8PYhfbGCSCXxKz4KPJcPsE4M3z9D+M3inaVNDe7oXg15rEq9aNwmrUBxS9Lw4jvRwi47muS3IYDR
AOBXGlHsmJGgkA6fL1mR+bxRNt3LFpzy2NfdCkZVz3xG5M3nusbHaHg3QYStkr2K3bKJsbdILAVT
STiYK4hPbDCU1eiuMzy6WWggxO/HEa5ZlH/eTHfjttJuIaMy+c8NRGGZ6UcIaOJw4g7T/3NPwmUT
ZtLcl512bAj2x8dE0BdEtFcjRc+P7krUctZgi1qtM9WWVcN7RnehbesAjsHXLwUD/ANyD/pEmxZD
VSQvloNGXZB44FP9+jLBlRXeSlx4GZI9Eqs0CgW+vr8Ndwf8VAerGpbALIGCc2fi4ZDcd9Bysxd5
3HAv4FD6y2sD1/IoBVI/AcZ3Erw9/RuNHMsJZ3qb4ZHolpC+6u/6lXQOckmDrl8VTYgz0o6Nc7cr
2u+fyu1zTTm87ptihez6WvSSHlg/1dRg8LA9IGUhMssUqJn03E5j1MGnd7PDlGlpvrn8r+qxJDXm
WtHIDTZOGsLoZ6pvrl1ws+VcTP9zZ3UVU3o43ypBxCj4F278vXaMGVbBprKFYo22eMM5nL8kZHQs
HewjyCv3+7Scimn8dtyl7HQ/WPm35yYfYafwGmU18vmkPDMm3DrKIBHPegFLh1SoBOherZoUV0Yc
WMAXVgrOq55HYed96dTjcCKZHWKkBtP51qLTXCUwEyLAY+8odyLaeQTwJVUUa6gajC9tKvUvBTSX
raCF3P8gXFZOU5Ftdn1Bcuu2BIe0hBDzk83qh+HY4IeSX4LvBkG7Ye6tWnyKli7s6+IaJsSXc7Aq
YZaYOQNmr6LSj8YUDMvFCFkOeRv6Ouj5y5hEcJXys66LDsemJpZZlWBlfwvfzBKFsviNvOEEKbE3
5GhY07hI4VuD/SqAOXlxKN8VmAt8AMNCoR21xRV/GLs/shRJefxUNe011S1dP/6rwMNERnKB0G9i
zCWRJpaMLksJwWmGicyJ2hZzONgH42XMRXFVq6rCwhdG96/7hTZ2p8Y8hcAph1atLwvHIbmtlBbD
CGKujzqyz0g1Z4cpLYHuTVIjwpTYDctGeQKRmRhUB6YV4sp5F4j1FcZpWOzl+S8jyl4Dmvqm6H/k
ioWF6PTLWu4pA3W8tQCa8y31wyWFdIRZXbotNVsQkCGcyil4DIiBU+VBX5DHjHFdm1iFZPdvMUTI
vW7nn39Uf1QPfFrZ9T+1fYU/C1nt2O4PSUHYOPqjL4cmzukmt3YDiI9UouySeYKdc1vQQCycwhv6
bAk8ssm229mhCNp0pIy2c7gbJxL6YfbzeDEmMpXOnXpYlFQX73qZ6I3LhqV8ee4jtmUeGpATqBj8
32ZSu0yg6PG4TzRnsKBBhnTXmm0cx+e8pmTuA5CMHFz6CwuH7zTe+23hshL2GXuMTbMXwOBwGNvS
sLgdwH1gcwmo2KZdlRzxf1vpOTtJmO1MOu6gVe+SZSI72L8slunnsiOmm5o1ngqhM5NYJbejLvBz
iGQmAOerq05S8uXL+3jafJqUtLYAktdf6QVt71CovoxaQYlN5zD7FW3MnVclmB8ejPvvAFY6zBNg
vUjfNY1rI8HOA7INkDKlXyykZaIEartopNPPL+H9SUkz0KyuUTR6EpJEctJwmfuqQvd7vA5XZhtu
WfkvIuOnNax7Tho34jY69B/OiBKI8fNrk++VF7dsswDrydBJSLQE8Woo71pQ/vspOmQtG4IfYtNq
EzFXH1eVdIRsbHSxlp3As7nr8nxvPaKquvEmp6S96QkIFy6DVN6sbxp9zTgkYv0cckQhhK8eX5MS
bch8TVGpfRxgbYXCPCwmC6UaNm9lHmTjBnzEM7Ipk2doaqvfe+/OvaTAOOfUOTFyElNpnTsPibEW
+KoJBZNCzoZSr/8kM4s1HV6OlYv1Fkwzvz4yie99JrIQRRStvkW75S+b/AOPOJljSGdKh8OIA0jZ
cTbncmo+X89cIIQG1lVCUbyByP+r6pL6CeN9uLYFDdVG27cm7zHf3PIze3Bf3t9Wu6QUJs7i1KTN
ip2Qzojyv/WKQmrj02WZpx1flS+q7pmatcPh6VO2h5difcYZogAdxXqTbV5M8GaB1XKcX2PUof2L
9P6b5mTc2VOowdR67yecdcTc7/7uBCXca53cQ+eRuegnSIu4fllXllGf+3q7bCLbm672b1p6kbVc
nzFwqffgi1tbS1GtezEdUVY+ghBlVSEhRo/QhpH5EHzH4tG8yv9rBysKiZpD3XCWqnl1AFU5DaZl
OidMRLj6TsS3Kf7fCbRKz/pLKV5ywJfkYuwpoUR4NLc2aT7wHz9snCznTLTjcmlQYnm58G5Amn1x
SqQmiOrBALsam49kow80+ei6Hgagfj4dDHSX+25ijsnprqE738VN9Me2wUnCAXNFGJhNXRNM0WzY
SWLh/TW5ZftZeeboa2GYsZlEW74wCoC65BYrjVak/NGvlWjgn98a5xAM+evQTYxVqLtKXvli8VdQ
kAFCFtLqRPTmD7RIyQ2o4V1FReGEVDHLtFgnfc0J07skuoLROGwkre5pSgCHAl2Hd28VK8z/Wcnc
aqv4m7YdrJ/kXi2L6Lq+WIjQgkBhYCEzJ65OpOOnEgpmx8MCm1JaiUXBy0L/u3fV2zGL6HS3JW3C
kDWazlCWRszXlr1NHDg9KF3/Fa2BAJ9I8jJtJ5FxJ5p66W1JVK8OX2eiedh42tdw7m9LOPgvdVd8
8uFpjuquaApccyWWZ+2fcJlhdC2hq+7+DfTGNXTXgUS/5q/lBjKy1b9YNkC3GcGREnv/j2dvkKML
zXE0yWlQheX2dlE3riukBbFo2ftIfIylW1j/PWQT4DraADXUt1j9YotjpAD9RLjvG8a4iDwxCMYx
lhKBNbOtgKNagNW2L6wwxruKxzHhHGv4es20rwmqj2JeolLPbPO0t9DJ8yYdaKH4sewAnYT3uUUL
hE4bFiASQgYUakOr/bWzWWIV3SGzFgWYny9lSYhgEaEU7/oywGenypLXf40SimiT/U3FYmJR/Hc/
O6WoalUqUvRzzwygx5n0sdWoLZKMCfGfzHy+tj1tsQnT+VZaFWD+qCCX2t022dzQIbajXEztNrMZ
lZxGXo264OFEMA3Y+xs7XvDg7s1ed/Mz/YJAkT+z830nFgEPdRjqCyA+Mr7BgpWP2vELRn2JxYCO
rordzyOs3r0tDQ39pD7mRxtQRPMz0qDjJbMdI8nEt8J0sTg2tw7BCAntvHFKHmkqRjgt/zAkopyH
A0+/rknSzJXwvSSVTd9K3CbkYa3x6Mc6OEE9pxjVyV+YCJ7dCggsl5Up3QxKdE2sNwY4zrdDkpwv
5pc4RBjMug3sFoprZzTsbWEE2xk4GUGjsirfkxUj0PEFBUtvwE1iEr/3X0SAcCi4IhNihbaEr7ls
ccg7VKtw+yqzZMLIeKkZPShoW3XdBrKgerqghzHkCzMAqeWlUph62udvZ3rCFodMg0pc4iwvEcgu
M51KYxjHj2rQ262+LghbdnxxI3tUbyIgw0J23ITP/b95dlwBawk2dMiDwqe7kTZq+l/O06bVBkF/
QE9y3SPlOsBrMqPd0fwiNoKbv+eJgGMGKIBA/SSav7zVAh0g0pkoyx48Apxbqt+coTK1yUSPBEtV
3y/3sMUrQhoEjeRJWR4v78v2rMtUB4pPmVevwTbApoHB+BQnegjsFZbSsksWL2dQiY0rlGdowqLn
1VJuN3vyhSdk8UFb5D03vZazdC24DBbBkppgTnQtbKlayCQoaUiwKEgX4+uQrweaz8fk1iVCv6dV
LJB24iOmYqebVG7i4QbKt50aCfj0Jur172pmRnTfMHaZY6fGXHdHxn5eToYehgZlFCwHLGk4Zl8U
+wrfs5+oP85utHfxpwmw0FnG9m8yVMh+6kpXA6m/r50hBY5lLA0PYYDx4PS6h+EtmUFPxC4op3Kn
kaMXVnIwlJJcmyYswb9STR28H8XPtiu0OJp9WoEfMwGH/DekKKZrleWuInWpzaax/YxBrc3ZiQRj
SdzjdkRJTRDkzX0l9hlfH/DIeysB+nkpdWbgpR5S+ERec61GFC0FBHbtOkjwsz2aA5e+cybmIh+b
U/54nDwn26sTF5IqdYQ/B9q7fDQoSbW+a1tX0Jp4miQgGgPUwbxcYDJnWSIC4gErRfwYRB0FI9NL
xdTj0NlSN766msyPbp7NO6RNotQICWPM+OkY5/vys1/t1TiUZkJXAcbdRqzvX4++Q23cwUMk5Z66
Tyg98JgE6QR7Xcxhb9Jx2JlrfMiZ6x0rFU5WuVZXWXyvZyZF7ynoOL6KC4I7xuwpYym0HHW+AKnf
oSZnThM8MV4GR2jNDcSga4Wqg9HY5DD1dB44x1HfQaFpwhCj3txQhgQ9kd5WKWe+kwsLRM4i45ch
bcw1PRkZo6NOeQru1s3nHY//5xStl1y/E2S+1oUEmSNTomDRDpuBfGYvZDdeX7HwS5jmgOM17rzD
VTQbVQeW7SXWelsso4+cnQOCy/B+e5Zp0y+i+NgEIAZ3Yk2C9Ti7DiDDOdJlMYwnS6FVHRXveNJK
SIff6tOxpYIehtcKZtGnBJ9lFCdiFqLR1PhnpdwUJs/GhzvokDlT9zs2GqgMNCKh55gYYaBk7oE5
ntf0zYj92QX/mSlbZ0VkniceHoymd0Ld94eAyhILegJh2/nGZHA5eySVhkVpVH0lc6z3TfJKCx2R
QUbAui9VaU7S5Iw8kAjJ+s0ktbh5IlQ8mUzg9qUYI4cA/30I5/XBWk1k5RLX/nQtfR6lMrssI+vz
ttGNTA3CXYovc4hGetrVGQzALWIfrF+QyeygPffHOn3YvoPzyvhdeymLASW7hzJNuToaqwwd9gdy
s1C6UzNj21hB0lv7CBJCEa3DNv1F6aRhPoKadhfbaY+RriAju7C/3HnvWoWoFOMaDeOE6OcGwtyg
Cw2oZhbB4rHq+qiA78e3M8QOKMbw4q588zuen/XNGBXGyCdShA7B1KrGvYRN/G5u13jMsej8sVOz
2j3uc+OOIxZ9YrDs3HTNXKl/8iLmM5pMuuKx0ugyA16oQ9j14/0L+kV/tvAVVoTy3+yWycWfhm/4
MurSFnNbE3rPZEVMYk8Izva1SzlwEcn7ca5jVc9+iLXuRaBRSZyC64uYvFhuIwrWt+v/w4wefYuW
89ySAReQK97cwL99o6Z8RUzso/LMXFcVmbtPmPU7yOIka6fZe7BMWlsOS5In2dya8aotaWLKWTGv
/QE+evNdvxkFHYgU5VjiIe5lzqtwaQfNknvf+iOrFbqT3bcqrEnCAQw2yTeVcUtZel/W2kle0M1Q
m8Y7MMNP6BH3sn1Hg/enWx4f1Q6nDxj1PDuNFay6voyYMQeGKuaYGsmx3/czzDzAssgjgzDxzwEU
e64bH+nhCJE64ERBJL2OyXtks1na8ANhTfcOPMpNN61jljPbe5lRVsm37d3ES8dWk/ql2uFhmrVd
7vA5lfRe8AiBwWV+AOdRl7ZoG+k+BPLkDdcG7asnTRDBXa1AzowaIROF26Zf9AQ+h7WuSRQEZbfO
/GmKgzrP9Tb8oWqrtK/Z60rpNGnq4kW9s/lX5vZchOMlyxqBycHBDlCSJRznDQ/b2MJaJtxi/zTb
n7l+pQgY3gNRYVkCEUeEKMpxTZedAFPulVq97fTQyYc4Kxun7+zLQm4/cyRRpCUhSuQUcYFDzyxu
MX8c8CEcad2IAPRUX4Izvn/479z7u6zYbko7+DtO1BQuZbMJ0/9OfycgynlNZnvIwlLwJmev57eE
YIS1Ad+6ZGhk1kXCR/cACBEZJgZFQH2T4FV02/SjKy2gpiyH9Xi1HsvMuF/b/QN/BUtys5Y0a9as
SDxkdAXfb0hFPoEM21JvTIxNFIuxeGvxdWyXpVIh95cwid5tNdoDxidCqV9+GntrX7caKMRnuoi/
LcS3bkZDyU/IskN3+IvbRtN6f4MA8HSkSHRO5dF7xkfNZR6roDKKefZnC+NMr6i/troYdAEJaey5
JcMho1oeJFEtLnSoXzXCySzkdN2vqM01t+cnXyjqGhYYDQrCKlETbWwScDTyHBYROjqZNQgEFrch
EkfiHlGZ/wLoPTaEOIJYfosKPl6sL9Y6nxsEyuxBmnLBE3CukFs63k59pAf7thhEubeXjQf9GHR7
UF32UpKvcALYAB5vnAhYl0sJDXKP12yavLWndvUbwFpMBP3VxWsc6ybHe9smoqa8uegpxG/ypyzO
cGvxenPt6nZVT1WFrmVeVBLGbsK+uFPGPF26kfSgpaKnwABsY9DpIrI4HnyFfgr3SqCN5U9VABbi
WJjELkzO1ScPtS12IGY+NDr/naTbGDE3lCTuBdUjcBFeMoopXPHcFo7i/rDR4a+CjnzaemrHJNya
0thrmkUircOTlXy9i752y7vPrGlcfNeXhpr3GJBMX8GnfvwPkZL37VTvszt5+ZnOfVL7GbarEmW7
bc5GNlvwt5yZu/SO9eoj69pSy2mwUzA4LtSrS4YieTu7Q8+eg0XgC3cvhXk4HzCeDxE1/XMplvgw
CScOFkz7XI+yfAOb5zWGtLuioc6zTalJwlNQInzPk/BPpD+fE53SjiuRhypAgvHv1PicLL8n+RjB
C6xH5SU/L2/z7j7v0YWH74G4WNzUMfGBIZJ7yVbzDeoz0Rw16RTUgZUqoXEp8lCMF4MebqaXxheG
xSkI9LmJVOyvBp20YRD7Z72ExECcXTQy2NsrVCFh36icBKZKulqM0c9lr/BWCwMkpyIPBWKChq0D
sxndfjff6tDubIsUJ1sJ1S7rE1tcD9e0v7GED5MiUWN0r19B6v3k9kPUYkgsACA39y6Y0vtr3a7s
BsuLv4M9jRkqatoZaC0SN5ug86H6FrcIN0c9aJBBBYPA9rzLi2rRSMGlBR8KRZBz1Xjd3CV2RAt/
BEiyyzWwLWBvuVAYXUFIHMoJ1HcjprOLTjOKAGuEqj24FNcUzGWSA4aQO8TeG0F/6iG2uUPmsTA8
d622/DWJTzAng5vOiT045dc2RVEVJ4LbPBosZEWZCvJbt/Y0yqA9hNa05WyV4H5hOT94yEDS3wc7
Cwy3mcjPLc0c9514KHlF5QOod9af6lM4nO04v8SEGpPI4QfjtvNeMb82gpFVoXf5oKrEXKhNSjsV
AVOwSHFpl4ocPRksXzra1waGi0RLU3QnWWeFtssok1XdkYodkXPEB6XQ7ao38IhxYnIZu1eOtNF+
Sa5Z/wm43rwCmPcs7mMxcmXJeB4G3D17f6miRKgxdUcB+BpUwFBcJeh9f5cgm05B262JUOJRNN+Q
mbm7M5GfdYVLN/ENXf7N93oFIzwEfgahZeeg5LtojMDUiaPdU+teNr4Mlj7jt53g3eKYCJmQPEjY
HQrv0+HNx/Z3E7lNMhrny++P3rcI9Su+uigRtbs9P5tteJOYO878b9MYwr9JCbWp54v92gIXw2LK
n1QX3QOw9A9B787EKsOuqxHOoj8WTeVrbMZMSF91IBDqF86tLr/M2w1Lv/6Wv72Qo8v1k8S6Xl3o
ejIZ3SDXhoenzrjq5mdCbljmdE58Rnh5MXiw36TJOteZvhdLGGkzom6uO6jm90fHuy+ldk/PI+mN
zltn2CJCmXZWWazoDtgsVIjfuB3A6EsFGrSccl6O+KQBzpGFsR+hnS6nmoTr0XKI/3v53R3m0X3v
Nwx/5ShNXxbf7Hxh8Ooe7kdYm4gmyMVP6bXdvhxwsBcEJhDPYcQskQmZDERC4q0bHoGGYEBN9UFE
fg9F4HJzcqRL+jno7iWG1h/NRRc5C5+k0xTtF4SpfwHqpUHT0uX52Et6bHyFYah+TKTABmuVb3Al
yQn5aOKlySJ+WAT1Offm5vw6Biu64SaqKT8PkkHsa5tmFkgqXNuPnp20IidrApPmx6ktB8oD64PD
PTdVW3Blco/sD+G+NWW7M1Km8SuupEyZNnjH1U3/6WvxgzeiRN5C3FH1AJ5w4JPbIQ2m1WtmegdR
+cNl5D53TBHtsqQURLxwRy2Q4BEN+f91ZScp27kcKzhRskAjFQXSwu1vso8DqV/7cjUzDA3XaZfz
MYHIFKsJClGvRTrZNIDQeJq20gV4H7MeO1V6VVupsg+7ES3mt0bAawCFKB8IQIckHXuMJezyoLYK
bBfNv0NwIg8h12Vz6pvu5Pa5G1kB6KaCkDdcTRCtUkd2A+AD3ieujINbgvu2ZA6T+K+IIn+UKBCX
VYxDcjgikW/sRm+TJ+vY9Ptl9fw+1MW7IS0VKQmaRbLcH928eQtnenUt5v2oigeBYjtCOGmzTAjg
jIaI1fnQDHx+Iyrx/xoESu+JXLSOkruLtNINfYV4LbOeopsZrnYj2nVEDBAQOKWWXPk8EEPUpB2k
29LYTfU6l25oPlX8/NigfiiRLkRbI4KWvfUyd6Lo6wZwpPQu5QlTRMTIsxgsfvFpUhxGvvrnEkMd
5Ra0qb6kTAXy6xvgkOYVB0GyK4tODQZSj63c3rKiyWn8OL2cjOtXiGnpG4Wk80atope5o+mjuFFf
Zgmfx9LlHeOMtqgCAyE3uxEEt6W1W3DoBbd7Jk1W6RV5Sb1bHHahUJTmk+W70SmmAThz6ftz10SP
fjBso6Ns9r2jhVmu2VA2b6ghz3EmWxn59g6JxjFITu+04qPSb4WEDGgo0/QWP3oVzmcd5jBguhWu
WllPSJVVwsrGd0PQUmo3TWhUXpjAn6j1ItgLrDcZQM6HKnx/UCHSiRnNmm9uWc/2RJcyfmq8JxiO
EKvptBgs2/PpQSTle1QRRfa2a3tJOYwAcG8Bse2eS5mwlhXDP7psxcwyYWWVuvrOjCFEIxKkpb2b
sXfoiDOUKBNzoUehTVcga2TE93TVuP0aN1Xuo+OLDvKPXAHnT/y5m7/Ism2kc02NvalPSwpU2Qzt
nWlG0I6VfeRunvCTurH5Tz9o+NcwHQUAD8sTxftUaZQzjYLrT7LiO3RJoLa6pap0QV1c3rLMsSz/
B68FE46JwOPXUy4/Pyb9xqxsHoKaNSsrpz62fHYvxjTzUgC+s5VexpQ6ezsk6uP2DNM5UBRpd9kq
519ZftKo/dUKM1zd22aQL8KidtBE2iiSsOFHIPCfqpK8+hVeSUZkKE0vYvrjVBo2NWtdSrPb2v4+
tdCUB6suuF98M8oBaV7uOAiULaQXF7SdqFC/lfuZJZIFw+NV6VYBECiFCqXPxOd8O7//olboEUsJ
m0FaAn0DyCuqLtOUxNYoJHC0yBJGEmr4lhtj9i6RURoVTqkZF+u/FyyKO7zxH78RKi8GiwpxHZeT
BLtd3SuVMK4jSLsKh2Lt2Efw62j67CX9pipKlOCc/rerdTggBwv37LSufaLhbqJXNwBFzXt8KrXr
2dCUWvYmR9WHj9yfRfm3+9htCF6hd6/+JgZqYOCHZwVwp4crsTXiuGzJxvW14dWyyhZGyVEaRW89
NX7K95w5EgarnGFiAfBFdB+twvqAxRRELI1w7smCsMvnE6pHbWsA5yu1avvHiJOMgYKcC5aYGT05
+ODTwvdut33iw9ptoRvWWRh/ghhskMNQ/7TRK11arqqEym1STaSEfUpkyuat/bTVr7QG8f2Xek16
iQLfG0cHDIPryP1S1mupbEAHy9GUynuSCT9ojSPJHGGkjzmo3H+37HcRtjo1UrKTEETjUNolJ6CI
wUqRuXimllqWieCP18nynexv4Qf2v6y5yjDcB10xteX8ZaQ5nCvKAGda+HRm//RD5IbsN2s7AXCY
nYtNYLDxv9szsNv5paqdbOqK3vaKltRsce9buWt5bKgiGch6B2fXg7JJRG0u/FwcC7tSrjTuIBU=
`pragma protect end_protected
