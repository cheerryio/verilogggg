`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 155456)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCahs3fiyq/876fXZqyDwf+5BbIuoKlNJVBEiNW9mMuuib4kVB4yOdmIt
QcWzJU/NwKP32tAGbEMDLBL8PALQJchlSLBoHcwQctuvWSHbJKj1TNCoudwe13iLf2yzabmtHjJw
kDpV/j6ZOje+7AAIdtUfXC+VLdGII2JW8QZpvPYljN4Nrc23PX++Mye7LMLR7doE0T9TK7Ftlp4H
veSLahj39A7TriNlWixN74PVfdgYV/Z5BSF2sYnfV5p1HV+ecpG35iX5VCXhczg7g7jvyeMUnq+g
yH81em/S0r5SvqMO6VMVhb3DvG4fkr4jE4C5gh92PKwq/ZLBy7rLSBaMtPvDJnE2UHWFP8rmUAVO
vDh28QhXsYqVhRTkraSsy2wGdfakybHaKfjh/ZVZiXyihe0kknPaxRRevAmIBDCbEzi+7cn2V6TQ
lQqvEQAcw5a1xVt5Oc5VSws+4wrLuUWuMLmz1j0b7GGvp0W3f8LPTiLXHIoT2/AW5jlrGJri6wa/
2f+zepuSlmWJgzfsfqGxnRQ5SmzGOmzzde/CDBhtgT9Pm5uEVzulE7b3Z0xrxY0NdiCmFuZ+vJr3
Vu7DXCmOyCDOI9N0vOwG6tjT+959M+Vw0UVLIkYQuqEBC/W7U8XN4XOFeKdY0uGTmSCsYxFvBUUD
7dm/F+jyuZpzSTkG5vYU5v891eK8CpK5cRLZ8OJc8U4Kzk3xTgWUWxq0gsPbbYA3LK1UyS2ZOTLF
bql4zrXWG1zGx+rKP47wdEu+raYrz21VNlqEA7AXa0op7yyNx9QgJjSBiVpdjQUh51WXPwF6lK4t
hJ+Vmr93Wtd5DyZXG02uDxp/UkjtH/qKopWLP6xrSX63b1QBFNXR1hBmSCQhpxJ/BAAa/QQUWgUx
sg892uhlQfZBVi6MfjdwjqIBT5y3IGMgdamlznjrpiLKGp7MKRftB7KLR2OeqGK/QDnCvdfwq3PE
qQNnsdzhtpeMj/TZFfB1VwJ+QqfNsTMkXehz0+qxYZarigN1nGkDgeJtQlKbWxjS66qMNwikX8H2
+nlVH1vXfDU3iI35AVm1pIzNIOcG2X513hwUGU8rGy0YDYukP7w+t3GBshnApwTxjzGnzfoaugcZ
xuT0fm9IgKODtNI2pIlZf1w7wq0CR9OO1wbCg/9HzPxsOXUYoEqKqPc7c6cR1lII0LknSPO1uFYP
cxrAbP9/aOfmJ3ifOX0iRABNJspWcJCMhgw5u+Tceh0/SOe9NwCIv/drsnWOTzszjhAYNwgXH2dJ
G9by8Sg9aU4vQeomZqyG/VSFz2TuOSpqONWDxBPe8Z3b2lJNgTfVHdLdyLCLbMFtXKNpFjPmjWo1
WknpTK9FgLrelqGITLvGsc4Cg7mCFeMbGN03Yz3cXq/y8ROsT94B2b5uiC1ItBzu+4NMHPktnAeF
2b97ZcpnOEMe8J52FVjb4+3xGh9BlY81lkLSKs1q9svrWLrdIz5kwyTwmGFl4pFtnI4wWjUfAkrU
m5A3c+akg+CESNK2hNlktEDyldgi9WF1bIL5NybK+3owtLaM4LHQpy/3+xYjSPG+HYj53g+iGeVl
ZSZgPmcErTnpFTSS76+uVRYjYdb4etknB7AXrQ+nzzUTtKwPxlNjp3oinwL8CZv8HMKHwjiW7PfH
klx/N+8bV2mm/IVuRyidTllNf01u8SmiBjZutldcGhtAScnE/QlF+st7QL/CoHQk7BaI/yCEq46U
XoVSeKI8sICbgiCi+bTtv5giof/nYNC9Os6Z2CklGQG8lDMplckzc7Wq3uRXo8pfsk8wwNK6muy9
OJnZqMwTTjlg2P3K1eK68kvQ/IsVplGxki9W32z9B7FGQccbje7Orb6PWJLpmLt74axGPyvLse6u
tDM47+s9XhXz8jm+mQ/DHM42Dlh/2zw1ikNQxnTeVjRFtTj9AfbKAiJdmX89vh3FL2CZL0IoQVoU
kxSMXaOngFIJYXqyxiampay6RT1QRn6moAFktcret4xXWp9FIpq/oY2fBrEhQVECkd01xjNDpahG
o5txi0yHr5c+92faKYV6erSUNzzXrBEtpB4a4dNfUWfyU55iJ8nMRL5w9B0YO1ZncaCSg0tLL0vU
98d4JkV8PqiODxGpzsrX3PdAOwEuAF0Lqjasv2q8TBm0p80hgKqdk9KVKNVL94M9d8D69Vy4ecgI
xbsHcz3xQS+R10b643I9ldxwVbUKD7F+JU5ub+QhaNHjFsoISh7SCSIpbkndXcI1aKGXqYlfwTec
ruHXF2jd//409CbzjANHx7JFRAeNlQGEt4b6HVqYB2EnX6KmGP7fj8k6HmVtEjdJ+vV1W50CstZk
78iyLxwAFNiy8L6wL4DEsJBuhWk1v4nXtPzaV0BIqRub4ij0TZxySCrWR81HqdYtLh59Bkt/aSBx
PtLfOUJxuyBqtXXD5rdwKg7HppSGIUi4VVK8hTuTWnHSRm/MtEp+GPtGS5DvbUKumAf3kHCl3Vud
I3Tjtf7n1wjdZH+wQiGSD/7XOGlO6ZbQL82GdFid9+BJrbbhO0JHGPgHDI+pSppfzyVL/2KEfa12
FpWCCpM9eYm7Cjcj7X/zwfdxxlDwjr2mM0mPIgsSN37B5JhylavVsqIZBqB5NKDrWl1yQgnydubH
4GE1gsrq0V5m8sDPSn+Ul3WwLFubRQgG6pDySLmYYC6DRsKpKovIIoxrwemHGfrXtpAFkwao9Czv
PO3qt8Tn48u2IXyhH/5CIzlvzoGQdW65GIHWx1HI/QCj9r9f/oyHhUHJv56IhftFvd2Xo/PIyELD
1OaQax8Reo9ho8MzMxTKz0Bo6BU+Tlht6xTfDjlqVQrpVGASzgKcY41Ah5AlP7dvBg61f/I0C0Dj
VG3SN762bP3ExIjKrXHcJfdNfB9TVtn5Ttcsku+XkpL0kGKDm+QS4R3WX1ZgP72KKrKRcigoDYnX
aRzBgqzvChOYxxwgx6eRmNqzHi0m7o5qbM/iMbWpO1tZeJPh0mBYJiSY0OAl4dE2jFUCqT1K0K+6
+gjvYXCzqSY4XWrieQNHRuJMH7IXERQROxcDH7kenCzeDMTPm16yzaZkpdmMGcesM5Oab9LeHV3z
CQ+LQBKZRLkcaBpcmrb90J19JakAcv0e5CtIBOgECJyw1+U7xOJOOecW/Tcz2kbwMM07e0RAwE87
PxcJOE3E9AWXOzEOunKuzBDmkF88zrvnaMJpMCpQ7FMoERlchg0UmDzOUitFYaAiYnz5tqQH73ZB
KQWvp+Sv5GrenAUHKZNTuDNFIQRWDnqOPLdP1BePO4Ga60g1eBwWuSfCMG1PR2ciQeIWaY2iR/g0
oEhtBzkBHgKLBgPHWHuZMsLSv8agKgaVeCtdR24/hQVD2KoVjJmZ8EEDV3LBWN6SPl3+8XzOCGvq
eMxK1eO4i14Qhdr7LM59WsdkIdTFyV2hu39wOvAZNqxcqYOjvQgZFJePmv6lDZCZKZZghzagEnTA
+Me+31hqQdAIWFVXZEmG66liiqBPY6LjC1L7YxaAVtETJbgvU1H3dA+krX0Pfj4o8ZWW6nMuRGzR
76hdR4MXt4C2F+9dspRmoKaNEAjct0DYPL6JI1wTzdt0cDnCufwse2hVAjFTDqzuoMxDcJ685D5T
ScCZFA1kYfSVupca4Sbwcz9NYpirX9ymCb+OYhhiXetB1Il1Lus3zfxmGIpfZlSU1snRFskmHlT7
JM/A6x0Ns7evOMtREm22J6y3nlDuIQzF7ZyJsYLingnu3UoCtoP1CMxtyNnATkASWopfFD0JCy2g
FuWkpaMet2MU8YfyPeJDbdTn9S9GDW9GO3fS2JQJtPivW+p92NglxRXeCQXeAhRUv2eCmBr4/6TW
5A7RkhfdEYYFGErfTJYpsJlEoEGaSN123e/QhLda4XSfrLFiBXvARCjBR24rWBJ8PwG+ZPCxy8rD
edzA6/+JAjw8McLsKEtlvgTv211S8F4HBgfELpl8ctpxSzpDqHaH3LENd5RbVFsw9op2FCEMXmvl
QxcBLnEMuRIpn5QFrLqArr3P44Gc7+yB0PyIGTzWGKr3+mCpQw3y/Q95ESAU2RvvDmVb4wOJKalg
Ax0fUrfKO2Gn+46nXz7No62ioYFwCJtA2+vuUezpRl7+/bCNg15B3bPOQAEjjZoFibc1nyX/mrBr
p7Rbda+UEH/JD8W69TGhwaDqdiGgSYO+c50T0EUgbK5a87nZPwvvH+PtYMSBf+yqF/7kqop/M/7D
OwGg14nrYz77kSe9uoEoz36bL/hXEoqQEhJ4JUzVkKHAxTAAEtuvTjmE8I3rWttChlZQnAOKqPUO
XQfXKTT/+8XmLS8d2V3vleT78yP88eBb5e94vGgQCWWC+Xm0skk0w2SYydZBDLu/pcrdVJjTvGI6
2lAhjMM0KWG7k1uYguD/GzsT6h87DEu3Fv0C9LpZJqj4raIIfj89WZR4cLDFrMb2W3RCaUcZIyKo
ouRV7MnBv97WTNDA4DXUW/SVKTT71hFpFg1ziuRdXmIALZJbl/HnQ0mhfYPsWXbfPJEpcp51OHx3
GLnmO+F3mNZbE1XL29kaazCdg4NCg0D2w2sxowyYylP0nFg9wwdPPuCucdy1FO2fbxjgR5MkVOVA
EQ3QHH3Ix7ytC2ij++5osiqf8CjeTnp1o+Ge8Ls6ZXkx/mIW0vz5ggg1ef50g1V3rU5kAlGrJoB8
8gXKdQI6bTzf0y8mQr8sx3kgQkRAmahOt5NTVLe6lgoN/OaZCFiuzHp7+YyCZmQ3HiADBxPYPmhp
SVWHwHrpcww8jKrviOBl1kBe4hXHQO0wuO6UxZ78vVEM7CCfacvoo1ZbANLRyozJ1MNrFekXvME1
0+CNybe4ogDptTakVZF7tw6q8K5zxsoTBZbr8GQfBiA5gbtYIQInHYQnsMVbaboMl0+oIfQFffVE
M+M3+4RxmECU11CEk7WkknenVT3ARmLU18wVPK6yK8iB9+EEU3EGEF96xQRsSvy82JsRwkLTLlbk
PkK67OOx7mQY4qIXEMhnZjWAF9UG8J/Ks26asuLHBRL72DzbPFer/bkzTiL5ig6ueYJe076O3rpB
w5hDSBoBugTDWm6mQBtg4R4Wj+BStHXPt2zwqx7d0PdCbbQspqxPz9ECiwwGwaDS607uufYzQJbA
hnB5KXZs7lSbfuWGtvU929s7bfLF65TT41K9KrLGmcdo46PEAVbACj7zOetTjlnJV+7mPCnjAsMi
ADJsMPiKW1VCWegiWrSpaneSkXrSSzumBFLKWw3CNFYFMqjgkYQ32BeCe5/GYVAiRgQDs6PSrnUM
ONDbiJtdD0+pDlAZZgFEu+fMkYKdk99jU68ob5BmQWJr9E0FKEPuuQ6gERxrk7F26zgS8OLNnD0D
qzM/ZsTtf5SmK9DoXENRwSokbivUXN2XQXZmIfTVGSeR1tXwPv37AJ/0FcU5aTWpP9C5xW4wrlGN
YkamRn3AqtmTDdiQk918nqeckqeoRh5qB93RHGl+dS7el5Gt29T1gX9ixaAsPuwDM5c6TGBZWvap
C5yuoTyykT3hzCvhNhnuPHoTuRVZQTro4G6/H0umq1e8LdgnVndMSszLjDs/CmCMz0NxdSnmSHHK
r/ydjiLxejuvt1yeF5CSnPe9i4sZjUnEHPrUfhrHhhAjiWbmW/WuGU+oH5bibQoG/92yX4rQPkxa
l/uJh7efQ3u/bwanoFCXJU0lnGDGSUZGJjFyF9+yH7g1wkok5rMju6nfMeJDoJMBfn0crFOvfebg
zwo3aPrLr5f8/TcCFOfHBR3pJW9ZOYGLUSkeLESrUVXwyKOq2/wWW8YjRaBsrohHWaiGPVf42BJB
exGeFWsquWgcPMhJixxc7jDLgWiDBPDg21TNx/N82NifCJADNztIGTRghfG2I6s6EoHDu7InaKmW
XW1RD0gKGcU4ZkPBWry8JkympIpJCqK2hlMqQggXEGHPsHxXEnHBTML1QYK6aq/BH8ERblw9AOCW
EQ80A+QkNWQCVw8qHB6jqiDapA50oUyM7ez7rG2NI82+mBHkaHBK1o1lR9ge4vuBzHaIEp7VIhuV
+Y1XADn3dU0l/KgA95xxQe/ieVPhDiNQoRoGH+PtpaKL8AVtSIuWUfg1dFgSZ/b4BEytIljaillC
amuj5GpxuM84fGrvIYKVDivzbV3sWzfPem+ijVfMNGBK5wA7klBSDgDW6xMoPJPZvnAThcJwTs8X
JrTgxuqZ0AlCE81r0BGLs+k1vICA/YJ8JWUGGhZdWDM/qTC6RpbIzUeWz8Of5aICx08xwtoOz2PH
Xz83vJH4Rm2sLl/DaPLgp57B6YnukOC+h23ApJ4Ggj2c/rcV6i9/kCFbMqM5kM7dqWqFsa6sXXqs
dzE+P7xrmiNY3+0vCx/PvCjPnYHDPXK7Eirwt1/zRsREjdCWGHoe9jQvkUe5N+jvxgWubtpZmqT5
9wlIOvzWPq9SMHeQE06qhicMAylCR3odHleTzEywMe6gKAzIqbSFZnGa6qctzNKYjncRxIynxgIM
C6yrsz5LN9P4FEpLdbfyfjiL+H8Tf7o2znjf7KBwHlko9PsqEjYeUKfUpTUSSpP+FuXDNSRODKnv
neZApykiMphR4XsZ3fP8hGb0JeKCskeQp0z5q0JafFjV6rp/qUM3THxGIRhQGoyHGXqu2SPTS7SP
N6gisJ+BUxHdeCkk0L7iRWPcwpCCWdfse3ke+g9rj0nh3W0TCK58UFQTuCnWERwDrSeoErTn7//T
zkgsApqSuSCDw8U5vVKly46TrI5WgSqKpF+GEx9ffbrIFkcUFgNBdiojsMDL96yMYf8mFbK3zQqk
psqlDPlryQIH2GhE8Up7C/IkAIpjKasGx7F96cT44Jf2r3BfWjtb/CO2Nu6rYp1NqdIeGhCTi7dC
+qrxPYBEBrbRe37UomDHrl/2NcAIOYd+A28mfEc1prXkkNJnUgvIJb6xqW1sZgS+T+L3neTmCPua
DNyabqSBDbsmgbo3OgzNc0EAzv1x7uBYE0/kCLSnOVAYXR86ezqtKwyaLgdyieupYMpNEV36m4JI
KrD4f4tfXoReip5xCD7ufKtzuiFw/UdQubtLJxe3VRqH5hjPtNKDuVoAVeoUJfv3pUPnGyh1xa1C
FIKTR0qEtlWU1I0zREFxlRLriLEJLNo7ySiafPPwwS8T4BkIXO6uTdbm0L46xk8d39uFXznVTX7l
SUJgby8HYYPsaBzhFStGL+5Ntv6mwU9qH1gy3A/kkI5xurzUH3HqD6qlEaa1PTBB5hcvpPYam1o7
CiabIHmSGLRhIjOnt0p93500738IhovgGcHtE20jyfYtqFIQ0far8WlHrgGxBdAOsxbZTqlSmxvd
7Sm2Gk1FpTIA3mW66QiqRmqxAaIzUcZElYaDIWqADpZWBvPykhjgt8mAIz11OT0ftWpbfFlrL0e5
N7SAMBgiefreuQzzpFGb9tQyd1wJev6k4yStfj0SgA0Il6Lt7+vH0WXBVpfoBHae+2FO9G5bE75B
HZY8pIeg9A537/Ab77ocgp0dmmJJwW/wvOXMuzhCxgVSBM2zd+SZpOVmm9oLPngcHuiPKfhXfp4P
LJivl8Jtkp3IviY5a1+uae88JM+djY6WQ9IuQf2+J9/BWZAF4s+TJ4kieci+NO73ScwsTDwdsO8k
r1XoE4y05++Vpixg3EitSCWgMB4EMYs7zzrdvU7WbwP1SigrYoCUW3V+yriPb/YKkFkG4I00ADd9
Eu2v/rjxpinRgntfAzQWEmVhfUUXroJH2OFhA1cie3vWny6iV9Wj4fQ7Sql7XCi8KeQ491jmUzot
vWbO06ba4eXXTVnvGqq9OmIXjmFbr2BuhCCuuqmEyY7pzGUA0jmk9QITJ2kNQ2+vfh38WICoUqVt
ZC5w4JnGfHY8SmrXSIONcXVneoRrzohrtDJ3OgAguvB23mIEtfKCIYQacPRgeCdU+SDTS2CPFxWz
mZuXJgn1BBqsn/koPaBjH1hVJ2RKQRowQooiCTGjZDMfzvFqW70Ho9vvkPwFYr7JImh3nhcOE2mE
GxWPLJ3Y23h83UIMSWrnN0+6B3a45mPaYf71ndJTrR64aegmDOXUoUghPlpv3GFR2XNOrjdtPDoO
pWtd/yLllUWnSX+FsyQVr0z4HN6G9RNHCNPQSFjWOz1JHD03Un7ix/+BkFRYmeeZFT6OYycenEuX
X0bkpru9a/0vB/Yc6chtT8/gmu9TkcrI50dpxWSZhqLOK33ezuwx4ygqFuUhBfQWXoIzP47XIEIb
A5lADDVJvJnwaZN4wXyzQRQHcgVeFr2es8/I8NjNYuW4o+JkRg/rdJOx3/jg2nQBZyJmJAeamr+0
1nsH83DG5IMjfEuq3Sm9sctvQGQkpOOY5tEPwwPuIO3Yn/vn21Xh93Xyor+woMiyfIqA/zj9/k7s
U5zYgIX6k0lO/IjQGx6dArnu3AnaeasgSLwRPhPDaq8tLR8yX9qYizl9bS/f+Wv0o0O1sTByLPNp
MM4iO6zjVDxn50NC+iGw8JIastzd3QFWi8SyMq8P7ZcYhTlQzP0jYzT7Am7oQGHk1a0g0jhJBhSG
pRTkgM2SEpc9l+q6i/kWPzEpLjK071DVsGsXEcx1iCG1pIi/l2THrBPAZKYEnT+CGbkaN4WM4tZ8
8jdDxMbajHPood+zvI9hP8OTc/UCnAZb27ESGIuz6eY1y7rhZsmXgI3QAlAP2e5zyGbp4vaFECcq
/uoVvvVUSxESE1L+7HjiOT6PxhPnzIhHJnl+e5rE9NFc27JpGQSQzfGegLyW7SrK+jZixpq1x9/5
5MlW93/Bq8F2hh/b7doiLdvHxC2hCOjeVD5mFsJMAM62lW0zctOKkZqiPxkmd/8gytzlg0XLxRds
/jjchsmmpavfPlOldmkDymGT6Bx2NCilJ4H/i8H/7u/rElDPWvxMbV6Wv8SJ+PiUbXB5tqGT/ewl
v05WpAfB1D3RQ7OAGHg6+wKiKJ4tumub+ZmfJMOHgX0AIx1wuJnPeqK231eLQ+V1yx+cHP1oHbZE
CX3w1YMNuwu/lpgTjkpsbva5SyilkxT3qfhSEIUCggmuOi8HgOtcHRvfnAtP4b4cCuun1AI8iijd
N/1l/GEx5VV9bXHbLzyHA8a3UD0hln5Da1ocbAqV1/kXCk072EOQ4vtROZPjhLKi1xUYnR+nXRC6
5iu4zZZI7WkNSwmDL/pwPi3pniqX0O48T2BdfrjQkFlgkwvUYkv3ef+40O4T8ROsrbUVsT20vg1t
hxbjkvd39HvpaYOS0A5gCTa/Gwx+m10ioYeUa6D5vsT5xY29/Pk5njYOLNR5mzdDJuJQ/1Rrx5mu
tCI/Pt31sa1+hHShkqm6OA6wOSBzkELkH8low5ziVmG1RsRTLd2UYSx4erVJK+91qS0gV5ZkOsSp
NSYJCAJEkc4qSi7QgePQLIwPO6jlqrg9b+7EDYyPC4SUl+8W0y4zckFHHu2KQhjWTenWWm7J2w4K
7BtWYuKiCoPzh5iXWh43eVD9bXBV60xh7mFNQUaLxaTzAbfREZ8gy+0yrmKwVpPlI7zKyQ6Li72i
30Md4bbxlQjKF2xzLiJeDx0RGGBxHoyan/kijRpf6ygAczJJnvPKyTpQyfdinPx8Oj6g7URsmKGH
3zvlkqQCR19ORRix525hSJ5q9DaZN1tf+LfT3clgeUEUewRLDGc1d1XEzRmEULTQTLUHBaujd1jd
aAy1o3ahPrT6DcNJB9Z93m9XgxyiiWwl7P7HB1WaI25T1d4L8Z9ffh3/+JoTthVzfdabHXAwyGgg
sqfrhCT95vCk6QkWJVpxWsCd6Eorx9nW0YfY4WDIGhcYA5XdFB4oR0iqZDKyjAuEqi2jV6vVqW9G
pSmKTmbjmKqDp6dZV6YdlGXmODh7GOOoeJZiB6iD3dTE4/tV4MpSU9UTGVcwJ3TtcRggdIgYbbaJ
8CAaIMnQJ90u6rD8xFHRtWMGlvwCGrYUniQxhzHHd33LMgEo/Hkk5EccVWAzFkIeRqWPTH24nxjX
GWPWokycV84mvH6OrhyXcEPgFA2rhPVxmsrOQlAg+ail6hGX6eKebnBeg+Tl0UlNgaEEhSg3yGNY
yiOOI3Z3HGj1/3QMNeubkWlwiz61eH5qcqyKrKZobX3SmYIa1pCr4aRzIz70ER3UA7LF+o1/CRN6
rZkvYKruGpQjgaE1dIHME/nFhOzjwzYwXnH9Jqh45u5nROyevneAUZhuknDto/Qzpl51epihdJ5b
6j/kCy9LuAKvrHZDZjasM/QhYdonJhdo/peaM/txBDyHspkI1S13q9J3QeD23fBrKbGqMnwf6Bku
ag1UF8S7gzMV/HIlKkVdsCYH5P6JYKSFa+15vZbs5Qwy+uN1xs91+3OiIcuytFpKH/RoAc4++BRA
wptUGha+I0g8AEZZkOsTzcMenu2fWsBkkZRSwttgzY8UXGLhuyj7AKotfdlmjwBA4d9PPtMwbzHd
UXAHDYgKMYPX0UJSz4PYl0WlDYDC6FUGyAHYkP7GYso242APZreVnWmUbk9wJ/eabeOUqI0gaP5m
PDP0lDRj9lNYl0dgqb5zhgx9qN65kDdITdlEBHuuTnBTJ44nhQFsMqrLAEDsA4VgQtSekfYxSP/w
+zn+f1PKtMYPM2fRSTkwWYil994WGKCyLzYITq3NihfhZc41I+N5COC+UNzUhFxMqYfmK6Rba82M
oVdcMiyErCZsxk+8mGFS1bsnzi/+ZYh4YJdtajguK4kZxPhVeLbMD2wBN3NLByjlKejYh4Vbhu8T
jnUT77Z4JwXIAGJekIl0W4iDg4UoH/6/1r7rukDQ9bsmU7UXNhZ6a7PoL4gRmsFPGfNUrbBe8S0D
DDheTfXfG2xhcvKoO21QdVEOTPrxxGGYlYDnlWt1WE3ZaSS9oOnuBz/+EMIs8Ghng7R+xCODcS3K
vi62Hz/4kstJ3qXX0OHdwpEocv2fsucKeoMfiJdnSFCGw+yQOVkZdm11pUUdTixrvyPkq5aHCK20
kPhRN2aJKxMJwWzvaU21cg2Hnh0p8GepoCys/WJFG1Zbra6UjbNuYoaSIrPZZ6QV5PY2T+9OSuIV
7bPR+D4lyegYb6RY3oqkjqoE32hZw1D/o9epjQLvkwPQY4A+ue7It+OE0Pm5Qade/Ssyd7fKgl5e
6alybEzeye1x2C2eOVI4VCv8RFJ9S83rSaMXZXUpgnln21wlMnkx+Un+YHf9iLhnbIhr7VkTgQEF
zH9IGRi685RNFGn/n3M6WHea/Ug4lMkFN4eOZE6QZssd6Es8erLkcmSCr155pRzoNXwFyYEwpx0p
NXHJj5Pt9WzM/Cfx2ELfn/mseutz0Gq7BWuwquYKQHlrLzkfNpC5fTPtRDiGjCUIqyGnIxMAPbus
qNGRorZJafdKSPmon1NkaBIb3dEp9uuNPXBbefGLWqUVwHygHquww4GG/A9X2QdRfeWtI0xAucCO
Ws1RtJ4N8iKyUY1il3uB/YOM1mJmi3PfI/UZM//jSovBRpcI9/C3cFPnJfQWSaKnLdDgBvrHvl6p
0wmR7k4kXG9nLDTKYXVpYUy180OvJcHoxmC7DpF501KSy4o7TpDD/cneI+nu1mbJ5ftERCkg4pvM
rPBqCIuX1rrlEnR1yn7P43inm+877vVNbDQ5ZAdvECgQDt8GdORfTMSUHxd2BFcq0oW6JKMOGVr6
1OIX0ZjEpGUs8hKUPWFKHGvWvrb2tdhZrOpnWHiYTpZWv5BdV3LRmZZNb5YQmYHM2IJKeSvPEtU2
R15WRmwB6bdy6ZyAaJSpLICCdbXPTTLVb2FW2Kxw20D7f+YjhFjEdcE4TgIU6nu9NSemJjZ0T19o
5fYcI8foae7r3z4Zj7yyHPxRDrTgJNMst14bw1/lhpDrCXlrg39/Gw4gFBQI7f21cjKvH4853xu1
UlTYwCZfsZBDI6sBW2tZ8yGIG7q+AWcpSSh5DaL81QZm06ho3m1xak4MGr4eTttCQi8+wMK1NTN5
yKYtAuINBPsMVv4JlIaltFQoQcuxtpNxqUXMhmhbPQVPLsWa0zQBI+f1AoOEbUGmqs56dGHM12Hf
q74lTZTbMlWyOoaLsIv/b8dQUEL1EA5vg4ibV++qM1qVMlpSXYv9XNTnNop/g9hrRkILLJwyUlyq
n7jpHj3qHISkZXpJJB5z6qsy0YLjPzjOPVNwDXzrm22+IDe5a/52nJcTW7kn/yWVXjse//f03zKU
G/vYm9zmrwyBL7eAQjBiD3Cno1O2vN61IKdO4sqkLr91B9qfSlOhiN9A+u9yqJgJg1Ltz/soqtmB
1hsHydmT6EKjt8MtXtu08SYnrQ9WusNkxojBvaMmSHdiErs23JCG+jpHFfALVGAaAVb1OqeNxcmk
gE4GKNcV2Wl+FrbnJxUyvu3KXEBpQ5ZlEad/W61FgJSLI/7S8GKiAeDBEh4YE5z4OMr2PfIbPuPb
U0Tyunly3+z21PzG0amQOsEhJdYQZQAvPpJtZCMZifAZC8DoOrQ0AjDvgcc8BxXch+tFdQkXSr6F
r0xFatxbv0Tg1N9QcG1A2Z9JW3JwtfzCuShtwCfFacelrt7MPmNclO88ECFVp9xSPuqJ9yx7gFIx
VdkRo9vIn4cdSZm/4BVcZfRsQW3jKzpf/ux4PzG03Ye0sVss5KP41WGYWywHZ0fxiKipCbxjpPhp
JpdLIhwiMoLvIRR5aNlqljE2kPyVm0HNfNFIaNKfcm/wpUFSMGIWUiqfFz/j+O0ErMDudADZUz/A
0AjoaNgYiZBmHnhXPpvrN60KZSUtkW3/Fpuis17uGBcnpFtRaySofDvahnGZlA/zG03Sa1KfdCHX
+t04kxiEmDKRysyhfAYaHz5PYMrslxsgoR0JBUJD0ZXFff7UAk9CLP7QB0mFI0U6H+J2ddJUSGIZ
hpYcRYAt/kkbsI+zqv8sQonYBECRKGXCGYn5ZsHzS6tfr4TVOJrSZLoYkHAjTzrleX8H1XhJSnEn
5yfH8/CdMQ8wihT2JTpPoifcVT74xgcxDHiui99kDfi4n/6aXxOLgKH5jbvIVQyzITtcYqErgODi
w3nQ8RPmk92tAuPQb+7JtvGSFJu4QCndXqqibVw5mo4ArZe7Zsx5H5zrB3xQoqbE7gvY7AwVzFay
/7Rn5R55rWE7NKbmJQ6fXuTMWuCxdnro2aR0eP5kqPGo0iamOKiUoKu0EaiR0C9GPlx688onlyIg
Sm50s0p3eePGgZYpGDddp+yVtkaGN9hy93C51siEC675kkb887tEd4ljw7FF+8EbCm1jNeuNi5yT
W0wlFJXi9GrfnuZm6kqaD2o9chanv3Qy5J4QDzSt5rTf0imk5sUmjLCohwwlDTYoaEyihu6TlZQ1
7mIVtgzsXyxmyh7BTgAM7ve5HiXtIaSbg9sXmjYMO5HwL2nuDg8V9i2s6FIGkW78oJlUJQ8iUjdw
M9DmlG0d8rW4coSs/TA+zoMVQNhVyCljyp2yHn/a4N1zU34yjMVW6uxtkD4lNy2AUxlquVuENOz6
GHZap48SuqCzFIxR2/fiAAD+ldNqt0TBbOImhLHg54ZIIxNVQu3WuXzqHPP2zxtgJZDXkRWf4LEs
jqnib7/iEluU3Z8+R8jjBfXRgXQhXjmvfF6EOcDNOXzQfB0Mjj1IWurBkUGN4V95Ai1cqgVCStBZ
SgKQiKszPLcqAlPiLfv9XfIZ8iTuUmxxRwx2z0rDFGumapOsH14fHEMaLFxk6VXZE4sTsDN7zGUa
aC6UVjWcwRLeRwQPmM+28XTysL4JbMtnbzAGG3wCzD0KHQ22KpEPK8AHwGrJw9Ypuqi8bw63spai
yhlCd743la+R0FrVAY5A47xvrfVgix4I8R6zZ8L/ztqkEP3PUF0ObdU0QeMvaZtBtRNDMV8rLgwf
3W9LUf0GbM+O6zlMUgzaxB4yCBg3sTRFhKyu291MAlsliGqPFL9gRcvgj5wYorDjuwRXEIMvvYRc
s08ba2OoEGOo27/Ve9abIEJNk3riySV44L6mc/PwjzYdGpEMvaTCiuXorrv5m1RlErjWmQ/OfcOU
+DPH1Sgis4SToehOQ+UFa4gJAXqLo2+UB78QvWbykDWxrQj2VnCMG0+Ezh4CHAYYl8LpcFs9HFiF
131EgmjAmSTR/SrPa3NIooMDPy33Swsu+BP5uaNSCCmD+qJ3/ug11fIDoB70XJ8/Qi8xDo7iknjc
wtRPRpS1M6Ts33t+Gj78PTO6iMZTzPEZjbDri3j/vygZdotdiQTdsgLhvCpn+TY6K+i2s/3rGOQy
j0Ch0D7SA6PS+Lss3aggQ+tRFWr27w1zHaww5NfabzjanxPYi5A6ArmDUVFnnIrMcaz9enD8X2nE
phKi1k5qOITYigeZ5ub1EH2ECrWt3twb9Y8v3KU+cxkcWrFLjO7R0JGtnLu65fbr/cyyCmeT41qJ
pZfdSth96nQ+/Aumy84RKlKaKhfYbImUeVH+gNoQ4l/lFAqUL1uEm6O3d2dMfepN3sPN8wPQpG75
VQrsXOvfatxBtRD5gwiVwTnWtefc29dTi9uUSjf0h3Ze2KgG6Bv28zpECwUhVTB2EDXYQwyPKBZ2
zj2QB8oZwTnbbG8A+O2OvHDHWUEzEGHbCJcHKVVnxYSNiEjs3hY+zkgYnf+y5KQl5LkSbM6/ZJuh
Ayp29IHw/wXUQqprnscg2New2Z2sCtnDlxepbF5U9akIsvtYRz+jm/TYs+veOvB+A7668Wc4/r85
ENmaMo19yrp/5qVm0VFVyJASdQb/USd1q2TyzdWTkBwLEJa4FIsUOh4tTgGcrM6sb9fCIFa+NWwl
Hlq9rTrC12xg0XUhTUVyhwkMyuECjZOPn7sj8Uo/2sH9tkcX6fhfWIzcvqBP/pQAmRS16QOIQ2Sg
7PRAZqc2yvtBhsVL+6ZjmO4rpcSQb9U7YBS3cbIhbgmGNdYDXdW884pnKbZOqpBkSDLaHxHFAxLh
1R9zqimFS3JTvNiM+mrG8g84M6Ma+n+xLy9e4kDbMjl+6n67l8sdLUIW9VMB3r0AgSf0Vh0L7P7k
/7bb590BmE3VYr3yIuilaEycL1BZU+3Ed61Urm3RljfaLMiRpoKFY69FeAwlMjrIr7OXVXeXwQRW
xYR6SR1ZsEthgV9YDhQQNWwP6JlWkEZwU5ESsn9707C2F52wao//JuQQY91TleYKL6LDEuF1eyPO
VwISN4JQjUyLkTJgv0FLBsnSzTAaSeETLc2+Jd9FtS/+DHttZJZZAEV2wN+BK3sYNHpKoDO259jC
rbMiSbudUfR7dXWjPDJ0CsSlG0IKxuiEmpqAj7o9FhfL5WcmpHlZfaXTTKq57i8X1XBxlCgojgMP
sOPkyN1ctV0VotAtdHEydt5G25QftHUqj6N+zd+hydQWizrxAldGQSIn9klsvAms+MHy3wbBTAtC
r22Jr1h3mGLsCqpStngyqL7yzyxaIYEA24gaxqdvGKwME4UATzTIAjQ5Kwp4sGFV0mebuq+dHofg
jFDXzEyVoXkVbBRQNieSC92qAp2FxZeKWybtSrDclpJ76W5Rs1JtU1EicLw3zlttxfyAroHAvQNw
V4ksNHcxAbG05aw8TR89ACfcv0LK/jhl/4VQFNkgbb5X/8xCv3XUMjI2Sy42UQU+zXt9r9rl8obx
D6sWt15uOUzeZ0TwWCKJ377SPgdxr+msr26s4ampZP7Bnua8ppv3HzMxE2hlzy12iFRKk5QFrZeN
PcsSQtOCuwlW/V/IG2UAux1zV1tApDN2paiHs1LnA2H3bNOMXc2ZcFuiZ2HJWvnkQ95c+gj8kH/h
hr8R6z/1RzzoiKxbnY11gZ3eUHOMMYYDpuk22b/Mx4rOZfXw887vl5quaR4qB3gGmMo2o6J0PBXd
Gmu4EMvs21Ynh+TggfYCObuBT3VKHkj76gV18Ip/iqYoieymRwnCsP6skRH27l/+iLvQI2M9WRUX
SGtKr1TZ+n3T9HKl39xwmyxo2XEAEz0jEsqM3gkQoLDlgosk/vDT+2NudyZdMIe0A5436enVFr7o
lwYlCwIUjLa/dESkpuL9LU67sqjineCcdg8/IFy+te33+aFSHid/WBK1kGIInOXjtWieCdZ8kmQs
3stxWqwlhXWMcCrc7JZ8J6sSRhO5bOU+JYU4t7bG4E1Y9Es8+SbJKcmgloaDtTGdSgEBvCuZOKBa
OkKxxpQpAvWDbQ2/mkpqfJFiWmn2r+Ko8v8wXjB+PRcMjmN6/LWd+FUTyGR57YX/URisEgfKbWlV
BljnByTfg6WShd95uZvoUQ8EgXjRBgTJg/LdyHTyZNBq4LDtqeWKaHEZ7gQ/SQwJvqN+hRKMNDwm
4ZrjxNr8ZlOkRwwP5z+Hxa1w5Sv8zpp8q8K5IfJAFvWpaF/zT3Wh00sN08HMu6sGYsqPGAchziQy
vxkGlFYGte97uwj5afq3gGygdWl6KNqhh3mRqaHEw92f1FctEmYrcdBtCQ97rftb6lEKfYI9ovXb
UUcxgJgtCCn2QCze6xEiMT88LbHpWPFzA8YsaRzd/Xysowm7Kj3tqYWftD3GWIfw9iA4/YZBG+vY
p91KXGFBbRPHXs4vMJ8K7mgSGR+3GMWJk563kWhbURWVEQcYJ3DV0mept8q3GNjkTuE9nlxz9rmS
WNS1s1CfpGE7u7q6cj3mxcgAisYK47HuICo19px/V54myggW40E0xN0o7V8bfAhDRGSUTaJVuHkR
ULf6v/WAgzEQ3hcspEVNQ1dMOg72lhK6HsOy1aQnkey+5y/vaXYHM7sAxGB37SZpg9ufKjzIvub3
BVwHrZQl7w6FfQIKIXpb8PM1uB0ff80p/jNZ2u2MEAnueVsdkea9KlXt1P0zIaBo7v9aNAeiocJq
HeJoaaboMJzFtpWFtjnBgEWcnNuBszd2IuhAAN2SwRyKeJyDfkWWOWdwQg2IqqrzTHS+yMvfhG4W
f+5s+BDyqcH3+0YeNKEVFU4mqA2NCFl/Gc5QS/97FrXtuR66QSXRW/ROyuO6VsMspsDO+yRiJr92
mFICDdZkFW0xiuRriFkDmpBA6+CDqC0tjgU3B83bb8EWcRX/qX0ZqY0/N4QWNHjrDeRB1ETBAc7M
bBKrvk4o7Z+cewjFxAi6HeLp8Oms/6uT89Fq0t4xJXQivgcSChmb1VlHRqdqGIIgGDamr2r9j0WU
sm1CnZgdi+CwCcgrExHt5wAxuNwc4yv38pRVW3fpeoKN5LDfpLdiW0fhDGGw5X7cZF7tSIfmQ6PQ
k2ZryLTwNHh/IQVCjreK9pjpx98iMxEUQ4ky85Q51R00wXm/hkiQIZn95ZE8Ld0ykIo0mC4DJuNz
3IseieyU/h/F2e6s3OkbiDWtMLo0HvCAUcGx/xpRWrRC8/EvhihA7oGIv0gwvWL7PahpjdVRUMOy
EGb2Pnxqlq5k1bOfGjLlWHbtoREWSTNMRv5poTGNgz28qXymKoPwps/aTagIJRjCuJrE1w77n9gM
Uyxq013VN1Q9PyUKEFK4GeP10tdGeqyX/bgSTrQ5NfR15AfO8jbnd0LCa9aSNa6OIE51Guu2G8QL
CLS1GW2DqWdS2oHZiwwB4vPQ0TmW+G9cKDHDimODHqt3rGYZy1kz81BohBG0w6qYYFqgyb0zXtDm
4BeEJ8F6ukXmijUFJwqZ0jGI53oinK5nEmNLGW3AUmnniGhhNRxY8rNHvciNJdV/M5NAgRcf7YhG
7ZVHRlUFAR4JECNwvLgpDOgjLvqCZJHrOY9h6ZePANQqILGHg4eTM00zZgUcD45duwApKY6xSKNp
zsY06C88QFPxS0MlOwcOmsrGfLpfw8bOtLoG7sdY/WcZjWsGE0h2v1FLa3+QkgA1FLel+k0sWjXt
yJTAgU7qOdIjvOL9YfVh3M4M36KfUcP3/xSxy49HUpk1aCVyA5WMAGM1SLhKiAyltjSJP/9gbTcO
TsW/HoLT+Juetcufg1Oux5xxwigjiaep/Abqj57sMiz/R0bglIpveY0vC4M43fh2Oqx7SmHn7Tvo
q6LZgwFif88L/btfh60a/q7PFYhpHFL9ZPTNBPN2ad+CWoIH0ui5P17LUBwihCdFe6sr0UigZXjx
2De+Mg8XYPjCkYtExCUKT6mbLMvb3l8ishW6oC8dvYOm8AAho/2F5Jk14kii1spiuVYMeSkYaSgl
th22TUYqnpzzo5LKbYgQv52kWuIV2mN10jlrOu+z0SALCPaNmZLwal7xtLBcx5T2DEeeGYGlAyIj
ZjUMZ5EtcFtRITqXgt7NNuNOXxXbfq4kM+Gb09nWP0xN99j1xFbE2v3pvQIylTCaRXaUKu7z8xmz
+jU8Gs4Cd/bkd6Qc9vqmJRJwOPTtkxBeSh41/HcRdyvQleSUXno5yvAASBog2J/V/Pa6TdD77tS6
tRRV3icgnbEWXPiuLQ/xpWkeFsJXFGIkUsvxzJglc+vs2n2k/fQ23JuRjOitpGPuUw/GnoQMS0Fa
Of7hHWuwz0bvBOJ2JHGg1CDA5ONKKQq1r+jXEKkvwmrh2gAcwpTRdaUJ2TdCK1cUKWdAAZl6MWWD
6vI0Wiq3aWevLmoqN2w+udzTt9RtJvb2etRexZQ8szFZkIwQy1QdRfoVwb97GWJZIYNkCOVOA12T
WkWsxyqlaRn5rmEZBCBGq+Zbl7d9q6s5S7hbpmXLbM87p758WLmwwXIBVRtNV1IVpFY8ebPUwl0A
bCdzKjUJGNkuUgwxYio7KpE3ZkVQwo/gBRn3ZlVpv5CC2lC+bHR2TIF+kR1SM9wJtPbyQtRg4AnU
XxsaiG+q4NIGVcuEd45KqDiR9V5MgC/NxSr4/wAg6m1yd3grrCtIht8s7aU9PT9UsEo1Ro1Z+M9o
wScdFiKGh1jgPZmN4ogRrGYXrrjBMOShgQq1mEXAajTTDn3BN8ec3eCbSHC0pX5KSYya+R74CDMz
4Y3tdd1GlPJSh4wIeS4o5w5T6Qa1btEt76EN64+aZq2RVjMDuTFMmlwh1jpPUBjQR8QixTU1ac12
eaejkFT2Kp9gbSIo5NmI5R/0nRsv/UoRNA3j26qV7/oRb1laawvO9G6ac6jCaQbNqwZ48T67tos1
cMi2E8X8991wfv+RkqQnPBoDrIceUj2KGJNbt6aOEVTjFdny8zE5BUNayEFjXq+qtiR/L4nHUAvt
mIQF828AwO3Ev4F8+mNCLjEPfPNmD05+MFALY2drt86iHJLSec0NUT8yEGZqLu+kKj8NThcWkCb1
vpQKfkjbpogME8VaqRvKpHQoD7xm0dBQUj9S5H7r/1JUwfQMw1WEab1UxD14IhYDfXknXCzGPywG
GyCpBYdQogEqijoJ/+Na0Q/imHylsFgMLWzoN29F/QEngbCnECZksyucsdnbvli/PCXpY4jFYtNw
JORF0KdWFyBcEMQPLmBBYHOWD+k2hFsrkbLiNik0tUQR3a07Ub87tu5Z7lx5OrA1OdVa7e7vaYa6
6xj2KehtUJ3+Eosi6nPXmAvFd2sRI1freV8O2Z5oGfEv6FBlsFL4MjULHGAmM6/Y5cmx0aDlmJwM
0+/l0ptdU0AZqBUELuCbVfOCX9rTDT/9cNJzTS0JPaTgFGF1zQVgV9/VcuzhMW7hzfZcqXMUGqf5
AioXWQq685WuXoc+MDghgpZ9JT0qEWRzTZCsMXN3RUa+BM7/Jrg53zJBYZzvkCMYIQj3ANmjf4Mj
G26TmO/gxW3rkiHs43h+8kwimys0zJjarQQivRI9OOHEenQbcZDZrf3yuNXvZxz640o+1F0um36P
bsUfd4q9reUp1254RRkC8lPU55DQp1bg+1l4UJYSU8amgLJfPbQcyzzL4fL5p4UeOpn0F67Y7oA+
voNVdgErBo1j/Ly5Sb8p7c9MDccM/tNwy/cTIPb0MQwzdqo8AxcPx1sryPKC4bqLQEESUiatecG4
rY6txdgPqh6Jz50VURSLbt0VGp2DV0lMmT0+uwH76A6JYrjEWNJzzEPumRzCiNN/HYksvKZ/o5XW
WufUBpu30gs7sH37CmzV6wfu0qX+WOjks78VPP73xPAfDMKInoqLSVaKsqCIj4JbaSgVsS58nWD0
PDT3LO8sbnffPNRQIuAl7W3Mx15JWVvQ113SnNalyD8v0EbGAkK3xmSspdh2ENajjGANppKYHjRP
Rp3lvUdOPeBORue9LeyWcuhfajhS0jdoXBD5W2Zy6puOgruSzC4zb1wk0lGUs+uIJTrEhlBhWxnm
lfBvRjo2jdsjatJZ3rK+Tv9GrBER2l1n8F+pm9cY8s6VI4xKM9phzVqSxcqd8DixmTr8w9scl19m
/Mnwd/UC545J68ivKT4bgn8ghdXGLkZSYcnewOTcBEp7prgsw7YOE5TVS+zMRTyLXDglfNKESZrb
6NMIwW0H8j3HB/k/6QowZ1VweE5zXnXI+UA4FEzA0dgsgLcimNep4KUjwzVoD7kHort+w/jxQS9F
n7H1rpDbe7GfjMu3TTMMzFFBalgELG6J8gPywqhXAdohd5Oau1bkRbf/W9gY2qtLElErcvk07frj
4p7IsDzY6GyhfL1N3vyPluswDbAD0TEENvCyaux6+7zK2l/6NB4qOIqE32CU0bu8gm+3DG+1+qFO
f7evf2rjPJEkV5Lv7wVY3N1biofJE4F71RNYZS4CAGrIAah6h68Vv1l5/r8lku6LYmnEkvI6Yjn6
lFiSGPyWcVG67sYaKDizrJFz/lAH3cxut5+P07PowZeAJHAZ3yHQqy0hILn2kC2jur2a5GXnoGuq
AH2BN026Rk/5HCEwZ/xXe+7SaAK39lx7zH57nzOtW0v1KKI485qED7uNJA4hZ9O4morNTjFlKiUI
S8WixjtoXuAfWY85k9+0M+zWMSCd/3b/vipd5+Fx+yNasBAqQm1VWtsyuKBqBajQxU+OYhRkKsQk
j7CQGNT8MooF53jvdeltVKIonR579IhlTK5xTaQot1M1qyNvPvLwF4tLDMqPMlVngo8wSBbS1WRh
ZIWdc+zJgKzmyIqujNoWuIY6qG6YlkynyQe+kOzKkYgsvWuvqiimYjmjL0qq10/OYjBINePuElYQ
Oypn3QmdjtbU51+5fzuKWfHS4O7YsvnKCj4XWMPhNY8ZWO3p9GPMTgrjr+gjR26vbuvZsMN7lNqX
wlwshWtrpDBdZUtdOR7ADHdldqQ+3gKpohswlPCOM9ehulRGzAr720SfVMinMXk8r50CUiTSGL1e
6oUIO73XUaNBxouGI0o2XQHEBRuSsQjblvt2XkqlO0OJXtQqGq10wjRNBP9l05m7Jfbi1KQu6HwU
0tboGH/qW5j9uTJ7xaIMlkDs63toMki3Var66EHJsVSdikvH9/2W+C01zD233u8TpivJH6yRL4SK
pdRbPKsoyurWdgKaYtRQudVGw1FPBpCM0NlOo51SsNzZla+utVtLb8b3SC3F/sPPOvQUp7fBm7Im
5CYXEcZTNDE0A9Y8jFF8SlSTIVpRDwLSqzDvPKN9u6GnhUCxeQHASG2z6cPSvLd8qLXDSsrmdzEz
09U1yAqwsukUkKUPccAfUs/DL4R8rXqx3tdKOqBiEGJj9jv+bMJZzEMo6syWWu0QIWn3Lf/kf9fR
jb7GTCIGnDEP4bANJgy9QG0QHytRy0rFi0OXU/aWQNBY4PBGQoM8YzIVGyLotdRV9qsk64geUk6p
TxlGAhr7kFIMfeZm5BE2F8AvvtKGFdGdiklJLd31LhxDSbBtxyIbV3iFOY4XyZ3SmDG1OV6J5nAV
vjnps0EBuMYPzuna/d+XJRSo17ee2TMC9NsOrxSsOC72d066EWw3/d4CzPdDoBgvWsAODlbic2qa
8Vzfs/4AieAiFtbcVBZNVH1uGAP5vhUzVJoRBzyl5MhwnS6i5WqgCm1CrYCMi8dQx1SK1aSjlcJu
LK8xK9PhHuTnAOOaFdcZ0tp/c2PLUpnTTml3t8PQVToHf9zMPt8fvAGFuikCNb61ZTpJE+LU7XrQ
NIGkiK88ivkKoRgmwMyxmswHSPSH1hAZDjjCGI6bE/EoqFistimQNO2aDJAor16GFDV8OT17Jj72
jM7XNV0r4Shf/rxnL5iCdD1etlRnSoBVm6U8gGmQpH9owd7bU+3Vec5xGDM0JP5Ku0VZaXlec9Kp
8N9MUEP9xCdW3Mh3zLrHu4s/6u7KzjnZKMAGNb8M/JjfK9bK2jC5nxE5JepZtij1rioVEOCEPz42
ydGRvSL5BO53J2zPxA5N9uVWpp5DTYhyJRQHvN+nmzRH+ibBJ1PheX/3v9baOiec2q4Hau+NC1IG
t/bMgIufylj62hW536fwSGhN1DyZIuYuvEM7Zy1J8GUE+84ootDhBQXTHIGGa09Qv1u/F6X33Lz+
4Ey33yP8IU5eVNkqDbGaCvae6EZJ/0kAspmZL24w3HK0Z2I0oTOdZ73jES01F8hgSZcwnVCj3bFL
zfTo+m7b3+wPopNBtHSPiLTAFESoCn+gtxarj4O6e8NuVQ768RGAYzFUBlDaGGkL9csGFbSa3vLG
TIUKjOfGC2YUWQCm+62hoB/gb0b5MhQP60EIs6pJdirVwR7yfnAtZW+EQ1knkLztHuppPmrIV9SF
beR3ot8gMxoXolBwAYgZ0q75WO5nzDRbcBJuPrFE0ezPVuLEnUjvxncQ63HmO9tNZ7Q9Vv6693Jl
WEyYqqBifz6qZN0puwIeCAqN8j7jWcHeJPPKR0P3Fpy5zCq/Vv2ZF8JY/miQcSEccYz0G6hRKN+R
VrLF9bQCJMkJiWmwyM0v4FEvoWZJXGWC6Nfm32o6662OcQ0Y0LJuVEX0GafwoIkAfSxNYMtW+iL9
w5xQAO63G9dJaPeLNs033HcfdnIetz9nIDJosh17pTMyy4q3Wr78o/rrZRIY4lrPbZzRAaHNAQBb
cHGA83DSxim+GmFw4joj5oM8R6K8Uv+Z5cHxsl05Hv51QMELE+hAGQZ6P50mJVuE3kJUrpDZNqYy
PhTOJn8ceSZQjAeXbtYNLWfHhIuS4TTvoGEEVfMUX3+vLUAjNiqqQzV6+E1EBq53vaFLTZGnAsr2
MORTfC2JcFM0c7hll6hrpPmqmcDF8dwJAJkKRhBnlk19Fx9atG9IcxBRN8A/T0E9++TZp3oH5ylj
l9R6TrPiY96Ewjbb9j7OxoQvpkBoEJCrIMK6yazqET9VROoSHIAcj8rFyNeMRyLngXS05HJMGseF
7FxEq5G2PUXOv+XMw7kUO2Q5WMToYZZoVGbKWaPyQWFgXtfDkE9E4nujHFJGf9A82F5FICMJsbZE
/pUZcrZdF5h/igwBGVh2al4pI2/sreiAGoMKNPIxxf3cyzc2Z5vt987w79vO6iMd3Qgne3tbepMk
pEb7f/js78cdPZDY80TtuY5ACmnCPi7mWXvS2UWrFAw0Wx0euhU/bNAujp92yZDbqbizQyhonk76
Vluonb0p4asDD3NAdyD/NaoRee0ZrOr1I5bsudAyQequhAhZ6VBtezDncc80MeGRFVeCSWWQFWWr
tncgppIFEB6ZiSsQINHcPYe/l/SylMZ/yl7i0cFmOiBx4xK9sioG7BrrwZj/kxNVNENlIXDido9W
bkD2VVCiPvfTaFH9yDNkCj25o4JPLywjtfqQuwkY9ySwdDeA6EUdDhfEKFz9TdPPrTtD41zguFLI
sq7tziEVZP4/NRFSumrDxcacBJ0vi5nTUwC5m7d/C+QIVBvscruHbsYfJ5dkJTyEO1KSspyfw/qr
nW/hPzA4FBFC8dRaFM98ny9nmj61h5ZkAXB/LcYP6R6IdvKy4V03lrypt5LqCZLF5cXoUePTFHtV
EY6ylh1kpcg7IA4RSUSmKY8G0WNjo3FcvaF/TSN+vaM70y1r4Xp8Ao4UToL85diVIv8M79rJP61L
xr9GBxilhVYIQIkFqrQFErcNNZ1crfOxaY4ODaXb9DIkwH7E/NzjUV1ecEz3vFdbDgu4iD9g9RKa
IHz9qGve0xSeAoipVzPr+FEJ/b2n6QaMpD8lLamSrlfjg2c43V98H8cBu4ksb//NZg5A5fo5TzyM
k7gDJNTbO10JOZ5KFWRh2AVt45R2j8Uis3e8DSurw127NJHpT7vrqWfrQfGqsrmq0HMfqbAAHd3H
BJHffbUDDDUJJy4rgWJhjgc7x/kW4T/iWTfKFW7sCZndwgVxqLIqsKS7QEwd86KIbR+ADKQcZBDc
qhPNAmfS8Y56TlDTXlHi4VpkEghLSvpUOhSFge5c3lfhMZbgdbnB4E8OJyxcC9uzBEyY7tW/uv2Q
34gD56Dm8O/QA5uoPZ8V3lErA4OwJAxmLF7d1h1kcjLb+SOVecMKsAO9hVmKWzcex/hQodsvq01S
E2W5lCrvVpzKk5I1qhQCgdNnCS/DcAcNxT2o4ZpWVseucAqjXgB5EXpSt6a38busvIZmnTv4/o83
f0U1LUtnauTh8Qi8QvZ1a83avOzJvSjLOU79CYEQpHI9swQkbDpRdHaYGEiRn+3oCjY7q2JVlaUi
PohLm/WtWHBf0kexQSsO1DEPWcMzSFtTsvdgKovV/XtAsLEcUbpLDoNvlW7x5PNZB1gl8QfUzCiu
Wh5aTQBGLRdRirinZcyGPydmBuxnh1qADI83sfItCBX8DTeRYUxSvP/gJdJ51QDA3/6V2RoizSlM
S1YphvylS2EMoG5ZyOPRA2OWyNAADdzoM+RpCjV/VzDT6iBZkX5Lbiyli3l7XgR1S2fFp6Q7VKFs
sfiyklFmLZeya4VH4oG99c7tI7Hib6RVOWNBB1y91MWSFkGPqsR1s88oZVr6L9Jugz4rrpRObC4Z
x9PByTJOl9EQr8TAaHWYquImxndQqG/VA5nFixWqgRvvFNvgeFTzCo7z36yoWDWGHvnEOlcy4/sO
JS3aFUShDwzajMf02u77FnYyZ4vaBqLa/uBp/+uwQmdGgTuomo8Kt4oWqMSVegzp0lkmMuvdi+yY
HJMQK7eew9BNuiIJdM0TSCTYiBKf/8wFIloKGvFzycO6o3snc97+nIkBSdareJbSCz+u66j+Rswh
9yjQjajMQt0T8vp+pTGRCKcab8fCZRZeCO/K7cs5N19rD4l8scJ3q9216IIoLKueK/JXDQNUNj6a
gRAh7bSeUCPrrS+ItR7PeYz5FO2UkbSjBg8s0tqxvs/iaE2QY20zTqtPBbS9OA/B9brTiDpFE9l6
OCoki6+Rb4dZF4YWXyr1HV5airxO1H+XeNJrfdK8Irzq6w24nsnhaYxAoT0YyTxXgYLd5kdPEIqb
D8NtCpvbx9scb6t+EuykYahMIFk0brXE34lUbzi2o4V/mZgamnteO11kTMG31y49l7oenI0rcpki
lKr2HUe5mDzwNKO021wRVgdyWz5dddjN8InLQBwPmVqzvIzVtkzCWHw2b6fIQHADLFv0vgnMRBk1
B2Geay4soDpoB523MiJnLfuMZaCft40euvbSpyo2T0/fLI9mly3dXaouEkEVpIIhqAyEbAr2s8ru
uFhmhKfMzy6mHbtDqhBj6/1/V39K0nWhJrS+JZRg9FV0MZHXcFF/Z2XevVUxhQkr8hZEQEbWPe0t
vskE5gL9Uo/LduFLhegQNPJvKUeCXrhQB73X0I9omMH5FVO7nWzUcS6kZD/Fx1k9JdcZvwCMgF+x
AqdqWtPXu5RI6A51cYUJy7ocjly8Mp3j011rGrQRvnKpKwES9DLKyGxzHtVlws/ul4HQGLqFag5I
LfgJHPhrjGC/yZoc4X/kNsdiOLHra0iv3HDZm3DpsABEv+1c3b7g9vdR5pE8xoZsrV+1EJlsNLUT
H9+6CdZ8Ju88TaTHYgvP3LAKcC7ubbArhDucYWf20mYH1nrBZ5NWWqmC66ueJPG+LCht6ZOX0enE
VwxQqITtJDrcXv4r+QtrzFs8zajID89to0LjaunJGMYWCbBQHaPvQbMiYYcdP3gIUjo+rXnHUw38
LaurKwbuy5qfVCbMmu/tyd6WPbD7xo+jlAcRz/Xpmt4JiPkUt8AMCPpjDjuCQ7D5EdGXsD/hOt8l
csItgShkWKr3Du5T6aMm0WZuq0KXenNvmTGvGR2PxYklLlHg5rhnsJYDsOjX6M1f2p1d55Hl2ItH
LMcTtu6zbmSyU8VgrMXmhpRxca/ZzKAK2G6QZ/dDVWu0r9Enbwt80Yc7prilTCgBoqZFQNeyUeKB
ZxZURv9+Dx4+konnMhbimH99s4J17otk2/dz2OTE/WgR4V0XqugY6h16rY7bd32l2obrlyPILLw9
JkQzUKoBY9iiruJ6O9i5dZPCJe5Juspizfr5yTQdx7sp+EuPo2PmCV+KI4oQKKDu9MlOGeLqL8Ol
8JQmwjQ8i7kfohsAogPuy0wGmSWqi1re+C13EbktYWUJfPfbZ0WJyvbYBwUS2+UKG7/yfkAjkD45
7LKi5LpTTT5+ZuB6Xe9vVVPOtOgODDE2ldQvbU0p2I9qkRtt6WyoB4rRlDN+55PLeb7qcI73W7cx
XiaU+hlpIlW4qNBJ58wyhyPc2WgMX+zQ/tQeJ16znDLFTJ93UKBGcfRHE0jUisEsdx07mRg8gRFW
mKjRnPoY47PxdY5HDp9xfpr+L77wKhVM3VdTd7n0tu/cd20HNkgVENMJLmDqPUk25BbSoirfd081
F8LXAczzIsmEWRmMXzKXYp31crKN5SLX9nlDW+F4yF7UI1BFk04Z+y2VLSnW3d+9oojbN8Nfx7qD
g2YbbgaLQXVaUDfoIgO+sMEo3N24NGwoU2gc9w/2XKrUU1ExAwmaC236NHnesQA24+dwxpPg2tMW
+MN56i+mXpKbKk7O25ZVAMfnXfH/KcQVZBgT+wW8MvKWS9I6wNiwOR71rbKcV2OA3rkfPc/5Yu01
cxHMGOb0vIB//Oof2TRgO77KSz77IyPFQkpioQcrI2/VdV/+Esp2BVj6TZ+B+431mLL27fvVhyNM
SoSPP/R7lrX7Go/ZYksERfWatpeT9Tz5T9y1mWusuj9TY0ItRz2POViQrH3abQjsfdDlAX8xsX+d
9whQ+gg5jU1Ku0djsxLXS46R5pa9NtUt1ShA1W/xW+n52l4MOOn58RkQZAFArID/xi5RerUnS4/Y
Uqhp+qYpYRUo4STAOhM5szR35tgWcHLe8i6Ws6NQlnop/w0LfSBtNz4CuDIZyp4sBQ8S77JNHq7V
mnBuJ5/zu3EnDFLJCeZ4VC1ZdknbBV2Z7pxRroRog3I46QVRN5tP0tjiL7hfBqF4xvtNixWsTi8J
BDzS3kvv71CzINr2ZQwGQc57KqqR4jxuy4V7JKBtfZ+P6lXQIAfDA3mxITBrSNVqkYJsLnV3LyK9
HBz5dwfC1lf08ZuOJ0ypLfZlCaRM7BekfeTnCSvg42Z1wdWpIXToKMOIYaOU2S1ctavMjbh/+S+3
xmHVZZSJfIJ3Yr+e0vawxVKw8ghlZ5Ler8g/LsXmDzV7mIat4dxNvalXDR5/OncyHrCR+VTNlSze
5M6DMlPXVEwtoYFF4tpwLjRahnksFNFGu/oR9NEsJJxJ1Ou4LnMBkNjKsVJMrg/9neWyMParRbsm
hNaAojT7mwynjmh343VUruZVCi6vn2LpVoaE2Za/mL8hwWe/YWGWGOKs++uLqTvwmR+Wi0UxF+Dd
0pJS1T123Nm+i6Qj1Hrh7Nw2rcqsfwBi3JHtWYVJ4R3WdrutwktfO9/uXOCnbEYL+C57uayxAa2v
t0E+3Y3IquCmSGMPV1Egff9aW9wifWwZ+RrNv2smVF+MHgPZecd1ZAC5FsSJoW8LqYo9rq0bL5fX
1kOjoqtbsc3jedVupLc5n5EneDpi6ubsM62D9eRRyFBNZzMbC4QspvpZi78ify8M1bDymKpRG1U+
B6TUcFTgLFL7aXQogsqFq9T0N36b+C2htAXOMGuSrvi71Ul8lknpLCMpxOpxW3G+RI1CVhG6IJNM
55ic0KzgAIipywcA4dsXM/maZ5XMH6zqyzwklI7aakr7JO8imXubl5EWN58s4DkstoldBLZgzvtJ
PAsduFBP18YoBi42X55s4Hb9JtNH1K/x9oWLKNHqfrlIKPDfFIS7xcGp5N/6zIOdO0T577l3SJ/W
guuFsarxZV27fRv968IpoIXRxgYN9K8d39VyL/NRQwwOiyccczzVOw7dyQ7Md3Yxi/VE/nEoumqN
6ClFnM8HELKCRFwHO7FscIOlTmGcFSTknELseO/rLYRRMRqFv9yUvGs2TCPszMeofYrJCwKDgj9l
X1wDgQp98meZNGb0q/and+bYB8iX7wILPM3H06A2esP979IJIfGjRlr+Y2a+kYMb4WBe4WQjU8/a
dwikV5kdYqnL7jOivTkpHvpyj++t/6IHa5zbi07spa6BaKYdr+9dTiCDrUKA76E82R4BDrjUfkCw
R/zB+C2vfmIhNxbLwWI+a7wQR9cRXhm/nk2d/UCyKA4oECNMWEYOR0ROsP33dVRpQy3McPkcpVWj
c1aAk4kfb4SLOn4dVEra70K59bJ6+LIC52ZCR7+G09QdhYU9ple0ht6rnr3qADWlY1yWpGeV9Kfp
87Dh6BHA3ixSwZ1G1gMJKBOHVlxWh7pvFUp4voP/HUjwO6cIfIOy/079EVZjEo2VNjG9SjNfWUZP
JLCjVXkd+Nrp8BaLosJ3kcijv2G4yhfgttTbV0Lk3kQ0U1/63LBTUTVhbBfz2XJAs35fHQiJiuMU
vqyzuhlAzDZTf1xV7tsSCZyLgpcUFo029ETJmbNF0P4NDW4vAyvCx+jaaccLZ9bJhMcsMkK7iYu5
o46t+IAmJ0cPdUMiFIHEPRuJBodPTJhBAsxXoefYe1Vl2ZHR5zBsQOY0v5I+yJtYgVV3umc31qJl
SCLLhOMd8SAbtMlGWjcNNDfx1ruz2+rmJtByrMMaq8sFix3RlbuMHmhpnVx9TXtyfwi5vGnLhnFT
eHj9Hp2fO+iDJexKV7Vy4W9YIHXYEJskXqUkXiY4X8X8XdGkmb/+cPcMG3tRA90PMRHg9XsMLcXR
jdaXvzOn6GRCPmLTho10xW1y9Hpxo1he7LlAUqEvGioSVYnxhnu64GOh9ccHb/T0qsPzX2rp1sSG
Q2iQirU4InYAmA1KSGkq6ljoL6SrDi/kcxvu1XcucKJila8aTkguyH13jGpuoneD6b/ZIJh1juOg
Izjw/Grn+dTyZYw2biiIonkuncCKw8MgXBZEVTdg14wpABa+LOO5Ncd7oXe92NLxLU/0TqGihsXC
XAkb9MCYD6XjqSq42swo2S2WTbUTtjmyFN+jbWlf6iaZxv4u2SJqmgPXEpm9ArD12OsfySXrhQ8h
d3e1/R0t1W4ow8EL/dD7y0kibwN6eaFtNCSNjxy4UVEE2AZBpak7ri+ozeqRBoIgzFr9Hntk13P7
iDRvLmaJc11m+1+W1SAcUEXFlqjsC6tU045qJmjo8Fc0sOOIRvdz4ffgA1FRkvtNtDv9rK8qobSU
Ktxdcdc6BRsG1AALEnXAzoYZrbGgU0lbinsy4xIYF3fqbgb8Qe6i5E90c8vZvT77eNnepawO6rU5
Y+aO1ZCQEGqyAeMjwCcWZbrgzCe/+U/m7CfCXlWKBv+RKowWDDSPi54CNpMuLuxh9ijfJXB1E+Go
jBz0/iROYuvgnNvSMd77TEIyE2YwM4DdNfLSjj5MrQaXyJ1zEECa2q+ZcFT0YMvUyCZYHsJDCKU7
fTjW8LQtEzFFyIlGM+FkdOUoIcQiwYzFUHaC/4dGvdEJ28gOSX8yCwCruHTUhnKbJnEHLtjdRvIZ
uYJ80RaYLlm9nKAr9bxuEV3wyadRJ/eugujRt3IWvtCS8zUVemWWjARgB2qa1QSpeTV4z2p5avhK
0mCtNovJjrKS51iFsEXtii3UtAgUbj02KRd+KrzyO3dM401dp2mAHb/16Se5HGsT3ao614gWirJg
UarevMH6zCXP9KpFbp5MuthV8ZYOa2CrMGdJUQQDNwjqNz3HOrXRDKe0LIXYowkj+3aXZ7ckGv5L
FtRp+cFKmADAZ2hM/lMs1xB6XnfoJALyb5klmwP2hevgqViOdQUb5+kP5w5xdWtT2PeFhsto9LUg
3tgtYaWXEkBAbw0gmFOhaGA68BWPs9WRlmxea6TPPzLiIgLMOjPX/Zot4TDNGD35yLajcakfRE9U
8dpJ8d8w6CyYXxgB1jqBPji2cGLM3Lmq1f4X1rK+HI3LLJynN5sGnvLAeb8tn0gexlNH1G7c/ATa
5NxNgcU4jTPjIhdbZmbuqf8plGn5/uXsvcmybGcvciBkFdPn7hBccVXHiQ73wF+RkmbgledvFclB
t4Mly1smElUTrkKSvoCYsTPrJIG+Y7vPsQFDPS+gSJEGs9dYgqTAIxpWn+hM2BP2uMGvVlMp4N2N
FG8EczN8G5a2OTs0YZ0t9I5VOEtYR7iBpBgN7pJWLFft63Ztd/Jifmazjh1F3kvTq/q1OkuxCizm
2467piMH/pSuXJvn9L8PE8HZ9saxzqmlz3uO9Fh3ApbwbufaJmcHiE+xPvci4ok48w72+6RuFa3V
2uJy6EceoLXh+hu3ZGYEllJ1OdfIppzdIE6P3w6NakGDcEJjkgrlZkj2+PH8MJp/gPVKmwOQQ/U2
6647Mha+8XycRjOwpDov5KzzTCvHtrx+uAiN+yvqHbSw5qkEKN1zl/ba20EHEaTocYosAtGioxgq
kdNyo+IbDpStXCnyEiEak5wvKscQDKPgyjXWuUphprTToWGLJbQwPKQI5pwxWIROsqqUdE0TJnjS
Qj1WvTZ2ibJpA+yVl1cIo2Pl12Tmfub9WmAZNFEA9b0Ip4ISRsNU/Cgjoc3XQ4pH6LZSbM2Mr9TR
75QgwTAzyZl8oHNoMnmvRSHl647ziFgMnOhVe0nrUxmmW4s9JCgHRVL8jh2Uw0WrxWX/MzW+PDny
TIbMsfxoLVIB4vEIF/aCjmc0f1ZU5S0vl9+/yHzCweMvQMJxWHlMho6x1DEcNZPnhBJiGom7lq1V
gBdAyzgtfxVrXThY1C6D59vKJGDDiDuypcKDpqQTtgDlnKO/Fxusgqiw229vsE9H3Z+bzCrOQ9XF
ieGYDmVA3JbliDvMpcp3ZPQdQC6Xg52h4a+suKQ6zYVicjQ3yjT07l0lsauwZQNTPSPPNCgYrUgx
eO9BpJAOIdYYBUMomAtWZBhkUO0Xbshm03+vSre1TFR6rq6Jh2jF+1qTafZDBUpzmoKJvRX+MrDu
3yQXahVr9bMXV7U9iNeHpBL6hXe+jngg2JWywFdei38ARAX8Zo28NfSlgY8cWOmRWCjh95eNnfHB
E5ug/J7Go4sTtShIBSNIudTLyGw6dBH8x4y9aXUXWGq21CG/BFHAIRjQTe7U+0xhuso2pjcf9ry8
AsptthpycsYi9h7htRww181lCAlx6bEvuRGjHzyUnvd9cSuh5kf/UySRHrd6lnOhjvFC7BMYKfZ6
yRAbtZMdm9vucqbrq6Mqbc9ZRZj5MEAawP+L9qxZ2xNgeNZpYIYb6zxmQUaxoBlsi3+6VR7GOdwt
iWYyTZanDKvDaSkkr36Y+kSvwAoN8MFBYZ06MxXK8tmCFxx7+OFdAn2CHzJudtcWYOC+otnjEeNT
PNzzosIZa3Wwgra+yfC1eRiveHZnaue5cJPC8Zonr0/UHV3LTHB4pR/pBuebq+kCM2MgWk6pTY4e
I0qxy3CweIGP+Xni3rjAtI/dbvMdZ21XGHnKCfhTJWYhPACDZS6zNprIOXF218Egp/lK05gLLQLG
RWgqBmHpGt0u3joexILkSY7LOpbmzSDbEhyFXqYfFP/fhCtbWLt0kmWdif/qaK3dBDyZ8OxuD2gs
M6Kb8eUnFAqgQkNNso7kAyAMRHs8pSLPkulkNOYMSzm5OfQ4KbamU2fuFkzKD3yKaSym5n9Yokoe
0+pPK6EfkZeM0/BpyTYdJPBNbpPLwOFg8OuwdDjDDny9sdtQ407AN9dZjvMf3DQmHtAMcaCLCnke
ByK2HZ2+9c4VDxTBgtcWtq+QvJH2bU5sQhc8PQH7k5+KgIdCTpxU+2kgLb2CeHY4eAvN+k54Z8UF
xgxzqFJClUcShOd8azuAJX+DEwgdFZXI1nC1BEZ85iao638Znt5iWoitoUhO0btMWBGk0vq8n/17
aEPrKX6dA7kNXTdkqBg70bHs0WLUhn16hUBnDHRaGPMlKZPSthlZFJ8Q5HRHxmD7blgGfH4As8NI
GCaNWJIhXgmVbN7OgxtfKIo1l4XYHfAVxMvCQD8rYQhvNE54uI6NFW2aCiu7WZpCyfRujs5dRVDw
RM9ie7eeogLyETXBk8HZe3Pj0uCVIzuuXnlhg03emRBTckdIfP7fzpmKk0+mCBmbC+1dgAS6Z3nX
Z16dZj1Hu9LH3rq3F5hPwF8WdvwVyCg8Z2vidvZo9DiEfZk9vnSGhvTiGLLgfm37aIwdqFTrPfzA
9tRoB4Dk3LTTuVL2c5gTx401Lml5TNwF1oHaNvHx+kB3Ce3bW5F+q7r1nZ37tvSzzdwyx6IpRA5z
BGbAhsMWYZFNY6vofGrpRSDCNs7bCldw2MxXf05jkJ1ckJDj62k3WorIZT9T9ngI9b5xtQtlRkXl
H6Alnuc5SbTZlOLziYoXEJa/nJmxF3Vbfc9ZINVZ3Xe81BqBGed8ntc3XOI08G47LUZk/FrJo4yL
c3V9eHQDeM0nZpiHtxD38xxFCNqsdpmdW86A8C+88/uJrS8vU3sK28oJSjmE3MCbrxV+d54gnssd
qG8/lsHw/AyMj2Do4/PCSDeqr1Ga5r+E1oB2ajQM1q/GRl1uCKohn3MG8/+ORqoKNABnsVEXzDch
5nHZPspHG49nTmOCL3dg5Ma93G0YpJplVlIFlYdA3jga/nXJBMm3sT7pvBvgrQhyllEyVrWyQcol
aA5WxKquhIBsSW0HWPrlYtWtDARdlpJ9rBWExvKL0hFNEdJOdiOawRLkVgP+uZT80dhVtkpx4Nf7
qOHCMlpkMfdq8VOl494cBuLcbU0Zzuw0nQ3jwtu+q2lC5m1gOtvv6gzsbyW7/Sd6xwyd9wek98TV
7kj3B8ICKmjBVHKWJv05aY25u63QFJVoJ+9JmcGgsoE1OEIpBxm7IynUUlmwF8S5UYk+uzhExl5C
UnZvssbBI9rDv98HMaxxQQYYOdZd7lNRDpivdJVNgUXWIuTpm5PrqB9UWBiOS2XFWwUWD9894cSl
BfeqyS/cebMU1kU3m60v2gScZ0zPGaNSnyiF2/5QQf/8PZGciSnO+wZUdqRWz4fdOqlTpicWPaFZ
2oK4uHfV0vfK2ROj1QnJUvcaZ84NEzh66CFUp2OdnqbNFdfzg4agWzEpIbhyM62PdwdxUy7vh2Rg
ApwKtONUCavnA9LedgC3vR8tgSOnP09lvx223Hh72jnCR9QC0KZGg9epQ+/7YmrpmbgA2m7iRFXt
6KzL4pbOwT+ks9XIeGioagX2EMvl+msXHQSl11+tADkXj/EU4YQfU/Nw4raSTknIuSDC7bAZI7hO
ZBtOVs2WuwmnkOaXrffMtACNPqgzFINaqXPJDUeQE40J+U76GAagIbWvIsjeDidqV/vrQwzz1eil
XzSFuEyqHXbCPMDdd818AfkieDJuEBz1VNb2TnOOyxBlfLIm2WNO2C9mVL9AXSHaoljX0BFBQ8xT
2TZ5DwWwX6dl7inhnM9qBDK24fenPrNyOSmqjjwnye/leklgpkz6enTM0vE9kRiWzIGRu/j4TtfF
C2xHWhR4/UGJEyefIiTra4z9WrCNHqRC3qRE07okdDwO/j8HDDfYjxK9IjK0hbxR65QKqlbKNZ87
IYH1A/INl4asg12Tce63+djV8vzM0j2CPif16qzhQmNPEYVEJYMwsEfyAbIEfagbVpGJuyXWDhh5
LqcPTmX0bJg/LTbXbVv0zUJ2jzxS93zw8Ek0Cn90MUr4zPRPmuC5U3IneOcBx5HaO4WWngnouWVd
2M3STM5anVVXFyH3pyiIe+wBLUVBQLBiyLv5iUCa42L7kYTv4VhIydL4tfslwbI2YazFVElgdLZM
0cQ+1pp8X6ED9qFYzm98dLxoUFl6Kwo13dKfvTD/4Btjb3EnZhKUsXQTXsLkU4ReXXi3ZiA6A/+M
Z3CrOIUn9Ieuc+Tfklkri3347V1PPgcuYjiqIeuQ99E9UFB5iQwj5TuGWCafd4UsM91TnqtW6nNd
bE3py/qel+jrtnghrmcNDN1LdS4vLWoWhjn34geFhjrzbd2kZehg2GzHplh1VfIFU05iXpdoKXdf
+hiNhM1mrieBQ7OWCyBDgHjLKJn0wuTHfl5KtHUgm67IbujjRLegQBsRpDfmLG2TGNCbfeWZCU13
ukvr/vn0l6W2kqbN7C6PPzhXB+11ZlSsXYprAcIWKHjTJPp3TR88g7ZMDeidmsQUswET7oR4NLzo
jU5amzXxjllF5hwq6bdaEhATCxC5zjcHBube2yytedno9H/V1q2ju+GarM1Sieg+FnvJWTlE5FF7
kNXMpGvRY4f69RGW5xRQzQwf4wVdibxBuNQAEzGB/k+/128FvfnapEhZ8GxjPe4pJoxNmmTh2aLg
kxSIahGwfx7wxnuZaxiKm2G+UlRvQLm2QztvBSM+b4HD4Irve2YKD8TwLxxpNW0AqaXfuNF+UsI+
aMRmDPCUhoMGt1Ev0APj7JDo/AIjJQUAeOgKCT80aY06VFLCdWjHeINb8JlXEV/M72k1GtwNrYD9
gnFvYKM4Fam64sEVetV3R/MwBc7dKMhgtP2N37z1hln9F2uwhHQfC/rEJE3MIFFFAVLm4m4jYXWN
4Pvh4dEY0NIcR2PDrVQqOBGCa9y0U1qy7JSjNo2lGkw9gPEzcCTqXapPNl9CPzx/C2YwY3xlt6I7
5onAuVCSe7xjxXOvvgS3prmoZkQlp7Bgk7CJnfyRp6/vzTTRyI3GscGKFJ5iYl/zfHF8UXCDo+ZV
RftD1JS4V2jCxz7RjYOgyhHgJddllNLyoMEmxs0YoU3GcCguzq4kVx9Gmy2lpF6ermtr1eWk556c
RE4EuzaNuFIk+pKlFqaoaxKLWVKDTp2m6CVMAvCEy3mz6fcV3xVyaOre29GEj6DfMWgGnBEAin5F
UQUht30kodeNIKIgMeEuhFOY/raW5TptZRncE8J1pNmKXXVWSaG5IrtO7E//brNDYQCmW5GVYxhw
mkg/lWgHQ0JZp+9SawXrE6+i885AqeAsg7Yh04e1a3U3lhipetcpKgqJ15bVLX6RVJUTcgXRHGqq
pXPEqamfKPWhAGGdRGA2kZcfjhoEZtOqSfpDZURmi9E8lYmNf908/sfmx3yI2ag7SusThWAI2lFQ
9KJzBa4RXqmDIRurhJ8yZMA1cMWWmr98jOsFUahI8HOK9UqgZJd2h/ytTjOALPNyiXVm+cFWYKuE
VEmo7EvF1Pdl5kO3hnfXcNAi/a8c6A3JtnTPhLqtz7QBvBasp7YCr5cNggCc4OHcKwlAFHKz7WK9
vYPgSl6N/ahGrtZSOKskZq9qaTq7LHxtmvOOStJO9FlwgelQ4mZ8PKVTA3ijU0C5fwMFKnu6bQub
r7u7OTkO4oTCaa5RJEMuIQ1b/9rAdkk0jeGtN2HrqKu4NBKwYgWTD/tzA996cXEQUQ2IeN+qxOHY
MZDxjqpSASmd2d3wTkEuyXVaJF0AWWqI1TU23KiL88rAFy5C9kVBxeAoD7wJojvlu6xeM7wehId3
oqGMj8B9cEjPeIw4L8KPUszIk8dMj1OPO1MVUcYKm8DQMsOW+ogGjC1i1ZW3APxTpycoK1Dx0LLI
tqwoOQAtXQBO4pxmRi+Ymmuv5C4Gz1ezm1enct+gKWS3pL/OCTvW+ST4v2BVv4COvl9yJ+MsW4WD
UoN2mLrXCOr4YheI2Dsl6/Xr8M40QNRl/n2cLmfWKqJq+3kSUPoGc/Ad9mEiPBisBlaW6z0ct9Rx
vJ0uOY3iMOrj7QzoMOVImO0hwbNUi9YMEE883n5//hWFr5uVRy1Xq0xMi/9f3bMxgvhmVsTkLIEh
Y6BNr6BPPYO4UtITXxzdyBRg7uJ+YHI0pTknymSoanx13UhTtWt9n9gQjGqhuxFP+PkCPoZew8lO
J85SbVN6t3EQlsNDqpUgzrOqYf7ibzHOvpfCcG61oNo+cSJmf2eoiSELHBOLe9yaLw2N+WJjusBj
uggI/uwCKjd2UaqFphIeL2C1EY3+BBwp7WWe3x3nQfzSeKosyZ/IAviIQDmeatOt1OMcoqAE7u8z
Zi/y3Z1TlMCF1hzYy20B6yOlKqNthIf5Qah6c+YJbtANujq51AXPzy+Y0CoSgZi4lUc78pTBMiVW
x0pPoBGImlbpqWJoRwjCyK0xWwCma2mU8kx4GplGBiid2EXtM1qEXcvgoT2OYsaHQbs73FAzQ/3T
LGu5uq0BomXeuv/Av10l2ezOScga+Pkq2S0YJOmDyb+mv3c7qcqhD8NjWbLvMFADwbv6z+BLDhpy
oxJL1rqd6dSAEmkEcAblxztaDR8QU1BtFNk9wQ6jgFQz3zVnx8S6fd93zPTfZH3fdtOoJRX5+0f4
yGQf7GTchyL12ydzoYZwH4DNiVGARpv4U10kvHu/zI16eQCJ5KaWuxMVc3e3RAIAzYc2QawAsDMd
lFiKY5i612WZzQBMZRR78mV3ZjYWcHmYwGu0jPbumA++NEgFMYVPsHFfYj7yjOf1OeYQ+g6+fmgr
KaZkxk2jHEs4/nv3fSWbGgVcmY2GtP0hLSxvRiOoCBIBA33I1lGNBWFt5yHsI7N/FR6vGyD4eVUg
y9nvzWWb2u+6Mk7sgEROz1X26rtsakjQhEGUV+te8Tiw2cQ9qwkl9FPSYpDzxaBT8XDKs9HM0s82
lGYsaoghB1mnbtS6/90wCiL7ODuwpxYj/LRYKH0Q+sFEnJS374WAp6kfRKifNsotqhQvmSwe7uBM
L1rBwpivzc87kBxUD+7iThM5d50O1DKwI2TcX74XlO8betNn8fSDUP3OY0ZXTMYL8ywm7Gey9tTK
hRLFIjTA66Q2qbMt3ZExfzQL/iNykQTvHqaRgFEJ0aFjEOWe2wRCpT6GktTtrPQ0LF1lG/g49k3F
aKweSA50Cia9xkCeUJcAmzd5jgnyRFYnDvEeDLiaDHzmMRozM/caP98DQ9t7FrTzsY+u7EQ/+MEc
9bM2yWCiNI0b3sN7mSkfMkr3km5NpICtkgvC7oox2pE84J7Ff3oG8unaxqfib8xr6SgqwqpC7xwz
Wct8Yjnyj2TcX40TLw8w1VNPus4alMhKQ9C1cvpByBVTP7XB9srL8EhRGGLUw9kID0pns1DGUc64
cnU8f8S7UxbYQb/3lV+zD6W0IHEGC0l6UGhwrCJSYHuUDgcFswkLsQBL72VXwj39ntg3a0ag6Fqr
NWHNbkxvSFpksTFfi+HqjEUPntnw6D+Ca0ivTIdlFJGaahAJDnrbLiWTJJHbX0AqcVCXaIlpZW9K
/5U+vSaKiZfhyJqX97ZPAv8PpLLnmn6gvXwiqzXIvGZ63cBLh8LsTy9ZHE938gwpRgtmt1RCJ064
IPgAbHSkryhNV7Ui+nAcA603orqZqy9l/GIRi8VeKOr/wcBe8ltQB6OnO+oaW8YHwQ6lIzN6oByC
SMOwJbGIfke5BA5nlScWUWyg+D4bUBBscPaCl8krXKUF6gPqMdCsh015KlRfVu/UnyQJwfM1S9P9
Ac9p/Z2EMR98eaw4uaAtglPwtmgSg094Ew6aT2tSQa0dPi7kGgrRarWOLXVDRVryeOy5dIqAr92P
GLIkd3471mRRGsFXElTBYcIFR3yx7CZhoO13wQasLc78qOvH2RFAnnV3xPEA6ydz8gTWeVFbDynD
Q6cBHA9gJ365lwEOA4GJA9G51Qre9xPVpCB6mOsyBdUfs9dm0awJlSbP9xxCh7t32X83vE5iFScN
1SdIhRR+H+duYKLDIf4BKq2U85g1xPkmsDmVKAnBKeSCgZ22g/iNq0NwRkwBHpr93BNHZDLdYdR+
g9JeeIF7sm/qNF92z5U1PXGXpuP7z7jaInC3vgTWd/O/TekjeNIMexGdnk9SS/5HAtmjYOSzkpP+
vUbYTSkpgpEvVmL6VAfRO3QHgzTeTYF+Y4FRRxyXwEswi/LTCZGwWmg/SQeUmvNBIaiRO2FD2MEf
B2T/nMjeybBrupGBBian/uKVqImXe1BeDg/9ii/nofJbBtaHVu6SpJXN8WPTI7icMCemcGnhBX9L
gA1hIa1cOnm6ujy8FFTFThraEPTkKW2Ja9e23uvEOk5DPiiwXahxii75yusMWYugdoP50b9IajZ1
U4DULQHjDn975DanqSv8uLejx3q3Eqr9o1xPLklDQea6oO2S4s5Kjw6CXHuXV1Bepr5r1lcCY06h
rrstMQyZxwe4MN9e4k7CjnazrDA0X3gq/vxDrYSCxLLnSrI59VrvpVVFUbJ6RUXqzlyUReUxxVLi
0GhiezT5cxJDm3LmUCMsO6asX3vAlW4+eZ9Q5W2uIFmwkf6xMwSlfKohb08HawFmCvaNtynkDTVj
QRSGxJv9kD9R2YnbAhqOpk4mWU2t1wHkzAZcipjuwdYDOJ/r2MldfzTTNuUlPCkMqwMA0nl8d5mK
1VhND0OagRuoR4iDYpsfuT/Ur+19o0g0VYdNFdJNh0FjbnhyVbZ2PR4wW4v3RfDHJM59R+bmJpOF
uMPuMjCPOzQxrpK8H/xyxXJAPbQf6ftujxK2gliz4/2kdupFguSj4f5tilY3oOY0uVm/udLHJ7W4
1m0tHcpR+z6425W5r0WcaMZ07xMXVT/7CKVXNil9hz/kVIXPCAA/ajKFORkpzZprW9GMKi3tDrpg
MukRbLPRuEfwwkXIFm1Y14fpe9w2f9+Y2ot8HHyx0WF7evy2kMRI+DJr3Bxbvjsfwi8T+H600XQ2
W6mQh8K7mIJjujTLcCBb9COMoROw4HjSZ5JbuRJ6PXMMxAZpTG/ANLKbZEQQeUkRQxgLZs+4I7Vd
ZZ0BkL+UaPZwlz0pk5S21/tte79g2EqH8PMFpaZJWXSCCdFNnImbhaLb5Mm+x5k79deNP5Lk4XiP
EM6W3UO1BiZubmHNXxl8N3oiaNo8uzIc4313mSsn5WL0zbOY2zURfflpQl7rwQyQImvlrIDwbEcv
ea6p3pvnF+AslhcOKe3fPpvlv1e3sD/bRo1S95IsWPD0MPw+e8iAtqunae0BoPV7vF88zt89Z+4e
m8dBDmZN7oVQpRZORZCxkW9ShxQN6asX6OeG4y/XiAFMrqI0O8QUNB+zwcDr9BH6Qyb6nlQdCjz0
LBisN8xfS5fVVcipt3DbBPHQYfrObtflPXpx3fdcKAL5D0KOxRrb6f2msUmrAIHcdKr5MWK4+qcd
8cM+wdh68s/XPCnddL+vjNvIZ6KQ0H4k89jVmk8ywMKBRqnNJHn0J3FWzLLqJ4qoVmc9k1xpBeiN
n2MhjNuraO+UniZq19MFydw6t0X9dQ9N98O6RAbiExFz4Wot35NOxgrkf71FZ9NXjidkiulcA9VG
t4an+V/btIuRgmQGMeZ6L8nFAB5G783xUkkjwSZu79DRpyThHQxm5xR0rKfhMR8UfHeDQ4ArbfOS
mbWH2vjynMpN/hnkgJtZa7N9hEPCddl7QY6VmNNWjGFYHqd1VZJlV5kpR6v8eryxnkVeQXhQH061
hDpZDjESPiK1a5InMDpSkh0E0+sTFUrg/InZwMJMQ5aRtO8If4KEw5i+mCYP0VjxHgmHOiVcLwdF
nvXHp02TJVBHBpZ8e5k9nBNarbW0TVtP7uBcs9bkueM6qEwwfBcznpc5jpIg6Rh1VfNB45nyDR99
PvugZvXfuLlvM/TJF2y/jerGT/Louhs7+Gsoiku6fsX1RgdBM0PyFzk9Rd/efmIcONsOeGvu01He
qkI7qpHs0vWmlbYsB2kmpQPEWOU892l3nxfpOOSagGCe4j6uymrh2wKyz6pUmxn7gBo0eUuhXIvl
DrKrRPM2GqDr5oGBmt9nfdnIZL5+mW532kjYowYrSsTjdmB/f7zZfvDZkNJkuzf/dIfm4FuUEHL6
q1OQ3NnIHLSLKXq/QUG5A0f1IjLYaUXU4JjlWb7ecqWvPLPaIt0cEYqhI/T0+1EJln1rb6PwGUWa
79tjzOFFqe9tpb6Uh6KWLEUpp7HJEj7N3aYo2YUVrjLbKuVer/xs0SGWja9ml6m7u7bEFzO14Lde
iAfdGFHUQNSpmZVUlzP0EZCELvB/6Xaa/RvlNpdRyg0PKKN9jyygTX5/UnEkxFE0zDbOKTvHfv01
rlYXkO8NaDHgWxIvimeJyddjTVMc5NN4/zV7hb2mZC32wZP9XKVJgwyhjNjofMWzEvPJaLk28mL2
m/GKLvEyM5tIJQzuMSidCMaQtqXrmmkqotT7kLLuQLsYwMyq6IRwhjsbRJ6XCM0Bz19gQh5U8rR0
g0epYPnQAIb95pgE2gRDCPFEXCDhnR2DSHV3fCwRnwqFSsYR13DVykTRP0/gBw5Z4gsrlru0yHHO
DuJ02Apu/YeRljDWIRxc+/A4TH9kbETQ+S51KOcwUEPLgiG6T7ZfUDpw7QLiZaLBHbDGgjE4Ea7q
f7iCrMsdW0++g61tGgP70TwwmdD/TvR5sKVJRt4MpebwuAApnhWmNbc1UZFvvTAbrVbWNVTXKYaw
OjeMOSs0TUrkjxDSX/WVIMOwTUx77ZgWK/PvRmYg00l2Mf7qqbk33u7zMux7cmzt614P7P0Gj5v0
g6TYDIuGvbZ/3ZUCh7RXkhZ1ZUM6pHJ0wbSapk0X64G4PWAdq0xvQcSPmhaMdh27wkwDJSTqfAhO
8gnqdDPhqACy7so31q+NLHjBxG6JzoiiEhNEN7+8bifaHEe4aapdAAmiqX0gtQG1ijAGmDCqWb+Q
qt2bk+YyGW5wvJVbacpY2D1nIWgF/i7IYTPDLVNsPZaM0//q8XY1/wg+WzirM/e5/no7sAgqC8kn
CdK8JKBlIy8TFdOimdNe0h0ukwHJdUopHcazI5KOCG2NwtoCb0virk8Mgnxof6XukHvh1Owj8H3K
Xa/BLsQgWI1p75a5hyXVqCC5BClg+PytcitSug0x1gpiDL42MhthVc12u6Yo/1BlhPgAAIHM25WT
Y3tQxCJd9iwpc6+P+pA3XsBG3WJQn4T55F1pEjhXCsHr8L+FZlD74WEVakL8ASum7+o1uN75KRt+
/yEhPwSk/gVuRmNkadmvPDvevGH6fq+y24k4Q8i35WUyVu9kh18cVfDGlYP4MGHOzIrs5HBZYKfO
FXI1Umg2dtvK4nqhrRw5torurD3c9EaW7DUEISwQR3MnEv1pk98AOv2b2KBWK6uis9FHORXUmCuU
RLl5zyb0orleanwoXaPbzRGDZYHgWpjHnoG0IDWRd14KVe73mB3QkwS0CsrCiNVv+z0+zmHEeSGy
RIF/gJ441yxIPePfmepF2metu7iT/LqJgMW52wAcWUMXEJEsOnepbDaFqzJmqw+g6T8G9EyCZHwF
xBXE1Tzh51uyxL9Gd/VLzzJx4q5OlMOIYp/TrCclxKU2We6RvJVajpuoG2xWxMxTOc5V+1hQgXk4
O8pwOz9ru32QYlskSHDueR8i47TvWY+26D10zcpbiM5GNpFzucJhUQYltwL9ub1m6N34T7j5dZ5C
Wq8vg2ejd9j+lIoH0Jpbof/cPJrMLcRu3vMHII163r/gGt56GA4v972QXfidBtxVwRpu6aDu3+i7
QJV+/+z77B4y0ZM7fHmT0cTcdk77xopiqxp42v4+58dZ4Z8XnBamV8g1i6BECzBjc12lEoXrkxRw
jBMZ/ppGIv1ypeOtr3DbRwz96jD4NnkjKVpZVKjik23mU3yxa52hINB2XVyEhMyZR1HFvb5noXgG
vW1oZTyitgX7V4Wk+A0/002A+A7gjU6lZb1ryZPN9LH0quYnuXwcF0hXJ8psNH7vAHmgwAkOIiMH
Ja/EeaOVWsS7Fozpe4Fs9ddqO6vNbae3xfCTH30lFBYgjRdXey0MMNR5afuRny//Yz7XhvJPfoHY
R70IJN2A/K78qDwy9lRHbcxKnSSkF6p29Syky5jirYOVesV/fjwteS6pVSQ187nNx5KwYWdHnJGl
/KwVC4OarRFsDBcdODGML3GhaKepc1guraDFHui16xDrj66UvlQz5br6CodS1Cx6eKD0ntm8HmG2
NEakJPeqRgpwscLwOKIuG7pGlo6hsWFBWWOCIEuDV2XiZOqopwcVmr6yFN1sZkkMyHKbZ0HyPq4A
CLarLI+uoA7zN9/OYoUeLTQA/AxHkao8q1rBFunH+1m5PUloX9lE7nEVXtrx7Z3QAJXiUOR7SmTe
+z5bgRbpz6ZnHl1DwWwmIJU9+YB1jM0m33+d8SdYL946ixO7a25deuJBjvCIa5w2KXLT9Gqk3KCa
JWMkunPSSe5OQOd1nBIkNMFEiZ8LwvHNL0Q3pIVQjjcQzqKlDTNLK/tPwno2ia5ULzxKmg/ndiVM
aYHK47zuD5vKYh6MbmDPCZ0fSBdcLThKbIzcLI6HGRvC4gnh03i7gh9fqb5xLG4CrK1tPW7Rj+vi
I8V1J/8aGPJ4xEp4sUlj2ZUzKquzwXRmfJMlr+tNrRao8VVqGmZaQMclE7FRDvdhgGObdGsPoTtn
2Or1Qzk8KHyJM8rM9QvjR4bnF648RhwafI/LCmWqFzKUJXl5Dld8F9km4Cx9IFJS6yr1jMlyoFOk
jchpLljv5N4rUSXPOrkiBNSNJTnuui0WY0MA1BX/TXi24mwgZoE2Vpa+zbMQg2Wotj994uFrUYbX
l7fJtovYDZZBLmPND6fF8bLA/ojEiWQ5boppq46XVKX1FE6bgUKruJlZMWVFmibutKLxiTob+UYo
mtziFGXIx5TZzVPTtKRU950SbB7aqxUMOnyMyImEVM2n7BSrC4F0PDBbkbnKwekwuSv2aIBvxsBw
MtEGyxLsv9eju9+jVQ674a7XRwqLAq65iHJKhruc7rmEgYOhB4KqvmwyvZXKefwqibTrF/2sWUVb
OFbp3MPtgD7Km5BObm+JhlMhZ8pitrWe/qEVHkLqYyaxo7Q2Vs1omx1tIyh0FFe8aAeVsvxZRrAQ
lH7CPr0grAtTy7rhgoH2Yqx5bbcewN2shkcCwTR8pCl+IiMkrn8Www5tQxJd2lhn4YRCnVpsG5et
19bJxZP128g8f0P643ODcRLUZtQM/jcsXvIYwGBegDgTwf+F8RmOb2PJTAS2ySpnqGnSKEq+Iayv
0XD1VoT6p8HY+ntl0DwhxlQ5Ql/lb/CF0oWNjiHWPbZ3fPovX9tAj3jqMc6bfPfObBVRcisRlyMA
py7Hmtqnv2pcBUW/JFotrswvqrHkznXN0FM2+JFNQhBOYZgxtYBQp/5MEUwY4O/HXHgJ4qv6/0z0
twKMWnmh78AVk/1efemmVLqtwgq0aYaFlXzIAaGPZ07YIJUgsEpHKkMyVXHLZMaDzd3YKvoRCqPr
tOFtMkFplZ2I+Ei+0FkM+WkJmVNomuihQuJynyDu0YxWOfN+JtJReW9bgwGRA6CSV16W1kVz0RRz
FmEhPGnmhADN6vvgpVlLoSJ5RoGzD1b/UJw0WhtdDunn2C9oGnRVNNPs8TWYf4aamlAQ1WC7MzGR
dmQw0Tt+5gfpGvSRFFEaYvfbMS2N5Kgicy3ghV29ONvjgGF54adiIjvCt8QrcURVuNgIYPFIAERM
IoVsm8vUI3jne0cqIhy7RrMJJd6elz+UfbgW5/zP6j9XMEFyMDF52yWnEt1i/wJTS6sk5YeO4Jm/
wz2OA2myV/YT3eEZLbRWcriCCv6tjiZl4vYbaDIX+D6spnKZ3i8fGFxVazQgo4Fpctr0tMVMSZ7w
g1m0auhUWnIs0uu7RohiZEWeMD1EiQQmu3IBG3v4t4/8ds2AEYEpokACHlyT7qmElOIx5gddQmhQ
kFQ6VNWn3Q64aZpzJs5tLdJLTxSh46eZ973+MbnqXKThtiFbMSnMgXtJ+bi0/RxbgpoBKR/34G9z
2lxTeuxlsSVfvDOsECfxiwdmstWommrqvA2oINBgYk4BEYQQLUs1nGqX1XojqkZiQzFClN+vIH9O
l3RdGAYDN2WBoQO1t9zRu+RQwmmz6QsR1a5Vudj8iz3kQLfouvBzi47xRjW7eA3wZLpyxOxsrgXa
fiWnLdey5ZM3fF28M1ItJtGRPpxvvlrEduSk6Y8DZiJ23DTbwR/D1z7Do76w9kDgHJ/6f5Dji2gk
g150PwIG1wJ+npyZDD/HWcUTcIaBKsF9PDvLvrhIr8QebDNV6CnYx3bw4uuiPoSYlz+NSrHMcsQH
mELsDqbLN37OrjDWlszzdRlIZAq9GNT8+PQxcOxYRUGs60PQrphfRYd8yFQQ/6aeSNK9CbHn6E4V
opaU/7NguQ3Lg7DtLl3ssfS3FDoEGR5kiN65LiNSpK5dZ3EiPa0PpnJXPneue0aN+fymTu+tOr49
LTsRnqQjly73u35oo0J9wXi49OjztVZ+Aumk93kproI3R8QSAmWF+CFH96fpyFwO5F7G6vx6bxaP
eB2c3WAbm+uTrIB5dotGNR14jHWHbZeKv6crHjl98sBSNnEPC2BDCSQXzfB/JURJ0+jtx7c9Ckk/
DTJjpy5HGwe6Y3j8O5o/u366qKoy9TOs2XZ25l9tkGvGpg1nb3vWP78zzBNlmRmYsXVIIxexDqEv
USwhf1wGlQo8n8/r4x3LeJEzzbGFgiup/djQK/ES+Vo7MW9vJ6KMF3i/xPnhMItLc8f0D5cUCupg
KWKxZHKuu28qfmIDFVfK/eitNoEbOpGcBdcaXbaTTPh8lptCoZhbI2bp9yyZK8URgZDTfaZZQG02
I0OWy3XNmK9WeCj2awPUzCMmCkNMIBG+Io13MQsGHhQfNRfqZmibsKUx36GohRgF+gUMduIVFPI4
+sWJljJ30KObNG/MSmTwGQZoutuOHl54BhcW431jYkv6PjxiWWbFDppXRHVtKGt9rA5niKBliKIM
kbsryy67VqTbrWrR1ScS2r6rY2o4e7jM9emTS/4TdgctF9JmsL6GFykonlIFSGaA8pQNU5Zw57KQ
AfA7n6mBSo473dUeTari/eKFzkNMzeq8KDblAvqF2wtx7u5Z31w3eivIMmBw5o4a9xNoOswvmQ5g
7sqKEY/OqeccPtTMfu0WcZ5Qtvz/36KO4VSV9EZcNB0GOnlyaePFSsT6WM5bFGY51GmtupPo/nlf
A0zyRV84VPoaxc5EdfrCDGaql9a+TD7VdbftwevKyOY3fdhC+q212V+r9MdpKn1Hm5UALz0G4Iwp
HIWty7gM0GVBDB1I+qSYMaKwt9Qs1ed/wDidSObCoWAlax5hazVLp4NJ2C7KczAhIwRqls31sBXE
43ICNt6uv2oZmPqU9+jZbWzt3pZ6hYffTKFWOtXGaH5DhJ5NkE+gIjSF3Y6JhXZ4VLa3mIeJpigr
1gUMjqNIoERQtLlF8l/Yf4rd79R0cqdGnU8T+lQtxGeacu27xjW/Hodhv8sDq7MfFd4CT8ZGuZEm
jHIxHYefyzPmblyIOg9gllzFqhG0mNGmCsK73lbT0HYTr0mpFASUYTZ/7lCSXKubHqZSKJvJK48l
fXvSAKwtTD4sOEOu3BF9oQmqex2bdR0TbEUNi+ao5Ow/404R/JJGJ3M9L5fhkKw/jVHNOPKglvSz
v90e3QsBW4prK2HDpgbmgcEA4XG/bBjlv4xZEjGLNdg8L94rlyAjL+BYDchPSCfCQqHAxgbgBW4Q
BUz409fQE4NhMW8X+ei3hj8WIShmsRE6udKXwggLIQeVian2qaujfcjMNds994JLRfxoIgUaRsQ4
+Om3Qn9/XLFWfQzbttcL2Hrq+4NCNr/i/nkhARgTl154QWgTToyZpAXFdWUvvcbJ+lPavSGZjpuW
BsTUsGbdypJNyBKdwZGLwbaIXMG2CnnBnFPwboMhIWo1ScvxUFTVSFVlyPYJ/A99CJy011j4Y8LZ
oPj9N9K5H01Hv9jXNNy19mbD6gEDvSn5GXDVMFxCB54chJnRYzFwW4DpP3lYqz/nXWBsK01MFMxt
f+x21yzmPEiVj4LYqeMjk9WnOY5uRYQ1OsDx1rFDjpMPb6/BY/7DxZBS9KWekHj3PYLxZo0Ruly3
ZZrpJ2zDj9vihLOFAnbe/qQuVZmOyfsBQwKEcs83XZc88+zFH78jdrZ7YQBsfbphuqAzhfhR0s6A
yPOk5teFVDGnrpkcGj3pp81/aFoInntLdg+eVNmCTowlZfjAsy7i2OeSHI9ycd3TW0CODRntAXF1
HiKqfzV++5vC77N+3pxrCoCINjpSULSw1bpLBIqn2Sl2lxg131ml+Bfcv69GHNNmRFcxdu78NXkZ
vS9kGxrHUGt4xRAfNCpE29sGHXN2ZFE6EwMqH6rR/mXiB2s5VBnJxl0Jc3Gv+pgmCiie23d2d+FW
B0scR9AL8msv8rJNHcvu0sXf+6vLrUaUOr+0NKOypZOMxbaWd964nW242fG985Jn8I/rKkqpokmT
WMRxhF4tmQSJIi09BP+ob76ED+Y7VwjpFxWKXI2pPWQK9AdPwgp8tF93mE14zr1upsJV+oivAEV2
XkGY8Bt9TEK4ZKvjrKOeO9/yYgQwfslVjkPNbyEX+ByMknxGtLLblX1lavh5Cbm39LdymeMawrC/
4E1fkYIt+I+RTEZ6cBTtqQMbdE2Zqn6NH7CeRmm+E5qZo2ReKmNHTh3a/waCAv1htmCXlpLUxmB/
01RdmPav6guysakOt0dVVRa9I5RHmk4SuVT2kENhQpXQMQwHtEiTxaw7kdztvde0oAHo/oAwv8XB
jP35REXgRUEtw7tety/o+SqoMStLOwHcGQqg/Mi+mzbF7iYhxLkRcoY/+UjAAMRtxp/j83kah9kJ
wrmrscI+Bl1+m3Iwc99ihK7cfaAaD7VYMWjMyMt0kHZ8YLEORgA3jeJKOkXseMlnjEcq3Ad1AtqT
7+foHIbWecRxT7NKJ0N3II9WRP515SSv3bAc+2YpZqrtORCp2BVvNucuo5cADAtMPBBIz0itLSia
Jq3dGnCfIOnL2jOdOpA1mALy0K8Iirx8PQjU9mgNZq7p4ZxWFcbdxroaoBIjs1JH7XMesNX16Sxy
8C9I5u1W7z4Wv/umiOaGP781HHwqRTiDhN8Ni/zS5UzZX2/iqGFDO5DqLahd6Ttgf51ixZHrd2XG
+A36nvJicBCV0t92j3+glA6gziCRgpQHWNCjY76Kqexw5R2K+87020RbBnZBX6a9jIy839WLgr+2
vi8MemZL1vV4KhLteURs/BwFz9cxgRh0mKqKeIrI984eIwL4hOq3URUCIwN7UO+qFuPJf1QvIbsY
nCZvVq7X7H30568Qm+FgczWsqAMLHgsMUKp62EMxOmGLVTKoHsIiyGIPQKg5RDzwf4WhT/690yXV
3y+/UsW1yS1fn3l5UtDCCooe/h7GpRSbFsPmrfKp4pzno6YXCNwoHxfBk4P8klhB31X6Aglh2ILn
9oqtAMiGOM1IQrAQEQvSgIr17BuBuz2m3xvwedAF3CA+kWLQrggwRgAE5NyvkwhADZptdSkbbQwv
MPlVRy7L459Jc05s3Ov+mLYineRkLlnWeltZteMaM5Am9HN2xmf7q+YB94Sl/+3U+pNrmgW+7Wh9
BdMjnomielYEABBwXEZxEpTsO5va2AGbiLDr7zqVAma99gWgF0K9+2yFl56ZdwjPrGbbklCTnJbZ
Si6KFIG3nccffcjs1Lw5FiqSPFoVR3nwzbanaR1cG+0a+tT6MAeZeJrRCzmEpFFMLZ7OiVmlPylX
TWmqo/RM9+huUPHCg0NNW9Y7nbz4BfyhAOEs3P5aWskXeNIVNfPI6lCQ1aNS/wa9KMYbd0K/icix
OqgI+suDu3gZ4LcGhEc5ods8SZIt4FEDFmpaGQJDCA889j+Ws4bB9pOsRSpMIXC40brhdpXAsU6J
1+FLIm7G5q1tqu3r73aru+8ShuMkXSZpzCX5PfFarQo6FTjUZu3Xtfo/zf656SDg5OffFfPOmH1G
0D0Y66wIYG+B7HkBQLRagxQ4mvdq5mdNeRai6zTF9KR8IXqQieiKl8bGBjXIpEQTAxoMUMgSJ3Xv
7C5Qi4o+6UhOppq1UiD4rfoZKc+HWwQKtC/xS54pUIQ+d4EMvzvzJmtGa51S6x3MludhMgR62Bv5
6iqFiPIzIk9v5TGmT1iE1izVBaW+LTKBOskonvOO2cWkpVuz+umbCdi2Vkn5CRobaTPU7UiqyhQZ
SgPSSizWYsY5vznyGzWDHBITZoCK24k696zu3IxDrcmBa56zdB1vBzZtZZToJb6Ey+6yaMmbEeT9
BkmVX0Zwf6cJkcuVirpRuuUUwn/Yi9qpjRKIku6BAVntX34j/8zzr7+xAGKaUhM4C20oSS8bq1Am
zwbnaecDyJ2qxQ2ONFEY7tK7qwnGy43DQIac6m3oRxJZocUchI3API61yZTy3/axB+i1HjJDLo5Q
bDT2ymYZfJPN/UbADR2rAZQiviNRQagEQvzJqx33aSOTBBQHPYKZAbtqzEDNap+BhITuM1TU7yKy
SRBan3rfy1GYe1KioasOgQK51C6Cz5MiktP90Q0wHohHd10HoQehS78Tu1PtCff6IQOSY8/aV67y
0bvayeadGvqP82P00c0J7Z52RIxXaTYr9wqsPqL96T2ysLDa+ra/0NcbZWwVUGP+Nu2saHmqSv+o
cXhsxRZGiv9pbVhmf6tQgYAWLpRg2uJh0Y18Lk3/GwFZapozoKdSdX0CgDPfatQkrsQ+7w7IxlGn
3uSZyB/Odq6OduE8pCOMUr1qt4QHAEmdnQrub7L3NfpCAikna+uMtK5AEghBUoNR+RpW7GkOqtis
prtqsjb2KzFmfoVqKhEqCx1KJF88EkmqenOXeDfxGSiJZMdu3B25KAxfvf1p0k21vE/s4llRalaI
Htr7m343MV13xKUFnYh/vsGfnX8aEBReS4QKu050vLQMMM2iDB1YGYU7XdM1IILH8p6XJ7UrWLQA
nGythSkmPrseBZLh4eBLysMCnmv3KYHPD1NkqkPMxjxdipQ8xX+0tzWvIxINPFct3nPUV2hSXSOG
rKddOioNsX731oT8kXNZ3WnMsImY8CYm82qkyZHvvl2i+cPRYcHDSX1+bcSFqpph95q2Ocp9p/Dq
uIRz+rtVJ5ayu68ap6/y/w45qv8FwEF86pQgD2Vwe4E5Ns2DoxI2FCOyLjWfCYXuqcxCnLJ3Yli8
nCAOXpSNetc0tIRMTSCFe0ipkKveRmfkWo2Jf3XvuZilYQCffs+7bPWdaFWA5JEQ8npQBkPIxuk5
ByucFNaIggYVzWi5lcenusTQbLQoxqY1KwZp+wa1FSw67WIznMVqqRhsEVyq3wOeCW6sgzVoVvPW
alzuLkXActtWg6SgYSZ1EpuOiB/aOgUQwkSWuEdPTTPa0j+V3nubN8v96NWduGIoLsHwVSBcCfhL
D57A/ArRXs5Wsx0dUy7/x2inabBJS8PhKCvJ7qMsHj/DfY/4wowHK7LSmlchvrlUpeE0xRZLZEVX
/VyjW7+M1e3NOxFqiGkOnrIJMfjCAHtYAWwXDNkBMFlNLlnayzqvsb5o6A4YY5I0Zx8cIeEKr9DM
WGFmt/oV76/1KXWWismpw6mQvsGj4sSj2XRROllZkviu2SfmTioGwk9PuqEV3h46rrI87Kuc++3G
vNJP32ZJ6L5SuRPd+rmdpL3kZKesYQN7uYkv73CmoqdFRFNCjawDPbCiGIUfZTnlu5maunmUBix8
5nxXg0H6k0opDzot9vGxqqVLIxHbQKKjf1wn4A0c6nOui3o5s5FSA6/gUo7H+hmmqtm1WOyoNFHy
lknA5P9QVK5JvDFH3aQm3ysMf9V+J3gk8SWqvQCkGA007Ze9QJ9H/1EZJyHr8GFuXGnGwil/ZpQ0
I26F/Gg6ReICrs6Wx50TwUM8oAymeIq4qStLOvqCLFLwZaOqZVITtbhdezZI+TisMZcaEpgn0/hr
2YBczE1iHxOq6TuXl4eg66cbgVtf42Snl8G33SnV4FwBawGOsjlUHdDoKjCEkSIps5eqSdPMih+w
JvIiwLqUbU59VENMi7OAvJWBLkUh7SoLaSfeArkHYLsuGWtRmnKWPYJMDaR4zA6sX+sP4wlDCxoW
Fij+OV5y3QSczM72N0NIy9+5ncISLmjV+jzqEkNImXcDCo+6vIH8gbqb9PJ08eZNGNGZcrW+YqBY
JG3HVxAwWoE/s5oU2/bZ0hD21Qklqny7PuKao+Eu3/iYdHGGDxO/9DPY31WiRH9aD7XJDZqW7OK6
GuXDu9qHV4tpbyd6u8OxCu9g+3s4zrH/lyPPO4qIqLXkpNK7+coENgYTuIXKqfN4yWZr1H3E7ipn
Z5JsY1msyW25eCXLeI8cP4z1zSrY5TinqQ1ofyEPvWfA+/P/PdilOSGkYUfXtORHjzHs5/QcF9Gu
LUafVTHeSaBjNVf25nDDYgV15u5Y0Isbm/Zl0YEFcsmqQKm6iVmlfDdBYfVLm6TsOZoOZlTw5upC
RBpy7G1oree/Ngl6iN16tYmfoV13SNphpuwV3dCl3RCpSkai6Y0vIcpmRqe0lT15n/bnLYr2jHL0
GH5KcQGoFM0w1s1zLuWzrbMBFMdXzprgcEZERphF/EYI15+UERXXqAUEA/yR7fsAPqd+2W6eY0Lw
6fSZMhV9C7/65r1GRiaqeldZrbien+e7m0B4Ve8XUQL7su+nPO/Nhk9+4+f9gkTn0Y9UFZoNsMGG
mK5g5FN91wIUfXCtRrdAEKoSEeJcbPZ4Ip78SQSOLMAdQlWR+UBMDM9nfjaHp6iz6YaZ92kom484
SyJqa38REVi2LpFNP4ddzLGDl6l7Uj4AQxXC5/pi112Gi9pGWtCMaHGcY+rDVKJLpyNY+M0pOM76
AtJjs0ubqMongDdUT3dGlJ7r0H5/Blnke4Fi0mUQNX7FYu39Br1vH1hQ6vDD6e+ykbLw103k2n5M
p/PuKFv1J3tKfJe5YwX7oRhgzrLrBgRZm4Vsd4vwYsgkfcs/O7b44yFjbO1K/AEtutZRcxzML+6C
gpBTR5Xxnm73uP6e85WJOytwnZ/Hwfj9jl461TaBw3wObQK8NGI7EYhmLJvhjzTbsEHYgpG2gV2O
ogkqGU6a++cuO3pBvt+o42sH4oiLso7UZf9W+K6cbwQG6fqKWQRkdTQRvkEMl/syYpoq7hxldhmG
Kpy7TPnp9sYI+3kv9tP/N/yrI26MBiFrUtUNG6fbWA6aLM2VMT919nP3iorXTxQZ0bGIiGUITXkq
uTGcA1MiQkBI+NP3m4f/U1e1i+Xb/LqWvYeNoT5W/nJu6Qk2mkX2RDzIpuQz4zQ1jki37+P6YOjS
L7k4ojic3hECDAnWDbdC9M8Qxc5LFrtqLK8ziXYZPWohvIgggthB4tWPcYexLUV0ymCTEj2vUUy4
1pQcTF+CprayjpDCjEbT3xg4GThNBp1K9P1MBHIjYZuf8e1w+WwJdjKJRTwUVPaw5NogwtnVPPEb
04RqsceF4AlwRh7VivebxaDK2h2rrIQO+5/F/34gpfOSnMeXEFo41urNqbccnbCp2Biw2BwSGykf
7tsGQDSJKSPL6Iz/LXj4SVsT3VVX5N7IVlUtdc20q4dAghGKSZ0LhBCTT7Z74XO8RELKOUY3umox
HkldFXh0UB/6+fH9MRd0eubt53G0gi3U+b5kW2eM/Fx8ViJCmDrCtRNMogbWbF8qOXPF+oCWsqLb
XNpG5ZzB7qh/oRWtF5J0N7K9iXfr+62Vktxo1V4ZkzJiJJhLZ1JY8Gh4igwFInK7ZdwMfXDTBKSh
eHlr06g9+r0bgQ1Poi/pjAkL/GzFfl4XV9Ci3bAbapELe5hSD8toFK9Ck6zp7WK/7OrjWcJxBK/r
i1aqhcKr0CAIhqkwdcUgh5Y450/qjjT9aAdsX6fTlvUMgRkwkrltuC0t/hBKfWWRk6mfzWrxsbTF
G2NwKPJzmyCZC588KBswLGojKlM15ZcphuBR3ZE8q+71ySDqAVIjmz8+RWWhdzpJnxHrjUX9cC0T
mAXFuCVH/e7KSA67yqwRlbUXHtYA0UBZIO+x7CUPhZ0dOJt7vShXcCZc4572B/GbTcY7iJwDcmmX
xtp9Znh/eS/yvwmDwO9aOwEzlbmf04CxGhst8bcNFvYQ6H28vUzTr3icVzDnd5VWst3USk8gMeN5
Bu+X+c5GY0ZiJMaQFBZUZxYLUoLanRE+njA78npcZim1+HuXkMfbOYB9oaJBxR6Ybkswj7vRyGBY
uMYYqIy7glN8f0MhSiL2YO9mJHWK6X+ZABwt4rnCaF0/tLnXHIgd4sBbKEgRnq/86z5vTBcmN/Tu
YcUpbCoOyXKW1OpG08pKRNqC+JmbrMlrIIMpAt8lB6XBziU2XQAHK5FXtu90PRvK4xNUxepx6FWZ
xIBTeC7jlnFTFxWTRRLY1MTlRgqfV+WAcRUXKFx+YvCj9K9bM73sk8WrTyb/DDmsAifv6heKvHQe
9Qanky1E+hn8HubDzZVoivuyQbUjnjJ14/yCofNsOXreeNemwWEVaBVyLfxIQaSL8OGOG+jV6K0E
gGvekAPnsHLOIxwHiL95j7zOXSwFmlcskZBbmuzQYhj8iV3OQ4INLf8Ft4AV9FpcWdI+8zsBWEE7
YdLe3clY/ljrrJ0h/T6bA+JcE6azRAcgfXO+FaUJbU3XqjITgUAQWh7v2PzImrsdbAwUtxwilVQG
mM6q3NjEjplL5RZ3gb/UsO2noSUhrYipatvq0DrmRriMlF0WC6qNaowqfGyifZyA85O8pJEVu00G
yGNCXzKH6GrXeSY7cp+QeDIqpyfR4/ZDkRzytRW93PgFsZtNA7b6AigovH5TUKjvWliHJcoPtSQu
1SalM29yn7aZy/p4eq+47zl76ZXfj7Bbf2j0KZ67XdEW0Xm3UGon4FRKh4VTH6ciszBXVfcj0k9g
3jiV0xf4HxKE7UsQVeQ2wIeRtqCzxieX/9qNeZ7dS7BMOe6O8uNSDcdtC/32gmSz2yx1I6D7ry8q
lP9ibQnjRXBihYIfaVw+Ku1a166VWrjwhVi3sRfJmDQz+pRjyQjJmuvJahMiU2o3V6COewHiZeY0
fU3BQAJ6Fbmt6JejcCMlW+zLMAq4vqV6EnFAmWeRgkubZy7m2Fu+LTYGQnuOcG6bDUmRpg9UG8fu
AfyYZRI0vTxK0bRc8kcZ7OoghpC3tiDeT1+x8dPhp9TDlCgBf/Fjdii2PlNDYHPyQx8Rlezgd9Qn
NjRBGtf5ILMNPdt06oSb07WDxVGMmkvuz5GMoUfpIFgkc+JSqK3YPGYWIZfUj5PezhenTd72SZcu
Uql+Pz9t+mjFyI+5tp7FtWwsp84PLeetG/u+GviWA7Rp00YuK0hUWt3imN9Wl8fjZ0zbizGlqW4P
RleuIR5XPyuQfKdrP9ecVJYuer5rKD3hrJYEWHG1AZCRzLS8mmT9QoeBeW9TgONQpnEtqDHQ8x/Q
13Wk6KP3A1qxYzjh9L9JXi3AQkjcuYCRAeCUeuJaPfyHf5Zv7NKkoLa25Ios+J0zVC7JI3VQBQrU
5h+O0Kcm3Vha6Aj4qICo6D35UOs3rQZlhRx20Rdvv7pp7CUGluTV/a8GXXgobGwdMthR17EFoHxx
3LP8axg8QDPJTI5XUglgB6eLG0426D/Ko2TFfbKhzef7S4pubsUPA1w7zHojph5QdwgaKzphWjvE
7B+y5Pq9GYxShy8T1wHHCfaKXp9OFjAMN2IU20NNqtvfRRZEqciEN+ry0Q4L52Mw3/k2t1KkBKoA
ChSLAYr/m30YJ1y8C2djA9J3u0kb/kdhXRgeQhlDyrdVSwlayhYAjHfGxLsxZqhaMLBXP81aBI2n
AyPPjJS9bJAQGB4EoiBaGvjgTpt7bSr4nsH+VINl2kLsJAHf60Fs5j9CkLMPHFeHB2tWINCEwztT
4dx24XwAZhkAmEthvp/pRDdR8f07jTaU9ilxOmwNIhAAkbioC+VEKY9waMXsiZejLftV8gcGVrap
KTGIBu6ys5gCkNEbyse1Ct8wx/P+h5sdZEDalXVWQ7B91LQF7G0KQYx7ArDilCgqiJ8dUzVIxGUU
y0HMzsj8vO/plT5Ctwm3zwd/VM2DS8EV+SX8Bjccw2PqYT1QrlgJYfU+cFOJY0yuxLE+cJCqtYfO
jpaHV0IqJkZVdET4ljJ0fSVwavmy3uqqSpZIbZFoeuNH8bH1Ge4qA7PO/7N/ZsdhwX08QUlorBMd
NETPNV8Zg5diI+1q+3fjMMZMXrdl9H5WZo6VuPSKZZhTHit8aaA4Fk2MPZzpWhtChVK1aI7dmKiu
oPEiaMqXJapPRFyEXuln6Xg42OEYwii9RUUhVZwJ1R8hA4Fd8Hm2l2VUZs7BI3a6qL0e3XIrkdW9
dRKi3LCHc9n6g8c+8J8yqLFx/xHaNwdOhEF1NmB48kT5RXMqV2zF2yt5psfoyI+d1pMlFrhxes4q
4ZA8BSTpKyFroVoRLwmoeEa1KLXzggTpTk5WHvcOLb010bUi/Xnn13b8e3asKkhSguXAcpwU3oQ1
VNXYjMZ3JorVhVmrgr54Q2mMw3sIkNzIelIgonYwVsofZheTlm97cQ7wAMQADnfhdm6BLifr+EoT
QqYXQ6tVo222fKdvrkFF5vFSbIM0ssq4NznnmTvoJr73YNwCn5i11OAK3sBkoLBNQLhjiidRPlrw
6/MppM6dYt2QGfN3qhxzQmB52Jsq9LghDOob5fLsMoHYhH+BHjvhhH2CZjnA84i0Z33cjMdWN1d0
IV5Y0g7/lXHiReFM+4kahh3XJqlg+asp5lKxFRhUVX51vJ0uq2RV6Z6gkovyJglYgDK2oY3eVBIu
lt53NbjdSDjwQbE3sJiPW0v3eb0Ec027XxaFn5Km3P58AZFQex/lbefBrliwq9zydGCk3aTSPze3
JuRyxckkCTRehb7mzUka5/d31r0BPwAVZwRklN5sXQ/ri/XWw8tC5JBOuTssCvCH4MvpmBjQ5Knq
eSSkhPzW5E2Ciyw2agqa6UJsqw9rTqz0wIObtyZA1tL1Cr5oDmXWAo7CirANTSCdqxGUfKBr6ndd
ymE3AxzjPEH2JpbQT50LVH8HychaBeBSrAUc3bMoaLiSEKUW2mCui6GubxCx9S5Z8CSjbH7eCimm
qfJEB+mzlOvo2XAye3dfZn9qfA+fd74hlqmg5txc3FLm8NS5lzKI/pzXHwL6YWXNf/3YoxAESesM
sykWD/5Zhr58Nk6BymCi9GxZdLk2ZmcFKeicEW8YH18YAQ6nCBeP+NfJoc1wF9g4Kfzl3iyjsSyz
MPl/Wq97/m5xBfP7z6Y8QRK38x8hT2VNeT8+xB0GNcMt59SYLWSxzPaJ+bTRCf1h0kclg8PvT3yt
6cqPKKGF2Mzu4TJ6D0wbGsOPHRxzxaSy0JkZvrWEcEz1jJ6hkWAuRAn6b4wev8j1muTMGw6pvFaD
8tJSvr7/+5j8PvGtbxxRdFoJm8W51dXWK861lZ/GYD7EUSD3dHZr4dU81tkf9QXHngkc2GmjoSwo
GUB1xmItEboigJVDlDoU7IXI7vLU0LsAXlFuh5vD2H0SL9HVR4ocITkIf+0QW3JmMgmbM5EA0GYl
HeYeBnuL4BwgLx6/yPldEmDdEPI3sNnvMILXCeoeh+V6gTZ4eoggDmhjC/cOR1WBq5h/LMihMzSd
8/Lnlye2Vkn2NDmZ+/Qq3DnCpG7M5RTKTtDqDdQ7F7Cc3t+UabWVlbzivUYuVtaAcce13AusQa6a
4YVytntHWCKYMa4otnpc5SlXOsrO1FV57tq5wzsvHhvgxQEGh7vxWZTXk3DVCQsVkuXKD6PX/M6B
4nKjmoYoyGlE0siC+7iqKwvjXlBEUclCrXqp1yt726w4SIATBvRMYb0lO+dR2ycKbdF8M+8MPvD2
SySXC3FCHNM5UITNtBZJNYGZkh3gLvmiviw9B7Grnb36OiTZpadHI2MvjpovW6KuuoZoQER9IiJ1
ockl4JEbBFG3CL0mH9Mf+FplofxP+1Km1nFgId/mUt+dYyMruLFeLzNqb72XiPkQLGvVfj7hYBIW
/9eNsO/QKoulqu57fraWg866x38vVw1MGQmBK8V0cFFBh5UDsYclzn3DDhEai7MQjy/NFFMEDCNJ
t8M4apGrIH9Hzm9E5DCtpaXgpkCd1IOUjagKwY1oBO1koafHA+ypPDyuvHI1Wm9p/x932b2BO/uv
/TXBAphKo7b3TbuEXjgsjjBXOMGkMMPPMjWDeTRNYinFdJ2ujdwsqfXNypoMMTjPGbMwXsKkv/oS
yB5xh1ilM2PAmZpAkqB8wHVncP+Bt2c/epRn6qGKde+4Uf2tUb72pCycwmm7lBEtTDuopj8gItuB
oDRATz5xwhXzzW/A04KbLz2ULdIq+nT+pD4lU/GYlCymkX5eV1pmwaDAn6yj4l5R97CjQiF5qIz/
CKTjshTr3VSk8RgjSja+2tRYuhRT3PFvdud6t3tnRzeCxWXaSqLbQl05qUik5KMfQlqW8z6Ew2NZ
NfjR8TGSU1IrUdqNEKKDoA8mbc5I4tFzw/u1KVZG+yv+RT298FrUY9p4ltUm9+mWPj/JjqCzZU8o
zj74mL+PwfShs6eJcjjBI47VWCH+pku4PNcHH590zojbb/XluoflkR/3WgxvIj9iBejfMqWEzUmD
mVuv45VpSIe0NEhbek4t2ZQDgQeoDA70553AtFcozhS7rT9Rg1II6dDa8lkWBRQHD4veagl6tXC7
aP63yUpEi0H4sBdgvuFZAIMhQ0KZ1N3I+dzr6jKsN291n0X8S2HngsXGEM5NoD+L7pIuEJ7Qswnx
9SWRAWIqcFYh0e39dEwfNycc+syy6L5CJx+SKFkgA/ZeJz1cEUSHeyoqYwBl5gIumY+EXpi+K1b7
N+oEaSp+knRirjCk51rL/fbPJ7AsEQrIt1iUhB1GFmSMYwW7mel0tEHSQjQStfnTtEQs+gs0Y6YZ
sSNwtYmFDkc8+86SINO25IkjF5nfMfCX03aKec5qeistCN48M4yMjmls1iM4HDbikp3kl0xiAB4F
nIDqP5fGXDexwUcs+7VAyQKAJZC5U7RCO2gGNxxmKuTduM5GMF96l6rM9RA5hb5Vy9NWQ0KhR+IO
etvObXae2WsDSLpMramH695XRozNHUlzsfzjLljZIffKNv4KEChnyOehGmMUbTk4ZMTKAsiyTK1C
GLg6b87Z2IOFnhP8yg6D3e/0aNpUIHfQCNCJzQSr1v8X9o8kNliPUdD/+tc0kEfng6JXeDr0yu4a
yQ2vG9JHEnc97z6+IxjLmO6Bc5KfriWAQS2CpgM/eNj0EtQ9hWMnO49lbeFzL6xuhCR/J6PYhc93
+zcxqTYQ+u++dY+0Hv8cPDDPbCUiIbOgZ+r2dhHWop8d0R11QSZZQVO/KD72LkiU/gCHKxrzEYqx
vsAcq7stb3hC3P3bHLm3s6WqzKGvkYHlx9fnq3SnsP/awoEU6GYHpkLK3Ec9JMrTv07AHfXokBjU
WIUTpghjMhVEK6YFFxBe70MvS20ZDKinoQrBWO69M4BeX/pHby6kPMmsXnZf3SOVirnW2FnPABUb
lI0o4vYjCtdL8qWpZs+whn6GDTW46BGi4HrddBlldrqs67p6bMRNChXiI3tYbnffA5r8MffynT3y
tugH1C9bUmLaXsHsgbxUdh+Ay+jXbXSu5eY2S1edp81WEqHr59DfHkn848Mk/a0bGX/oUIkk40Pk
uWPHJz7LQDzpcCuMkRQ/JMb5Fxx3PaBiQqPXI4URuAWd11QpbT1mP+jLj4RL+c86GB1FTdTs8tfl
HGDPaXaw25sD1UB0TpXD5NvfYzzKnsMQEnQyByX5mjVVTpEOrcH0RCV33xKUmjsH16js4pmevdcF
sxnkVl8rE2/wPqXMv4ptwJqVVVnksmizj7MPyfKO105sYntP9qNjbVDR9m17Cd7TPY0F0n9c7fyq
xAmthLsL8Y23Id7kJPDA216FME9H/IAiVodVg84Pw9FrEKTK3CababGB5fhxsUJ1OpWxESnzY0k6
kz3kLeO5noiLAWIZvYI65tHnil+4dP7Ef1QMGlhyYeRqjSWC6YUbHsBA//evNk1YdsPM8LjY/1HV
qGld737vHDgKPOEEHPyNsB519DReQJxezva1Po9hvLbpmQzu60OrCo1YIIHWnNEZl7E4VFF8tNeL
nTrqX1++++lEmuIV5fELwuIc/j65QhPbDyxw0lrQJZiUz/Wz/9b5hCXtwxHYOtAiYuBUfGiRk/ae
kg7u1CSgZX/n566Wd8/2BqTqsKMOWFNJiSYIZcLvFyAiR4NDNgBdDClcLBXZB56s64j+IrpAJp3E
XTRSSNFfucaZXIUFetNds4D5dTYmBhdelS34+inZUqh7Flo9G8uF7GrhMm4z7Ie8kd6j+AURr3BW
1EGLuc707D3BXMPdRI15hXL+pS2MQkAFW0dnncH19qNp02weXl9HgaN//sa5dL8oSzZ5Wy0Id+9+
aEvn7Z0tAuDGFhDyxTYmZRKZG81O/Nlb7HWh4ymuEpApGTvKqTwBXEkL8JeO8pWjDllf9kx/QFzs
U1nER6PCYyy6/8Upix2ZVFORLd9HDVcMrbv/PgxoCJOdG0MTT7ailV+beqCYFcq/zNJKAkfNEdhR
Te5voVRtXCjCENynzRG2J9kEX1hyxUk2MGtnSFYqAqb9ulCpCu6PpSbI4VI5paAQwPiWEvAs130f
tJh+1OxAtKD4WC15rimIcYUlA6BGqopv1sDB3TL2qt0hrHaUijpFQENqPAgWstKUN3HA4NOkaZVp
lkxnFJdNmx/QcnZbptA/DQ0V97WHvK2rACmgnlAguvkgHz3rhROwYJWHDu5Pt1UlF6fxX0A5wcka
NkrzcCZnbIRyC4UeDEVbIiYTlFkbWQ3+ueL0+7hJszKlFbuDdmMKu0M649sHUHENw1/gUCbxjs4W
7DOhAtMNxMs62UUERMisljDIn3yZ5YXzhbtfvFtPWlyNxhMC3Vv7K3XXLAIKKHqlMyCHFmNW9bFy
n09jXIxy7rVuf+SpfhzJ+7XPJe9MhsizE5EvzyuewyL79yoneCQEATlJiqeVu1D6J4dL0msoWrRA
ZgQy3AA0tF4VUxcBrQKw7itmUquabHdjAxIHGV4AjnqMa3B1o8V3KM+YbR4Ov4EE8+fVlWr2KslS
EfhaKBSUUEP9RrJFHVnU4oI5k43a5ftW+A8lAABBBJeIAR+c7XS6z83M3I9LmdSjmvtALvo1R6gK
p7iXHBFPpkerpDfse4xORWA6DN/3m1yXmbLHS1XjmraQ9ZEj5TqF7qWFRp7ppDEKAGFWBqPctZOh
+wwW0/925lZGe5q9NElj9P5siAFRwTkMFmhYLsf2cPLof1ITtxqC8ioxFQaSPwFt0I7j4q47NlGS
pRINz1I+ubaJ/2rpIzF4XQp+XLsvdH//04OLon/0GguSsZlQZ4RKDLHDi0XOArhdh7y+x4gF+QDa
3iSBcF5r1fwV6Wbh7oOTSy477W0XwU0fXClSoyhSKmYiaq+5lbKz052LSUnpyIxQVqDc5IjGAAY7
AMiuYFe+kx7cmVLJCKhwLMeAGxVkIWJpjMq7pumA1BxqYwJJytz9HyTmYx3Uhwjc9sSgHCHlp7Zq
NDGkPoo0exJ2H25mv6oKQdznZPN/NtNZHWV2/aoayNMuNP0XlWHzhBf5bSBOzk0GsFniyCKu0c46
GNNBBSM9LQdtntehxBNQwCKt2I+7Blh0wKPgsNGQ+KQ6W3oH1HYOfc8To8OoswMamucSZWL0ZLU1
SAzMXrFc3HPa/LMK83lfKu+UgCc55ERZL6LohQfJdVFubMZwU5P/HJ2rp2O/2kQzBxixtTzDw+7v
5kwbfbGl4ZHP/tMcoFgUR2xEWXaagJCwKEbNpeJ/UHEvo9lGPcNgaq8QuqUvzHYhp1oL8+y7+phc
uBpkJFOB/IRtlhtAtRS1VNvwE6/JhDzq9F8RWSMKgCwZSeJOjFvCdQBx86Ta1sw8bCGYXWWYyBH0
KvmBzKAH7PaYhhFdJoQMMaXW1kkVGttBYtfS4Db2Hj0976aAIrQEu/OE5bWBK5K320QVV6uko/QT
b+lJhdhi3K8KK5bw/u965OxkLizKAgsik12WiX6OFL9rUa7UHL++kjhU70Hh5s78OIzIDjHNBihz
GgYu2Y/HLyuhXGV09VhWTZeyGwmCzdm8CVvYjb8de2iOQLze2Wqb1KI9MPh23FnQUgaYGaGXn/m4
MCn9YvzhbHe9LIfrRzDnHRjWqS1wCULqDmRAswDfibNbh5rfVCb094KmUM0dBA6hfIM/xE+XTOZa
yuHxJgHwE5SvDhdUCgC6YpIKT4Zl1uzNy6hGhVj3OZgLNtWz+SeoPKHuW/k7lOsuRmTiik/9HE8K
z5yBFzHXEr5fwJAQTrLIJGjqa/UK/s5PMTc8dLFphL5ocqgaH76/mjtzVDwDcJor/jUUUbFt8nIk
n5zzFk/TGa6p68b4FwSTflr7/iYx73GJngIMJxfOQnjfShaX6ErBrMAtW6evuMAG6H/rkshGiplK
SbbyFpyeiJbSxTUDtooROyTj8O/oDyvqz4LmPoFL3JdEYyZEsz9Yq1lTGB3jWrT6m1vU6PI6afH/
AM3NRnCXrb/UsuwDYd2jmJJxOq7L9IbRyNrWFcR/8OD1DKW8FH23v+S9dhlDfU1mp4YtWk44DChA
dnAWd9uLPmlhjv0jSlYIDDijZTIZR8oK/c5Pl9SlX1VMTxOKi7BwyXtwL1wC1SfNL/RfsclhC9OD
JlXQ2KmDR8QRIibDeiQAY8ATfXZGISnra5gWR3p39OESpzQ7E4IJdS2Pzfl9fQJlWriw6SekA0IF
pYoPgM/50GRexNnwkKBHskTdUNq6Gh9NcC0pG3j8ymGvwVJ6/jxBMzGi5TIUvcbXnyfLmbH1Ll3F
LeV6i4irF5S08vnlXziUZjy8OKiUumY4o/hdENx0J6tCPfyNiE6aNRczXjp+1UUnWcSY3VlN5GFm
Op2Jqz/1/f+Zr4K+SO1qel4dENBasILS4zD5nxm5Cl6wdB7a3EGZX+1c/CfFWZs4VowkYq73lacO
jMZo02OgjvqjBcXYYjsehUKPOe5k7sJ8DXq+roTMyD/+eYknAbYZIViIuMTFwHcX4gPXJyLovSYN
/UbFFOCfraWXmFm+fti4D0Y0Aq+Jhn70q6EV94JaB4kI9AMB8Rcm5ClnJYyDcQyduDaQNRnoP8Rg
o1AzgWc59Vap5hfCKA1+pr7mP6fbb2NdHPaTXKSKBWzcOVdAmBtpgYC/Qg1nBvx95v0sRtlC6B9T
yZxn4OhWh+XpXLpZhzkMw04ZZkPU5iCtfCL7Jv9FoQfic2JinNzotHZyEow6dVlPPT+GxJN44Yq4
IbT/qlSbS5Vt6nuKORxy/t0gSdvW2PG1fqIja/ovNPCt692fMobC8CScD962HVDQwfgN95vs6r70
2KnUGG0pwvGRe/M2QTJimmS0afx+hVCRAviCbw+GioP6ev1axJxuGpLVSfMtsU375NdaFKzEXagA
GnXV1p/K6s2dFU9x3UWoY8eWhenB/+Hk89yAG+nUyGpePV77RbaTKlcX1AEE9chxUJTzXukRwrme
cZS8oenjLWXUeniGKiyZpUVJ+dd0FevPnCfqvxhyjPvbTdodNl2jXXCZIQUFRX9VXxBixM5MI6Gb
w+JN56JYYK8+emPEuQKvY2Vpehb3djfhwhBo9NBE+k18eYQFqL8Pb0CbqFwvr46nFnA3qLfHMzsb
3h7df4uIh7/y6ADNegFLvq0qOaVw6nhU8rMrDYdJaVgor58+RUTsk/lVy8Qaf+4bLLo+LCh+Yt8J
6dNALNk2uguCeKoHLw30QjSbiakC12TVhZs25sOH+zZAY+B4Z4CUmes3B3N/nUxC3a3DfjvbRDQZ
JOi0xQ6qIO5+Nf2HRZSIfmdj4XOYadGkAQRRDRD8M7D2W2sO/lgWClxh82smoJ+8+N5az0Qusmzm
xmPqWEpONWZLzciB/612BPlQOk58QbEEXgEEJ+Ad1vYSOuxcFmobS4POphZwM34gdEQS9Mc6RkQW
dH6UkZoFKyFNFAk8tEleZynGDnRBtg60lh5tA8N9vwaenftG3L+Jd//I+VZafdPEryQOJUVlDzei
KSVnoegtSsLRxBkYHHxBc6NxvoOFDmm0dHSFyRnC6YKKCUf+3odiT7ox8XJWj0qyBfTaiwDCZF0L
dFoILrb59WKmp8Wc81MyIUXAUKmFhzptDBr7jj2kx31EeCKG1kyWXuF1IjpZTuJ8kZXE1Uv8JUld
5RoJvQO0X+bCAake0M5dAYOvjynHzjklW1JFkWKGm0p1wFqjztwXhCzmyK3DhOED1GsSgKKYcQcD
sNw0IdwuNRXFN7wupiqEg7v5Ek7twlK8uEa27L2RHUyri4FupDas8Fv2a3KYG+CAjEMBTe8LdH2U
OXsmV25FQ6wguFw9tbcTbXc8ewKzMZzja3SRSvQ9k2E/edbeW0Bj8emJgL3+f0i99GZVlpuGwm2s
ZwxP4N+ugjgIZYPbgRnpUkkTVOlpkNeJaxFYk32Ugvw7ETD18DjyMD2uvMznPxCNV8DTNkk1hzM8
tJcMArcBV5rUG7Dvia8eS6vMwDfGhKv+pqXa/RqOxu/Yjl4hBKPSgGPoxmro9rdFPd6VPVzjW1aF
GdOwYhpjwWJ0M8/55D9Bs8BzTbTgTsgR5Ea0m3/zr87EDhRpz8xh8tKte0C0ATrnyNkM80i7374w
nsb4sVl6Erg9vUn5r3dsx3UeUsD+mCuuWJHzulfbrN7I6NfRjKoyOEWgZNAtkEeDbpjO3nqW9iXx
SnS97M9JrOE9G7vNTV53nbNxHCLXc/wzPpvENT8MfTw2G4CKwQN29Q5ONnvO0Cs1ZnpllL+bqe9s
RFoAcZWGHnWlFZ8xBsj0whnKcYot5up1siyc2vbmcLz8qJJqX7xSl0rhq5Ea7RSxfIjD8Tqr7i2o
uGKO7qyaH8MtuqSWsfxSTu4ojjJaOlIjO3A/GJZqk7n7rL1ITEZ5aKKKSFIj4SS72BXMcHZCna/j
RZeL6k5uaXFdqNTz23UN/m6phvMrEQObxhnNVgyJomZ+40UXWG3Zwfz5rtaGxP025jQOr4o+OIbi
DSjLSQSf4fGLCp1OKA0Ax+jOifFdfe7Fh8Zp1kB4p8vl8D1vF5b11o/fG25X0Gnmp7CKziHAKLZ7
TS2ieUMwzga2Q5JnP+qn9TjQIg8kzrXZk70d0YtmdfbDfiDtMFjOqSHPsvJmuVTIR9dVXL4oEFsJ
RAVZxgJxkMBHjJEv+qTasB7tY96fF9OONUDYbAF8vMDmS5UoLyk9/Ugo2/AxmXXkyaIs74betVo6
HImJ2xomilBfHteuELEIcGYK/1l7dgyGd2+4CGzhJcNcKgAxOlWyAlSO5VruAmQGyMuQSd+Kvq5e
y+EursIMLu3CqSHoCeQqMbWTyM/CqiLtX0ssfOQ5pt1y5zu0tZrT0lTuoRHO5bnGbAUdVDMTr5F7
nB1OWEeisFTKnuD9HOsIGvCM6j3A19N3bL5MPmWlgRnRXg3Auss+GQ6USLLd4cILLkyfvC+kYFZv
JX8ZyqBXq2GbR+zSRrX02jx0znlEzmexa7xjutvJnENj9P4StcWHpPK9comhsNaOmXvKHk+lXiTJ
49zz/4YpQubuYcfu6A6bU6N4/k6DPuKNMQf5xGHJoaXT6RZ+vNtczSdIFjHglcKmHhz+VEB4xRCG
gtd8hmejUbLWRpA+S5/divatsotzWbySGiH0O2ZpHOVSWgpB1E4/11acoVq2n52r0E36BaoJK4O9
W3ELK+7k2RtKQltuhORy8f6s2Xv1hcF7Cb1VT9bZpku4nMXD9ZKr08LsZAoh5XeuhO6VcBOqn8Ih
tLcDvAjpTHtZW1lYHaB7Mt8UmC1W61DbcChx8ApHsrx4IHipAlXx/KTMAx/zH/qY9pTnF3Jh9IE6
Q0ovocfEeALBEn+pYKKO3LtMxcOXlU2m7EQ3EbPSonnyyFzCwJP3BvsukJwDgqOfwrD4Scz2jTgN
yMtJaTeuIArf9KljEvKScf7/FBGk29/kWuddJVTNMsVAl5Xq6X4zxDvUf+A8D4r5kbKSM7POBuRu
vWjc1pxPSi2zoPBeLTeWqMtpr+erS8+JqN3I9vZRMAFDdoBjk1ptRfj73dWeeV3KpMHQA9T7Fs5W
a2Al1fnQYJl/mbjtutE+Rh3Yi1u5oP3RexLTrb1nAuYPsj+MEt7Cg+mumHJ57vMASHWbG+cctb0d
ltxjpchrOf0OiHghLQRi1SfF+n/nMtyW7RDoBIGYImmc0JUu/qf+ck4EIuNkp/ltlJcu9u/+rR8C
bpUTLLgIaWwbhv0/sz6OplyXqWX1Q0Iw9q/qNYNFG6DnQb1uSl2qJy2WYT3Qa3I7O/rSPXk5naly
+FlO92XcLEkLIyGFKihsHkZt2sywDHBepm2zaBn/zeTlg8R36Td35F2Bo1wygkoU92JLAQl0Sh4h
3CMD53hMt87LvIHpDyo3PozfRH7pt0hl28ShhF05RXiYDMDKHURbYXWyJQmNLNzt3aQb847WGjVb
1Z3wj+vt/B33HkXpKWU8A4ScTONpgTUYtyc9BVg9qh8/XJqjQB7VNHFcxm54yVR6dBHeUzNigXpM
siDUIrY3ot3K4SBdV/JeBtG8gfCae0XLtLerLrpmC/zsTTNZk7CU/GCRNNy7O4TEEmbERZMtdiRL
2mus4anaJXeADE0eg0hMxlkj0jiRl3QInKTUlEknu5DtWYIyTdnk+Naokb1ijolzbHOTawMq1Ubp
vc1enYCoJtFiIBilVdq/O0uwfbprSCaGakKNYYV/Uhxo25dwuKVSRwqXLv4ngG4ou7Ke5s0bqX4T
bMBAamZwBRYDRGsK8b3qoYWbsnD297SVNBGggxqhSZbtih189Js8gfRLE4+cMnbspBEUlJOUVL1G
qNK5G7YjJUqX5QZ9YlMCXUK8UrcxZOnzDwU8+hf423h9//7Z8xgvNN6ljqhlG+huHRe7wE9x0mue
GjSr+WAPtoikm/Rb39ljT1vbNaCO0swdYmhsuVz7e1HSMQYO59ueafrNdJ+QVjjXdfOvfIxQUwLZ
17GoM/cViWO18puyejF450/SdTH3mVRJZP99zHYd56k+0nLQMt5wq/9figUknrJ7tYxw5N2PQvv/
t3hSyahHh8ELY5tMLBNwf0YhHDIh3x87AriPHcDxbtjlQuPPuSX8nc5DWVHCLtuH7QX4yGOATkX8
qse6JkinJpoNWjXrhOrspYpSwxwpQ9ACEfdcfSXZ4hFqMCNPK/cbpXjyw60IWKwsF7wg2FtmZu3/
2UBl03B00yRy2pkYUur65ax0CuU+WNUqwhccFSAwyi0g0qXKwSkHsxJv3N3PHHo4T7U8k6eHCy+6
VErw6jLo98FiKcmAVHXD3i6qIlMb6FK88r1Nr9iSqHA2MiMM6BXxmbDFMy3Tbh9VJOEdrphcEO5g
4qImJjeluEFJX3/S4OPMH86arIyeMcQotf5P3/UK4k9ULeAnYKzVNdf5CFwAqjrDcynnTYTJgREf
uRTtabRtiUezELkrIU8dz1GeieV0YZpNJRJ8cteZZkbmuXBJNzhzLGViwGq/AMSw/Tf1SLqPzen3
R2zzsUay7E5e833F/lDWTc6aZstiHFPfaAimw7YaCE/TXp6eUQw0l/afqxPfuBAe4hjhqi8aab8M
obgAqnTbbNReQh00HS/2THiA9WnbSl5Avx4S38ztmya3ULXM+vvIOhHINJiILoRyvoL2LEifhWmj
ul8dgHHFRwgvijiyGxQtkp+iOSAzwygoQTnDxDJFbZXZKA2siltgQqC5/aagnxYH9VV7DZnTFx7f
iYdLe+rxj15dkQHoh+gPLqKdm3Ej0oiG6REMyHUGTiDRKZsPi91RCOeR9tlJIQW1Fhx1666KYpXx
q9kO8pc3b4eYJNNLNdGmZc0qzJceVBxUVKxMMn0O4FLOJ6r9228Z5Xo3qNqNqDkdV+2FP6xzIAGA
sB6DbreIsAgSS4uljTkqvEGVCW0ti4TAI6lH9s0XOsF48R0PWun3CZWD286MRQMcT5xCHJ4J3og1
SXUor043QWIBrEsyIQAkm8doU6dc0cOGtMR0ePnk6hIxrVX/zyU0shaQ5d9J9kA6+0OAAnBizaUl
947+eiZQMdPxu2/rCTivu9QfrQNmRoBpTMfgcawDL7R57XQKA1/jUSa0WTZRGCUNbig9qdJDesuc
KBEP9NVTybteMufyKL1F3RMsIQ7umJZNCkfUCeP5oOcuNoNuxxYbTifdvnAtbxtBkSTjnJ6ntkSp
7Xucu8/jTsBjdK5vwGaF0010ROFUes/s4U55aM8eF9dLAQfjjvLHRcPvEklEoG66cJd9RiIL7PbV
ZW4pgdO057DDc2nq0y/v1UpbP0drlXm6xuT30ami6RcGS7W1sbov/qBw7CLUHoBn4WmFEeGuxv9D
d+fK4oq0+aR/l1w62VsW4+vveWWc7fTIzhOduxR0PkigfSUoRIIoyVFHwlv6PxyWO/KD9pTdR4SF
6tC4mwHzjIHU+SkRVY9Msp8lF3RIALKYJtSaElCCxGtq6/rvrA/oJtag/tkMCXTlDQJlz2m/kpp9
gDYKF8/kwoK3zx29cAeRhRllzgbLOImhJeZlZ9fUJmcQzAyhFCBxnHWkpw2NAqTm9tPQ0BcKylJR
9FGTBB5x6icpNMZ8fXuZhXZmU0erqcd9KV4Wlx9I94syXPxW8h72a2+MTN9Vn6751dB4+uFbpzkX
O+V2VPealuc/3FAn2fAa8nbs9hiRJ+/rXW4FxuuqF7PS5X6VSqVVABmFj9Uhd/8krUv6reneWlCG
fQ1x5K3ixZZupErOtIrbjsKhrxK2vSp4ZFcKEIomj5VASinyUPCGCexwSjgrxuv0Et5QcFvMOJ0L
N+/vijOiPHfhQaWLsA8E1GgVwPXbbYKW9b0lsNY9f9lAXB1QSaBRYl5OPdEmlMDZ1Ro450RL3HQD
sjGY0JejZyPU+H2G6S2wJuuKz2yZ/zEno7geOG+80m3G7hWg+2cgoRRPRv4TVBC9tdCIGiQlHK+8
LOc5hwXgZ1MWZ05FAPkfwSBVXXUjZ0x3g4dtBGdu4KLGdsrms5dJcUqPopHaRao0VzQd+m425m1p
7BGCl78GwkReqkSkqeOlF877Zn9mqB2sRWj3KMy4YOk0AhMjX6XUvO1stOga+ROXgMhXLwgRY3gn
5yY1+mLuN4uSMAY7GXiQQ4h4dolYHCw/vl88Cr/7ToowT3ndwh8R/+hvggLojpC44Jr1TMl/Tihy
dE4KBD+jzevtLhoEdgONzAPghHwrdmIfa8L7l1ve2dz/fCGC9tfkJFIp5jYOq2dGsxGvnIQGWWUX
XFfAqRBQgTPmUZfSf2JcYbnkDDLhRd8KaN1xmsY8RK6f3pXezLQ0M6wR3GWevSHoPDIwIzqHA/LM
Datcrpw+yEyc7Gq7amaNXalBytINiX/laj0GpU7QysNJ2g2bn/6Y9X9FPqPaBV7tE9uIJc+JcBJT
lcrWNyVsQYMt/DtYN52yWwB4iOgDsEc5erIly1B2KaTMqEhcW9xYRWdfCIH6Q4+2xbJJwniu/IpD
65b2Xa6WZ7PUQpMoBy9cQLlceyMFH4FSnkP2SgoLzzVio//lczQWITyjEKqNBuTqCi0UVymQ1AAt
oP4aTwAiNbYxkTDDyesqFzjT6gzkpj8mMiNjyZDlM5NvBYw8t4SM8o7uF0TR8M/2ikTA3SQfe1AP
H3tQdGhLKd6Cc2ACwlPKHZIXWzCFM6C6i9ZDMq7XlkMK5Sa3i/MaiovVBcpsZ2leQ4vL28iw/6ME
8Sm0x7TBify7FWYwJP316pYN/JIoWrJ9d3/QOVVvyGydFZhAsSkQq4vFXcp0wDdDKWN1ZKJZJ7/O
e6cxUywL/UNuwHHeVsIE1S+sGVC7BBS34PB7Rj/MEVEm9oPiXtR3b8/okQrDwxxlLvCwlw1dQO4r
xrYHtpFBUaVHU20ITa8iyXUn0AlgAI+wxOI4jGkTbmsm5XKWQgavrAt9yQcMtiNccBw9j7VK+UHA
ETCQ8QMrjqS2IYozkuxttcWwNcQ2r1lTAuV7qA8l7k5IrQkw8UQKgFKzeTsWRUCkY+raVEa1sU3y
MB683OHbxORAVuf7gKXtALhlQCqN7AqfxZdqCNanzqkvP7oZ9XMpJSmfc697JpKh7Tn+jTLROYYW
qkRH8QMN59ozVOQ5icDj4Wb+klN5ajVIN4JBZP2tctFf/iZefe1jXlh596qVKD8zhLSEnlrurg5k
C3yGG/3UuLTAex/ZV+AaFMzGuRjFGRq/2moSnGkfmlVyVHnO5JpuRwYOoOT8KcJD9FXoYWZPYndX
kDl7FoTl1S5kUA9SjU93SUXG2w0WzxX2XgjX8dcN5Li1LeLMaZmgMKN676tmQnEN95JSknSf5WSr
ozrllFv1EGtn4h5N7AbSfl1A4dXPpOlDSpn643hOH519SjFdO+1X/9G6s8VesxsMvNfBjbrSKC9a
8kjsh2Gj/cvwbUQh9KgQC8gj3dVAfGNWkbZOc2FOWJ3YAOfDLD4lYzfn/kb0VrYKCyn3B0EDL5/W
Cl278in5ZDDy8ovtkSJ2Bqdr8sTXlR02nuSG08pSyY6yzhHlKxde3excqb/yov6wo7YkYZIAliz0
vvp4i6dAb/zXe8LbQx1/c4Zpn1gKpe+FKRQRUsAEApmtcy1QMtR5wvlKo51d5HeIhrhDzQh9tl0y
39WcGpaxj/2Pomrgyq417DmF99OonHkXuvBPtgJLdxh1LCg8WO+gwC1JhCN89byQrcIgWEMRbKJo
WBHngaVvDrB18TN6NAz+vbXhsyS+qydZJW0SGpEDmY5zceqEzeV8I8x+W/jB0/JY1+ZC/pLOU/SL
rbkh6X14Zbq5ZYsBN13s21HWglzbIPhLc6ZXIp7FmgUMLlG5g4uuC2dVpBe7MFZR3+jgMeyxEpZr
MLCm5+0bnNG2w9DQw/8XB25vwihtehOPud4drPAsrkPijR2XQnNveDnU7pADg6SuCmJKGDR1Ks4A
OkUxFRWrPYCsWU1dSWIn1LB4arzXR4SrTJjtLK+pYNx4/bmWXrB0b3o3QAceVWbZYHSUM2oTk79r
xg77F2h50ClQ6Et12w82Fl0SF0R4q8h2dOO0JKTfvntvYgy1zVpH7gZc9zTGKX9rXPJNPtzSuck8
aamSgOxEeXuNQszGNepG01cJp0wSjdjzJeoVt2jRfX1hIhxHlrvnwuodiPyT5OZQNmDRNcDQVE3S
nwD/3XAPeMK2DJTar5p5Tc5CiXelofwMQnSrIzcF5VOwwwPp8qN4ZDIYYgiGrFLTKlI6IfUM+LXe
s8e77lwXSjrRlOvd+AQlrltLOrfeXoDDSfINjtw6Kv/QIe4bMYcfGI96AsFjavDPE8R9neyIVd3K
ERYBZd0lJrQCuMCc6QYex+N/tFEF5UQbruY5w8vvUuz/5iPId4FaitIBJmMV66qvuZeNyA9oRpM3
a/sEwdD409cmw4ZHsRQw7m4yvVY5kPSPjo2tvlyJwTVp36vPIInq2MHSct4+I0k4xH6IdKzKUyZq
WniHyELKS3VAtUnhj3XKKtSUU0Y+iTRgax9rdhYgZ12Ri+/dLIEXjqI8v5L6yMMv4QJ/2LG7+sh+
C/DvYlkvQ6VJzMGd8507AtgGI4xjhCXYlpkFLK3do991CeC2Peo/VnqO0C72Lo2jAVysv1T7JrS2
1pvUxDgnB9HqNnxMWuhDZjSA5Ch3l6yz+d3OynTZNknjJ8sRt7/e3wM+HDqC7MpIpzOMAKuIWFpK
3N1mf0x5cq0AjPdGxxwLnSwbBziIX8o5ctSO2s6uweOi6qmhyGh0J5qI1nyzLvokm0Sx3K6eAFsK
bYWLyzhs4pq692J5wah+/yxIJhVmsI4UehfWzCksVHwiWlCwgSa78k4Gf/9DoPlwKLS9NlLg4q0q
lWt+dgJispeugOvQ/XFm7v2qIYvjVyoPchUWDz/l2ZUfK6vcaXykIOIG7dvDTA0rp7Vd/x7zaLXX
AJz0C0afmfLT9d63Ked0IcdfWcq7wIWqa9gxYm/+lLDLVfsMmp+7JEgyH1O8y6ewFzUrWdJogR0I
1aSxaks14uPp+aZkBYilHO7RCKm18p/fRyVzD2qQJ/LfY+Nn7YfGL2wBTxIvHhEw974v7JHMyH7Y
bxSogM5oLX6wC+us3SrScnLzDI6kZ5Uwcm08O6RG7+DC3VW8238LBR8lMQjY+eHIpgZIqXD764yp
cMElcGclxt321y9xquMnWXKcpleO8LGL9PpDurVs9PdcfX4imiKC74gbpTNt+baDqtyHM27svLOg
uUwVmFO8DqqsszvF51E+xfoJKbaiKWmtfPG0R63SDWQWFbeDsOnDMsxHeAbYtGSJZT93V/o6iIuY
+/QnuNxsi3H5A1o8sKQZNNuvozjZDYPcMcyEBHtLoy1F8A5TWAzqJ3X/Xv4j4inM8n97XS5cyYtQ
bkYx8SArCB7xMjFGflqeZs5s1qLifh8CdzrRoD4FbWprPGMyIE7VK88qLCMjtlCGInXUQCDyMBWC
JgMSR8hJ7twJxPBdp3B/EBSixP2LWfq8CHtZxDSJHcEC0FtaNFXp0Ix4iJP/OBHTJJLAWhQCsV0s
LfYVMJtYaUwgnT6IfvsDUI1+565ezvRolRoyXCMZ25M23BKQ64xdR2JqwBp1z8x7gc0pthGctmhJ
7AYwHenPOOSs+2L+0s1MBlrufgniIcFWMSMuANvAb3pFNH1tBZ5JD748VjC8c8lKEKPh/YhRntzL
QAe18bhfSeOAh7i9gLdQsV/RlBHwpxnStG91VFqV7h5IuOuOERvzw2en9R86mcBXWDHebgrBaGkh
/4mrESd6oYIVWl78cI1SkvA0bE65NZKlu4Ee5f/YFQN/ikNaVofnjx23miXuxcLZ5+F/ADtxs1xu
ZUDvsNjNdy/mIrlYIh4WdCTa3gzh3lS3dxu7KEVdafJybGYijH1pdAYgxuhMt387wFBlkN7Y0jtc
2bCsUbg4sjdUqgBO5OKK03W6xVe3cma9/QP5bEGWN/2Odn+ai6ynFy3YczeHatMPexFs6t6H8qy9
HkAZI6Y5ZLEP4+yfCuOPdwr5cGP2Nu2QRc8uqIEPEBa55WR2jns3VhaEuVGtI12tHvxKKwno2VD4
NtCbFxLD6hx4O1P+cJJjvaXCa3/T7J/P6mg+j7dDiuOj46K9Y8Z3JuEFH5eWw1B7T5C39BEMZdvw
Vz4UCKhwtguCoYQ0VmfCS6HBSEXQz3lajC/pnKm+LH77Y09Oktj0CKsnlniN/WYnxxrr/7JYSe1+
NyJnsFyO8FdjoN8IOwxlmzrgYqWzESKKAjWtk2lLgM1XbJyobmrP+OyRNKxCEXe7lNS7CzYe4tLp
BRCBjQxdLi2v0B6yD43/QYj3juuX+w16k8IEMsfYFoWR3cJgCLouUwIWMfk6jGUBiP8Zh8njFHHZ
AoIb8jl8K5pKCs+Ud5U7a+82rwnSOTOHHsMfk+cnbJXmVLUXrx87FKU3N83aUFWK7hHQkNztlOx0
BCkhKJa6k5hSm6aJarckNZUE5KzPfOrfpzR5ReJ3K3U9pxgOvnE1f+x0a9d7n/M8BZKwu6ywny6C
v8DpeumYwIZxf+ZU62CFuDBsyLRu8RJiNf9bAMoQQPV0yD15D89fCdxSEx/AB1H3ZSutAyd6fcwi
iRotMkZHAhgBxjb6t8yAqDOE/ZqtPm+YKRfGSEWdj2UEFrig5jfelZaW1wAt7MZHfzpJ0DNvURvL
MCXvcnVCXXrUrEfRgjlnb9INgk5M7t75roWZyTjS+uptS2ihXs6JnmS+Pqf9/sefR/c6NRolMWx3
/SvC/HO7rxh8QV7PxlDcgLT4Jxzj6osIPBrem23XMFgjJhZDQR8ebqKei097pM57aG7c6Oy7Igek
hHo8V/lILRUcCosz40weU9HIk7xSw03No82nhNBpaH7d7wHvrPYmJ3iquXo39Dq7OoJJSkFYT7Gg
YDipyRZcGlAyLMuZfS0ZqyhIIocws2nl8QdDCqdGzpXX/0aiCNUN83oT0Th1PmI+Dqqv4c1iTPoh
J8WmSfVhjhbLYOyDCZFdlaEFB3w4uT9dWYjsHxGHmtNec3dFmJrzuDabMQ+GgUqdboNm/BLfsLtO
ojDNP2ITd5hFVqwIhfXMjMhW/47+ROZXll3TLaOC3NlMKv+FxV3aV4/QMOKTErQeBxMtDr5qvd/q
1PbF0W1TW8N9hULoZeiZceIsJmvprp37GSOmxumIZLomotmGDHZE6g8paEI3lQ6UV2tbgjtUV1SW
g+YV+VjDVIdZj9Z2pZ6jDGl/tJz7EQzoqtdoB1lTkwl7hGatjEFwiu5mdwjIXfeELbIqxZrmllfq
GeKl2R9DIvcqNIeXMyfWnlddg1tPFKGjmx/cnkh7kzBbLw2qlcs5MDgrFGfN6cFkrVahZJMtlD+C
wvQeegNrjojgIeULCuWGYsJDQRiGNpfhE75L35JWf3i91dJn03QAB8mxWfdK5TNtDzsS/JI07M9K
IW4dknAFv3Y6LuQWe5WjtY2sbeKeKELVFrlLK6e79fi5oEN4R/aQrhBkCFuw+6misMbIVAxQTWzR
TyDXwekBwmAXLTuc7glK/xsG6UGKeWK8aVhuthvc4boe7yppRXE3UcXh7xxBcgGqbWOTf5mJ+iRP
MDTaBR4/k1WPXi3XpYHQIhtUukq2dGnU4G54avQm7ryca9lCoT9umZRXXXU4o0a4RsHqeDboPV1o
Sa55ST6BjnlepC8nMCnwdTfa8AgAQ0qVvVcecHSXg110IoV7hS5XPPRC+nItNcePe3c3nQTzEdn6
z8iEFLf4rm1Z1wp8DO2Z6aigV6QYis2yOacaR71xLdKaC+/mYHLZUm/CT+928kliEW7A4zdqJMin
vubum6AsMhWaJhj/OmtEF0vv68uwWkYQYjnVDFift6klNAXC/SO1iCEeKJE1Zl8Gh6vAJKAEDWso
nwqvUf/vyj/FbIDxVnWNCXYoblDy1pgSw5tLYbi/p1jY9Xb+c7Gey5nnL/oaEramsvyv3XwntQYN
06npFvPrqkY/dZiEvNEr4zanDBqIXoSRjpuNvrb1DsCLP2Tgv0pOEQClqJ7RPT709oiTXh0juTOv
/CgxMevnciuCwhd39qqCFPh28ili4qTZS+s8yZ+xso7VUQWWjGQLscIW/jJ8H9PNbPgNi2BLRtKo
mqrcSLZTB3dUv+tFljb9I+ioHlp/PlxpbCLl8Z1jAjfRZ+SZvBcslALvIGBn0D4MhhshIInFv6c7
g+2Bf9t9SvOUhpvZshnWUsa/W52ApPGAePOltUk8truvQa4qXz+RXY4WKeYlntLyvodXVDkI62Qb
8fMfcwBgC0dB8dYpjDyR57DnpxYhs0dL6kqpC3NvGe6nQtA+Ib1eNnY9MeFFIeojitUgLyVf8QIy
CdAQm/J0O2gw6oDPbvELQXVhp6S5F75Z2xvvWIDf/lK46e6nalejLLUVo0Yj26HBOJ588PKc5KBw
CwWCrksUJkL8cp0tY/4PSIJGqr4/3c+LGd5jzJMuhSi8tGYnhKWtKde3HvxPUFiHEVwR4uvFZRfk
rQT94HA8YvYBSV4puTlbueELVymkB0hTaW4yD/fYpANmDalBJNZfFTq55VNmkomTUkwaVL6rJB9q
tFJDEF95En3lLScoO2QPH5LLYon7zoGS7R2xuDL+Q5fuC3N9P+XrT+cnDVfMqHF5582VyRJDNGCq
AB0TeoDD/dZuve7eEdSidEf4u/xSzgEGeA7oZP3REejzygmt0lGtM208DC1YPeGBJ8lf2PeABRLn
KTcWMIIPzB0p+SrYCm6zAKfZ36deJ5gH8LzsRvM41IydDoIEK0nx++dJnmBTcODelNRi+Fi/Hhg2
VX9uNbeXxn4VwzXPmPhWGo9jNYEPK2zx+cc1jtdYWAHW+utBlK8D0IPbHlxtLy+u/6p9+i+tc1Ei
NcPAgAaKKYaQJZgUZX/6xwDuxuEPttNYBlengroG1lMK/gZQ9Fz6fcjwR3LBC1Cu2QZ4lOWYBF0T
fcg12SqHqkeFqoGDrWQ/sh5lQaGP9LrS80ueoRkIHM5ZoG9b/+YAopANPPEXmWnvWMSupc75Syyx
ar5Q5Euf4OtrB36uvZu0GmPgVifutzNjzxRR7pwtotVnpm4KfyHIvXuwzWio9mmM4iSa5Jx3G6Gl
i1Ba6Y5VxM3WyrvtXKpJ1oubyaGp46K7buXEwQZJ7EUFwWleeFdW2SexE7Wwir/ikXtG4KZvUsHf
zQwQodyb6LiHpAZfVhjCOaVNMwf0yE7DM5B2dRviMStj/XUzSTqGnY9V222Ci+jj3710BTch9dgC
bJLI7RTJAOnnNT+6m6ft4duhMyz8Twfku43yJNNJHQQy3Ksjk4kW9rqMuNEkPgYbrpbIEYPAM0Xq
8EeTCSf8QstraITR2nigGFcx05NmAkJOQe0m/1JR6OfUzDw3LW3GxHhCT3hwNI311RFhFrtUDJhh
3fs1lItVS+yHZD17pqxeZZGu9lWUmad0Xd/O/n0qw6RVFRGt6onhWTUSHjSMmT3iWqPI8043Y3fZ
knVO3HluP7prFCEf0/ksczF9jSMuK28ApbsxbNvuUvkvD+P74r7+o9UY5QlL+4bjF1kLaNg7a4dX
xIfRnroL4Zlj+UH7LxTQT1J29azrlDIB/oYTZrl5p62MVLy5YEll6Wn07wD5GaIyFaossvV9Y50h
MacTlElasxXYYsDxBJm8oLeXRwg042P9c/p9plE7c9qyI9d4fXD88KPmCqGoWigNGjEdnyWmIHvz
CUYCaC5QcgIEgyIiBsp8UQgha1MTi1q2ITjXEm2CMiw759Lf/8EGYX4y78ZhPItD0TIOG+9I+zkf
CP0Ak9ldTbXCpR/jAJrzROJnVJTjAPum9XGBah/S/EsZyb6i3YD/GKgtXG0FkO13TTzZ9FCug1uZ
TVb1bIgU615un7li31OT5Ih4z1h48voMYk0eXNnxbH9dPPVNZr4QXUGljswq8MSBhvbXyrMjXsJH
qMXfUHnitAEL46UePPNWbQI/ztAumVrwEAF7dK21/er4PoPr9fFxVb9qYnjbVm3p26PqeQ5S59Jn
pOmUWqruexaojbbqy7XXYuqBLyoZJT/lBzsQ1wHTJEA6XSfsveNCrZbF2sckJ8SMedBW4xYhRTRr
x+yDOhyyKK9bsnhAp7u/qOhqapqQm5kap9yh/ETdocvkcU4U8/vDnvre8h/vSUgiweLtmEPVHRQ4
bDt4zTpFN65/kM3EFU1STuDkIn2xiVtEpnGD1FEBL3qfkaLfNpKUtoirf4kFeRf68rmwlKMwbu0S
pBisdBfC0UbIFM4w9CuAlEd+dnIT38STVS0pxb3Ct9Wl4ja+2EHNuCsY79hHFeD+I7/GHuNGOPg1
Z0kAvp89GuxESqk0T7Uwnk+HjreEkdNKtQr05sqCjpZ/ia0xgxJT6NBhgqn+Xs7/wm6kOK8l8lQ6
tWVYrPMvaUksWnHdZE6QDKlHLJ0B3r2RNhyVhIyNYy6Ai0H7lepWbc1vUIEu3z5xZxlW4AVk8K8p
gM2L8BwDpwdUzKFWAs11z2t9TDprfBMyKarBgmc0puYBoK+rn9CZPS+jL74kyOvD25PFwXx8g+iW
kRj9j7wwhGv0r2BJDwAGB3wem+VxfN/6A2LtEchMj+D04faJa/XC5voCFdzk5i+CklEttQkMzIZm
PX9iL/WEvfFJ2EOWqgOmKYIaLaJoAdO0S7295mFQgYuj4erxx0j3whvaPPZKqSD9XyYMrHoJNlyb
l/hmViU1kONN72vwe7ldhEqE3mkplFE+SgcDgFYwcmwDMqGNOUVtUtdlOe/JBfsuWaKSLz95Qp9C
nFaNaBUj6tF9SUEDx3Ulg+uPENpj0tuyeWoFO2FCLAvUmPblWOK9fz+ULkKr4rsbVcRWp8Tw7ZTj
4YcgIhMQIa10w62oHO4f4fpRcAu9LskM6rnLE+ZmQqs7ddr5CbyQCl9wWpdPEhCgcCSDGkzclVR+
MP/fOUPA0zGtt/qkYIMo38Hkt6KqQEra+6OPK4bd4WfYVCG4xcGEPQK99JKw8cgkT4Oj07tc7dfZ
wwfs8p1PNpxEieU7mInPJxXwuoGvZpLe/8umdhsatjcXCHoZIfSbA3n/o6ecrXl9VnnOZ9UM8OhG
3LiFlpAXJQ2f1QPkuWBOkCdu2avrSTFwQnOHJqHIO39eizRyuQ9WqHKB+IstokzjG7ho25Y/Fysn
4eduf8cOfOb+PQgb8zbkTSS42utbeC1zC/nunGAgt599ogli4SG0dgWEGSMy0zk3XEzRTsWcUZt6
0gUdd/LUd+upWsxuiFiKsw/tuQhKLIfJtPTD1t+9k944n0sCQ7p5xBbcGC15v5DWNWic64LE/f3G
mUCVqfZOdbLw6b3YZSgHY6Kt4PvVFgDTQVxwJN+N2hH2rN+xsp9cvYnsk3BjFOevPLJi987iiUbo
BGsg0QARnizdwKMEoPfWeY7W0BgmNMRzWwrrF2WUAHuz3bzgBGx6EIzoVz6EBA/iC7oAWyYnVGdy
YW6BMWGrVBU4Obmcgv+VnBTe7iA6IW58fnfctU6nIxNcYZaRTiwg6XMF8MsUqwZhzQzu+nav7eYZ
PqwiEC/QuC9U5UoZDcxVqDbSMuFEmHDQ6W4RQZ1tEP3M03H8MEUkjMcSOmL7+WCIU3j+6Xy5Mx+V
x7Qu/p4nGSP9kFTxj2bDPYdrc9zR/PadLhFwBs38EFWvRxdkTOp5Wr8wDRWvly/ABFvOyYHjA0hS
dMEzmu4UMwoUxQycmgcyACUAPQOKwZUKJy2fOdB/PA3Tl9cSG/D7dLBfQ1VqsGi+uX0+Mic/bVOI
nJ8+RxiuI8XZbePwbuOH4GOF3vyYAlIZcCZ9MThvhZyc3a0RDvUSD5sVgzGekelfvA2UCLWLMzuH
g0qLRS0AAj4hz1MNvf8Vhgl9lCAsJfEpth4VHfHlZjwEYXmZpifbqL1A/09sHCAYhZ2kj6pQMfHb
53O8ttMXSyIRS8y3KtmgQGLDx2wWi43Yerl6Vn0xH+D69R1ShY9ETh3WqrKOjfAhc7Zyx8c3UnF9
wSxANEyvIFNa4CDN1ELdVGb8KQ7A+UOulsolCdlMEUYjfd6Cuuv+5KRQztI7H6vDTZyvUwu/4I2t
PZ2Hs4c+iYDJwxhKCupmZKqmxVZ4aNkCtX/k9WF3+Ot7nLyPeNsS+ZhnbnZc0lrBcOu+FeOI+kZV
knExyVn+k2x4M5bGDh/T4KiI+k2NCdd5yUkP+9Rx+89kd/K7R4bELEd4S+9dYnX5J0G0JFuY78lZ
jwen9iA9LOJEjiXD+vk7HjTbvqYfyH0WANfVB6K1XMvJkO0cKHNsT4xBpaxEYHHi+iyF2/qJWfu0
SZCvtsuGm8XkGUdiXVLVcgfpQYdrqM1sFXbat5+SWFMAzdRbYZZtcOEhKjW/KOZ04UGFEpA6Z+PS
xhiuXhZsIxYM66sIwah1Ni8yj3Qwei+VQRSLMliXsWMXQRhSrWRQI5xMHRSAiuT6Hax74PBaRTNa
60Mt9gl0dSarhBMIGb69C4xxAwX5vRu75zuJFxd56H3hEccLTpRsUk+tyTezuQvwrmyjFDNWdV8W
qjqG3g/ziWKvVmqp9E6bdMhaM444tl7zA1pWFVRZDOiMZAKxiRE3EDueZbFv3O5ptX0pGJ9sx4uy
uHWBM6jwCtKp2r0XCyuHvhYFZ/KgMcz6Ss0F5NNMMDM/u0E+YTJcsmb4dSOgCHrex48sxW5qIJmB
1rzPdfLVKwdrRjVuA+Yni1rHHzo8gWXL0fmDxxJw4bowERk9yvUK49vdXqOGNGgMOY/NmDRCbNCg
DXn/GvjX8fX+b7259AyPzFTeBjFoi9iBFu7JaEKr9azbFzUasTh5+L6p2xtAkhY+3k5/eIKu+Ujz
/Ng6D0yFIyGmOHZerKWGRdG3r7J3sssYjk4muHSDGiOw2DFjTSsfu4uGdKdejvepnMcaY1vFZwuM
qDFf/XsUILwDXd58dTTqDvy/XVYL15aQV8cvv7dGHaK9ip104wrtt7bcCEQdHgUXuKGqPMUtXGgJ
TZybLOHZRnVR/hXvmzbdITEKSqanTQfTLYuw9w+o3hBfI36W/QRTidUmq15a/hlz0cpEWeHRaUFc
Cq5IustOt+qoeRytaP5UmMe8Z77TLl0sHMgqGYBafqErPdkKb8omtwv1zbdOcmJritwbVMJtv653
jSBC/H8sNGjDGQINMo/cGA/dMagXjfYhnTxCg2kr4bC0qKkn7Ts7ov0N+oFV8Bs5jSdsiWiPVCip
BjH0SYCAc3i2WfVft3x2kLIiC46UqS6tipxhjUo4ILD74JO6a+JL5nxY9z+IdCGi/5/CC4AEUAKE
S8GZlXpChmq9uLR1tR0xUlLeMlPV/tgS9wd6oNjq1NzRRJRv8z9h9g3gt7P6YMrEWyG3MZWOmg9p
b70wN07nUICdFYiqDLWijzwZjXInBDEBFLsoMD4Yko6oMmVm+dVO8NyEjUOUuhOyCE8g046BcFw6
o0O3Jv7QuNLQmVbLodsD9nInpaxgtaiwGGs2B20BOgXDklvVwGD8AErctAwR1KrZ/5FT28OCe2fN
9/4p+uEfBoBVmlt+3f9HtftqoeCvxOx8AynuejzjwHBHYJplK2QRZRnpP2S4xs8+PindR4p+sB8G
FvT4wxw0W2VlBcAOoh26+572EozCukIije+OheW3+qrDfd3JGu9seADGb5ksI3+Vc0fG5340EAvJ
B/nlvPKa3JT/YE8BYtIzufokLYrML5OYNsh9eCHmpQSp/R9vKsVwprJ5EJhnuscTImGUqVAKc1qn
gKptBBw3Jh8je4NiY53uY6lDTc2Y+NRLDJeguWIjOXdrh/gD73uLj1drRum9yImMrqExOC82UaEz
rMbVYyNRyAM3P6v127rPFFabJnNPHenuID7fsQu79tsSb5Lcc691gJOCLSZFN8z/tWYbBEMvIqXL
JZCXxcYiw9yjHC6R5BJFcwit0yupjkA5Uqqgppijz0MAeIInELVdYZt/n45KOSD5mujjmZIU2MJI
UMzMIsL7FGoZEv++QeM1fsRCXjWwQvwmew3UcXhVdBUpkNJW0RwaVwAN+Yaia2JwIAHlruWR6U7t
1N54oGGxwJivVhQxHd0apvahn2SLNlpTSmNwb7211JhBFrJeCfhfGIQaAMO2liI8vwvkE+n2soiB
u3HJ2lDNifwE4m09faGjo+L+zX8Kq0Rzcai5a6t+aEoFhrH6Bznl9ODpkbyPEF1/v3nclt5q+iWZ
racCpl/wFiCQj91OSfBQ0rS5wpgxkgG31ZdsJ3Xieja410tLjB/sUVhHlo/o2ZHrhtAmAHm2b8MS
wNs7Ic3j74bhGd5dnW/64whQYNzTq42ApS3jY80vnaBxMLPKhFQ/ng4mhFzO/+kbSc2Y0aJouLLC
Bkz6DqE9XF1qlK/48JpgMm5Mnd4OQDfqPrcj4VcHOrnwnt08Ksl+hMn6VTFbmsg5wOKmgMyQDzmp
Ukqw9W9j7NodKApurpz6+TkLlplqumJJOJxlDPudhhiM/lC/pjx8gK2Yjo8aWW9FOYY0SEisbuSJ
sfTrj6nFQPshoqs62JIi7vCPLWfNgi7DxIsAR8rVZ5pgsQ3Ev4zvfSau1lqbqkjlUz2e7zh4IjkA
uvuDhbVrG/ncaH9Pyp4L2NseerdC7l4qE3ZREtiKD/bpESOC6vi722YATuzslawPcGgcLCtLU5az
ZKOVoLfzeNcdmjzrDkoQIb26PuyUCwCb/e0hgoYM9UVq+wZ4e81BzfJG82Tkh9qdunOL/qKatwNr
e1TX3JG5lhP/cfS5ZWVr0YlciMn8L2v4GEHwzV2+dQEteBMvijg2RevMESShYb+wdb6b06T1GNrl
3e+REH5cFXRxM2YbFi2WN5KFZBHm2dgKtsP8XIg9wtfwCjIcA0ZTDuhVQ88Q99LkWJeMYSX4oAUI
UE/urAavix41t26JAEJHnDcJvY1GMz5Oq3nVZSxlA4JYmMR6S6Dd80Bfy4r/KI7KCspk1qMJe59i
zqkmA1brHIYNlLUD1C9Ii3t5n79uAaHbHockDZF1JyaCZXCIf+GMkfCuKiG2SK1DHdqU7HjVigdA
dGuefNmIPpy2VKwNAG9uZTIKdfjsCOWHe5EnS+FUZv3QNqz0v7V2fsbPAWPyL+GltmHpazFpaebN
2Vd0RIOtxXzL7HPOFlPk5l7bokL4RaAAPQ73YKbDF/XAt5VhXSiJpthX7EOf2BJYWrTk6P4VE92t
p/vKasJb7gnkWiV40TjndUZ7mQlu+WzHg8QxvO9gBzpVzsPj0Qi2UKQFW+7W/GRFtghrpRu/naug
bQ72LKiirEGmR04UsJIMnIutZi2kXR1ytaCBLOaF+o6dv3Tga15avE0PgFDOSV14usPG1HBdeESh
AIZucUva7aV3WbXRoAfk6jpVY0dDPc2icO/Y5oyjFXCq9OwAjVTICugXOF6k16w+kgDh4ksQsunO
PeLNKItNnSZZljaTVJhYHYGzdr9XVMt1sVv3UJ7WbyA8f0cFSDwmHPsr3ALuhsOvTlb1Ru7y+X01
q4/A7a/P8TUjj8XefA2heZCkBZMVfSdqMTSoBRFU/aLHRKr+hRDC1P4LTLHZfuyN9xZhbbnAzQ+I
IX7Tk8tXkLwfBU+S0V0+E57GTGGqhzpnUqLrW9b6R+ogd1Cbq+VBoNH8F/7NtXCS8eppIHTcLYvt
FeFNlXLoOxjpYueHk5HSoQyuNkOKTN4WGHZA3WlmzRlGFr55zITOyjn9dmpS5c6kHBuTwlmfrUGh
NFZSXj2/MW/W1nqkzctYs9m93qkWn/bFj6kBumSuxDptNQf70qsbLpefw0fGtwk2A3HB3GYsMbK3
M4MaJ53Cemd8UJklAD7GaTrgJVJGjf8cS+NZQToD/PMszLxWtnAPArYEz9/f4doKFoL9zMKCbf5e
T+CECsZwBXSH4+jkGuGHShO/EtXE7zHqblxAAZ70TExdfK8y46KlM9GnJQFB9aTr9b3Yw8vdNIAn
G6mv18LhxxRV1LIVenoo/vVYYJK0ItICYCPvu7bL7OrmBz4QMt23NQ6gxip5VMxpJxoxz/saT1db
jTZoTBqLrWow5Tu6fsT3Yq9RcKxiWhOR/QllJEgTj0LiowUo6pv/b1hGcO1WH6QfQsy7R8UIdqu1
FoeAd5hJqUan8ngA0P3/IQFETO6t2L4FwvMTYmxgo7+FFGivH0C54YC/MRIq9UNwW5RTAnz/w6oI
kMCPWipjYeFhArM+tf6cNVEv84EJiQYp+k2eVe3MmVIf23nSffnsHd9QZHzJ7rH1nhuof/4bs0sb
EciVbO/kyC5ZyCK5r9mRtYM+r2B0wNbnd375Cq1BT6+t3hEF3Q7g4iBEjHiT+6JaukN3J8GW21j3
qBaWmm/IXHtv+D+uSUOIvKiSflB8hXsaBN1sJEoheQPs6v1lJG0VtldJrq11Opc+z7neYPijQ1+i
HxzJemhrp4Ehu+RKvRwcnj3uUYRuCG/urbuCo0cb2ENEjrlBLXheGKV8l43VRkTt2o8klEAbviys
llOxnBon8/JljZtVSktkPrsmAjy6t9Lq9hqVxM/AlsP10UQNf3pNKv2QOXaNVecU5oHXFibyvOuj
/yLR29GmBfLkJzfcrvndPr0BtyHBhAyUk3MgV/Apjhb3AMY3hFXcjMuT2zKrIDyNijsGD9N0/ikg
Hi3YMpbUL5tK2R8QOVPV/3MWRzNAttDLNse2IMrGLAIXG/GSZERxaDvxhNj+IYih4cE2BzNpufIC
TdaGSAbzJRCMOBFFkZ2VQe44dMyE5vFwt+yw/y1rOHn9Vgu4SU9eViXSp8SrXvswCPS7JU/dU6o+
XB1/gxh3lFE1GMIcOhrqQoGoiZli97ekLb4klEsTaBI+G/kmdysA4gbwXXbf6jW8TBL63DZZnlI6
UXnLrcvmlJ/rls91wmKt3DN7quqlgOm9Y0pIlXe9ShBKxXW7QiYrwa+cuvU9dYMrRCjaKeNh0va1
vd/pT/83dcJMDIDFwFTlOvrFQL5unb40cmY/MrYbGf0wXfXCyU9kolQpQ2XxcYU7IXO30pOK43EZ
fsw3hEBYfdU493sdPSxv5tX96ttVpl7QAisdUT45oN7Yxm5gSUJ3HHA+W/qxCHSHRdtFpU2GRh1u
GACSKLk0stIgSdmCMleb2qNEhjVwR4nJkzcSeP++hfjkoyhVVDHMA91YbiJanBc2ZPEphqDw4e6C
wGJ2Ln6OBdhKUXqAR9DZeYdmDYMU6NnRSXHINRRh6XtHMyvDAEIrSP7Cjc+7Qjs3hxR88YeTtM3t
v71TmcfZg3O2WqXiCngRbjSh//XMbeZndaTUONxjPNF+4/COcfa1MzoW5/dawuCVQ4L8PUkmYdNZ
FyXQkD0bXNz47g0rtQlC2/9sR3ttu1WWyXPipqxTeyXb81are+BkD/gqIlKb9BcoebEexIM3uhj5
yBKujHDhrEuTxJwKWjQZZgCnu1Xpr/eK4DrVdcor5x5+o+H1mXCiBwZBXhGmJBDwNb9/CFPRZpXm
fZ37UHEnf44cMqgqW1QriCjnwC4WW/5b/khtrF2K3f0rbKOhibSaaicJ/glrVsUH0fjUEo+nOe8Q
qYdvIQdbm/DKFd/oet+YfEPx1Jvj1rAnVUBXu9WdIEBAYXHda2sV2UJ90JEfyLYEHNAyhDw+C9/h
jstc9B77BmLz1D9+nVRNgP/GveQkFi+Ir94C7eJ4Ul84wYWjqCJFhvmPOrWUClNhba45ZMWVmqDA
81Q22GLh2LFl7QSIotYZIdbYO5ymwNhEAQ5HILcg2EfURpJUdPjaThKL4a3c0R0wTSl1QSRShI6/
eeTlxdnE+Gpq+gSWkGHRA53r13reJuiKP7QW9BkMsYqmQtJUlAD+lufjh81t91Q3+BXIWtGc2bIJ
WIoef1yq8lUEl9gf02MH2pmr882vKnaU8d3jdxQcfxrmc+PNSHXhuH+5wN9UozB/4AR8Gh3zVPV6
pkzePPPmg3hhho6GywjVlkonSginej0edT5zk6SiLXXoPuXoFXg9EafE5xI1OzB/pKIrlRUKiuCX
juXv5EFE211V4YA1qHJflI4em1mKuaVUFkM31fq4tNwsATtOh/nHSdBT1db9koya1xCrGCTeWVmz
v24i3Ma6Q8ZWvQWLGP7rDjoKKY1l5PPUyl6N1XDAdgLA0WgbLA9Nh1VGgnriRr56PlX4JfBebX8L
ZWYkEBqazJXI1bbSW8V4ZM1sdGBdxrMGnRluD2b10UmecyKuGzacKh69/zLA7CtKfsE0grXkq0bH
ZgKnL7ZhK37/OD9KtxSCY6uxbX+ix9l+csbayh6rqojdAtr7pHeZKQByEGQ9qMwzfPCmcdwCcgSt
MPasxf7r4QhnKo2Hzouu9mmc6g8a8eNmRaUZjrJ4o1eHlAq21/AAHSv04RTiCaZgiLtDGUnP9Q2a
/eJ5mvHeUQW9EjsruxfsVlNEC3f9hguSoLFbjbyPCBqi26SHg5UZmF6nKIIXQieIcG4QepbOARPD
1VNB1eJsw24VBYLq+CpqffNGv2GiDo7RcNGe0h498eoWd3K9JU8RSMRw/80tEHI2m5bJ9ZyE/2YY
/ZjQ7DcXzPTKs86i7mY2TIw5KM6PkdnOCNxDl1sPDh1FzxiZKRGjQ5JlwKnW7hWGYEHHi9rx1Mt0
Pr+5XogBEmNrYGNz6u2uDREaSoHRg24Z0nc59hvk7PXeSQ5HJQ4HHx3RmWipVUG6L/f/PgXIkdWd
0beDPAGvzLGZFP+ofA6zqsqAk9vmXLaFzFdt92etVkWUkfe0nXkmxMoC77byYJA08WDmZPeew16J
1+7se5CHp7N8CHlz720HaxpV8OfKz9Zj44+Qa439EBIxTCgM8PY/K6Hs46/tdLHUc8BXG0XtWxAA
DolfG17BhdPrATqCkDD9KimCQ4YzLD8cGgdy3Z7MpsnfaAgS2Rf/dxpWqdHGLQkmMBVfXtXFa4c5
J+HiUY8K/+Vi9w8fct/QnlDZJT+J+vRJb7BZxBkL9ncR3FU3S2CEkvk34Ovl2y0WN368ZYrUF6Tk
/MXEiPz1zCBNT/PtM0FsLDxfAXVrI9xhludSUoMTvk2LDLe7BYP7syBZC/75FE5zb8cxfRIvokA1
GYLiueRdrzfQAjBn1VKZvangAJcKsa1CP/d9Optxy7/mr+9WOEGiCXoKgPN7KqhN43YNkaV/aEwG
3+yQ1aW760BeKYczsKhB+S4HgSFqsTX6CsZ+sz3jAopoXbEbBKn868+6M9r8CNj768EdS6u13HMe
GAQ778DKFWcUduEDwWIr00aGMp1Zrv8Bg4pQwMC+Y9D0ZZ2MW6M6Pn0l3IPFHdkQuVgVxPEnRmpJ
MQWeZwpsEMaSA0irc3liZxoG/9vZnjouYj0+jItwyLF5CmC61eSKG94V5NSKwBXLfa7YDrTs1ZB9
1xoSPUU03Qrq6PEmjytnijpk1SueXRwSdEbKe34Otu6LwxPQjn+Kre4RunOcfgxwVz1QaW10dIii
ZMINfZ3hhjlJ7B6T8K+uquZKrlO1Rg3gGWdUglWTS2QrOje8dP8IMXNZryEhpA0cP3opsTMGF0Xg
9foYUy1F+wTGih5GhotYYSF2mJXseRyYC6umc+g5u4BQ+WP5r+e1UHmyZ37Y777Kyf0DQUlbMZLb
7vTY9oMHLUOP7xogDxJ0aMJd5Kr1mehGRSoETdOu5fFHrkIj7VpBYRSvlLM3cms0IhkjU3FfejDq
ArCyPkD/YdG8Nkatk6MEwhwsFUa84iLdAK5HEjDueA03gXAOTCxLlYNMCBsw7vIGUIjW+v4tvAH+
+OTUO9oaqofctlHYEu2NVc4rWyy3zD+uzCWmzcHpMo58BsHXXo3c4MD1XaxjiHbDCiu8yqSWZJ4k
uH30ClbVs11fXi1/33s6fJoCrQb61p9h/HT1K2ecAlMR90dNcWSrJupFanYxg9La7JNdE849Va/r
x6rx3Db8wRiaf3326kH3Y12AkbruxkU66TKqtfTW3bgq8DNOzB20zCvcCaFp3SmGUIRZLlHmypO0
RkxZ0n/qKZM0X2e5/IewtZdHauot0QlmGAs4Y7xL6Hvxbd+GyDmZgCQDyZ6OW2eCxcl4bE+U9bKj
vS+nG8/TomWXfEMdK+V/v8rZ6jO14NgtM3mTpI6PEXg3VYrvXz8+e4XU0otQi23PZJvK+purCk3K
z9tlqKvar+Qi2k28SBnuTkPafnJl1KwwkZR+f2RfT+sKV6z7mus8dZmNQelD3y7m/ivh5PWeRbyb
tw0Ch+Ux/bJIBIFUg7KHKyAUd8cjMVpt2USaeUpaa1lTGTih//Wehln8BczpjMrrXbNdBuAodxHd
kECS8ALYzE/T11NXd8e7kpVkzl7vySUqInBr4O4k4sSSOiIq8fdvnrfAiareCMB5xfmGDeDDNup+
GjSDeJp4l7QiNtSPbvR85dgRVmKLmwAj5PuPvVlb0E58jTzeGaNU/u8zwxelzLoeNJTalGoBtEv6
6lARenlgEU1DKF5qalGZn6mdkDWDIV2pqRQK1dEm2T/cvqMbK/lgE/0S2nUqwr95cOTke8GDEO3L
stePBc5YlR7j2qmK3/KcdiVtYVL2JYu9wUs/dpTvXbI77HdMpTc7Ums8/ySLP6c5qLa/eFAZ9gT3
ipmwKALVQwBSpAk/U/kOKV+19lRNS0qj3e8CYcmArxg+2acXP6vlbsxSavN2QNixofzpIHR0VRkv
pD+6aUPIhPO9WpxUbl3V7ugK+SpTlrz+HBgJomr4GbI5JJq4JBxzYuF+ioRdFOxiHVvj7QZjAYlz
4yk1Kiwx7B8WtT4AS/7MXoYW++uA1Og7VOiUgn/7gxfW1JihEqfdX0vKAkAuMrzXHvdrtJbE/C73
/Zs7qm6sIR+I+6RHmhCxmse5XgqIS2hrEBTBWbMc3GpfAdwBW+Sk/QyS3FS5DkDwOAngevzTIM0/
cwx7sw3F+ydyvT1kMgwLKG9tyy/QWu89Zwrq1xxK4C54wbkvWTVQimXTKyZnkQdNVYteHX9Kl8SZ
xPbQH8obN7vE9kRrbbh1wDe30CUBqgdvCofikwfwV+abcRINZCnTdkoDKJvUn29uIgPPq45QisU7
9bC4GJ2UaGIHXbmQ233rNBpHr0XOuh4mIqRdlM0UAMSL+iBU/y5DTBP/VqRRm3glQtsR+JMIBVue
4TO00tQ3N5ZOVD0uHm2gbLSzy8OZBRhqnEoNXWnoh6+PBuCl9cEqEyokA6ln1mUbP58wfKZtoFZp
L7Jrrk7+eySzBKkeWvp7Kr6dbJFNFBJC+UEqlYeb5OZxa/vRr4oNAYDyazHz8wHUMU3KSkH5e+mq
KbpsxJUAf0bt+9319V5eAKLJVEynpOB7DpR9/Fm8Y2KT8qtOASsXt2TsXJkf1HQrtRUehHEKvK1J
FJy6voLT6Te6qYiH0R1h71hGmMDXcVZoUad2GPPuZy8p9PUEdyuhZeeEUdh3UDpFN4Okk8tjGfK6
ZhjqSDol4d3gpK9izAzpovrjT8DkapURHzgn/nzjmCKaFsXUAxAXy/TdkL/u+WPTOnbDCl5Cu7ET
GjXrj6vJY/9k25uASiHfOaWeMT7PgFhrm545B6XzoDopwOlT6eDBhe6dFT0LTDRfVRBQKPmzrh2O
/1gpOPe/Ms8F9shd4sz9LWO8M3YRzs6uOPxUFVEwMga5+7FI7Ab4h0WzsvYf0RSOIPanLdQmXYo1
QEOccy2tv62+vusQh0ClfkrHLIWRWcypVHhnt28MU1S4VxXpD6298nFHriKpWKiWQzUbbDhKEoVw
Chr4vRP0aoVogR1qx/LwmJ484xYTer4ipbx925wlpznVekURaWCREIRcfr0L+F3NciHmonRkZKgh
pbYhYTp/hRrkywtb/aQQeUSywnrku3ppkbglZRFDwFdx/601ND6hSxrQMmfb499Y48+lGdD8Kwlq
PdGVpEgpjynzzJ1A1O+aslh1dvsxY1KP1z4xYeaxb0Rg0sLaFnGvpVxWT+BAvdTLHjbg0o2GbyWx
mP20Si/d6nznR9+bLUixrTN+8YuSENgYdwT2+hSKlt43vQyNz4/VtE1LOoMcqkC4tXRp6IZ4YgGU
2L1x6YP2LkLcb+fgJo9HjeS0LOLnoa/7kPNFtpgwWuuj5C8p4l4OQMT1BktuyVpRSPAff3KIj3Jz
sSwBoLp2La5vTbqNvipOU2r6X/TjNIzfh0k38X0WwRWR5KBhD5wG2NoeIJanu8k9n5rWzPm773Dm
2MfXkkdk9ueF495fXkXArf1V1yImBtoU5ZPEofSCemm3b0/Hek/1BVNxqmztUXK7N1LT4zZESPBI
gk9D2P3Nf9XzCn0zumuDdPPCOGA2QjbUrNkjIktvAxBruk3WmGi3s/b2FrCu74vUrx4q8H6JJW+T
KmeX1T9EKWAmHqSXiXqjrOBbBGQSTqEEvfOaHL7ld5+UUlO29hwtgPttNnbiTWPNYLDla9cyCHjQ
k9uZxajuhUI+xceIu5lICesmngCY7C2/9hlBezpjt6ss/gMHq0FdcFt9ib1WcpJ45vmp2SkJ4KIa
smGtzdWSI/jx8pTffiwjhlXHcxCGTQMolxeLvNGz+xdYAo2tRG8sQ451eeMnCNF8L3Fvi3Gv3uQw
yMt+3D1PZDw0Y3TMdx5Bwgx4RU8NAODAU76XI8QUyKQm+VmivmvMq3d3/1JwDsfP/xUCAyF931EA
Uz72lHhmaUlTSkD8/VRH04oPYzaejrGqoScEfCAYyqZQ/G/5kW5sh3HAotAoxCjB7MFx4dKQ5Enh
1HCRjCwUHSyCGUJ0qYaqvD8vUAICa5CSeLNAjo5k+pKbe4nRY3tdY/euojZwWVRhVBVQZpT8vnpF
1Lo2KOp9v+IWj2FrxkkFoYew0/GMUmjH9uG/98QJtJhAy7u2N4sLiuMC/ozolC1e/qmhV5yymC7w
J4CJeUZZVNe/fKey37mK3gelDMxAW8aYnS5q28Y9tzxaZS8pYJCzpPrdrghTttqVLQoMiGtFe/AJ
bv5oylWpJ5l4ygqOSjjvmnN/NGYv+azCFOj8NMw2JPAEEOpkvbE2syIj5P/+14EISpgzKmsff1s/
mOy1mBOeA8mARWcjSPSgY1rkR2ci3Srek/hQvfEGav3Cd/d0EU0v8mKcMmhWS8n7c+kEnyYxhEny
JiVpsZMovqF81pIir1VUvzSvle70febuIuRUZHPMdeLIo/LbhsLJVP54qJ3QNIvKO7yXO7tcbxWc
6jg3h8lPrwyIUc5Yng5/oYNoowC02JsSbA0pjlMejuUNaACMohelY8qnxhttr1ESKcIOjpj0lKsY
c30+2rtDBJKnRqVdm8wYGVR8n8qRRI2oGmst8daFt/+uT1z4Cd12N+fzW1bOrtXKhOzG7lU8bk7M
SVEZNlnbTtFXWeldOMnakEMGLgwL2nRDVKl99pIE/QouoOEdY4/5ICzOeO15BYj4Y5TdA/GJ3cmA
Bu74gDp6I2S2CGoYPuUDM/I7T95OrkfF414H5fpAKR8CjgelIbT8573G37jl/jnwS1v/GPtOthkF
Hu5xzNZBMR1Mls/s7FykrL+zhFnNhtqYazEQAjiSRMLZ5AQJcwoVQM31GuG+nTfLyooj1TWXB9PR
/QzLI8qqR2gNt1kmiBuHYnL4k5vJr7Zbiz2MCzEieG12uMP9PTlwJ8X1CfncCq8154Qjxyuexhfb
pjuFgth+uFlqKlTxtNVfEe0qX1ujAjW+B95iOdd677LMtWERgyvUVEuyN9WZo+2FDlJMlfW37kaD
mL5t7W6ubgpx/YahrCnzunKGoH1ul9OjDRckUZxs5RsgxMX6BeguUCR0SQcHACfo20hKDxyzZs5A
6OIfku5g5L/O/6DZamG6WyHzZMfONWtNtd0j+zYoxC5XXd+0MdnW5LFml44JrG4VwxGET728Usxk
IWpihS1WAe7GpopIC3pvto24xdR1OvZ0fnaCj0EXyIidrs4p0dDhvIdzpi75hXuB/WLU3X+S2EYu
eEhlU1nGNmeltquvhFdPhiQPCKXLmN1sC0ReSF49ShHiL/BVXxIv6eMtl/LMNjAWEvpS7Ur2vKwA
LlXIvu9VpcQKZkS8ZSjOglmKfr759cMrQ+VHpF6ISrnRpo2IenE83XxIGZY56q3rHKt+MxpoIg/E
S1kQuEWkQ3SlYFcCdQ0hQKnNfZ+3SB8ijcND868AX2Z0Rsoyc2D2PXXfBRAXbo+zL+foz/qDobbt
J9+NrPXOBf+hNlv95PAPeWr35KicYwEFTLOEZHSoLEMgrA4ice+9GLZm5OHruQ8icX+8749nak7U
EyeYvnZRYz/9Xpj7Ol8JdHcvs3js95Y0tOePu87tdY2wxfBLhus8PDYscYBkLYpE69JZZxwb5z1O
xfK2AXelf3lMOcSIMG8/5livz/7eUmbWmDIPfplAg1lQtmyK3Nt8UBuVvaa9G2DvjewPo7ZQ/qjo
1g3+En6eYN1PuFVErxZYIn0I5CyXIWZTFgjbFjWfupWADhZf3g+x4ys/F0gt5UFyl+rXSPnDxXjU
uLlloob2uyQKkFCbZsZL4+5dmOb2g3ChrkU/tBEKOhdy6vZ3b+PQ7RDNQLE8W7nN46ePQFlLJ+PT
yeMhUP5SjngxejQC4ua3gU3GkgoiiaM3ks0M0aXJWLb/zl58YZrVW9A6MiGdADXNWBGjUYqrGO9f
M9ATuU77sRiyFH2QSmqjpHF6vUPIsWJ+CTfwAWiDmdKHSQOToI4C2oRxUSECGuGVJRqLlHkh8jhU
/eE1ZeVvXBAgManLISJoUbOOTkiU2q34+rG3HQwza3oybvYmKRhsluyDFVY27xfjoOxvgc7MksT3
Ss4iK3dND11cwkHtKXZRW+WhcjVbPAH2MZk2GgGSBhbCmcOr8QagHeL62EwTGut3NwhD13jKLDMv
jDVpLkJwjj3mhiOqyoHKyZia87kPF6HAL1ICEIwhKRuSwqhV3eMnk/Q3sUxJfs9YHZbUQzBjrCLC
pt085X2yQFjTqUpuGPKH0t3nH2NgLSr25DCMEjAJorp2MT5bow6OGm9K+CQELpQPd2mfQrfdovsx
qO4TOf6mVwTIL2ik5l8vAqvNycvjiFQrvGnhNX59wjQM5rb1AVN3NJWlgkjVBRS2zJxsd/Ojxz+z
63EY5WWD72M/hKHgNZH2b8zfsPVl8XpPqHxzOzCruKdm45sQc2nVLvs637Ads1G+NnI7Tnht/oSr
UyQD5c7hRMOn5cNMMAZmyVuuN+98LMbe1ryfWsQ54aUoRvp+QejcIYwILIXKlhsNOYxQruWxd/eq
xtTwpArrLeYPxFyieTAdrtxwJmJT2eNg7sASKhUlzORUlIDQ8uYf63KDtJO4hFWLe/2kBXzthZXv
+c9Eg9Mkkp59plQbM5Y1/EjunLdZH3dksb2xVVj8qrnLh0wwBp2CgfO1woP32Oyj23eDI5TRjbom
8SNuA82gWFQQrjSWuw+vKlcsanvf8wET1EmYT+cmkTpXMqpvgM6C1EzSnS4VwfCIWOMcivWNmtQV
sPxJr2tCZeXukczJCoMcT/YbmQ1b7ynvEFq0mUTfpLS2oB0/PHSIgdDS613eXn8hEI538VyQgWR7
mxTmOyTvL1ygukz4UAotdA65Rm+Qr71aVYgFw6hkMR9FPCwOj5+VENLOalV5M61KCdnZGCeya+WA
kEklzK2Rj8QerJ7d10gvS23zmp95/tEwdwXmrd05Z/CXDbM4ENyrOkvsTiFEdkV+0tRH9+7+XEIL
HyeGsbUF1Ln1x4v1+y7j6vlQ/9RimhUwUvtZq4KLCHuU9V3Kikd7Q0WgEyFYb8XdiCG2jgWwj6Rh
+CqTompszLtUwzdVTWZj8anNFMUpPs8vVLVDYp8n1kkeWVZ1geqR2z1PgWSr0WeUmzLEIyd/Qj4/
og/8jKhwFmj/y7yy5BKA+yyBQPLN+RiadS8m73IUPnIOdNSqlStsgNpDLGjptKwJOuQCLG+kJH7E
LUbe0rqiz5GfAp9ep+uqW0J+1OP8nSOoIOoziM2KKF5jBrg8zQaS2Gpg7WaWu7Qs1FLLFzRQji+m
kp3hH6m1atniayYg6q84re9CPHEYiVriI/czS7HjmvJkIGU24rmKGXXY7LXlc5kZlTdese9fV6js
DSQijw5NdrFFPKcevinO4+WynVfcskC6/x5LleRnfmMrfL6ppWpp7mXCaPKtlk7wBIxHpFUDO3WK
JrRPdcHEOPA0T+CqFbz0ZBuxsGfU26iRJcITsC1eW7nWPkFp+guG6tNSO73SmtSWnmyFIttj5frD
zIBXOs1ClNr4f/P/LEIagjwdSltyoiLL+7APAkCYjndLdlpbIMwie6jCcTFRIMmMecnMA3tlwJz+
CVnJvZeIP/wYqTpbhMHhade5up6JDo6gnZoqh5N/ZQUjIZqbkY/6+18p8S6crhTvFYuZacnDYiWA
4sbDVxJi4AUgBnl4NcNwWxu2o3DeFY6YN2rRMawg7rB6YgasyrszdzjL0k/vYMaA94Ji+qSi+F1p
HRMDCoy23JBrtAQtTFtHBptyPmDlT8ORg4eQacdfMcEzrBBByeIEfVrStP3y++Vra6OrvZ+i8YNJ
rFcZDq4pNAAfE5vbUEhGtnUtwiSNcpbJPW60EEeh7OX5D9jQ2stRcU/Nmx7iF4ePwuW0D8xV8gd9
mful3mOaLv7A8G8J4//WR808rYamHcBICuRQpParm+i2xitb1e33tvHKxpo3x1aMwxO8kawf/u0r
ZteLicSB3r0fXifE1EEXY//2xIgJEMHFuPw5DMOqVgwz19I6XVGn6nxJk16bRPteKk6xDWPfE3Y/
nyWpiyY8lvHyqU2oP3o4/E0NH8G2Mh5qdpeyX0ETOEljRyxeDZvL6xNQs6CYh6ARDWSsYMXFg8OT
uyX74B0oIB4fSADyF59D8UZ+x0uKBD5Em5dRsxWEjHXXc0VaiGaOT++GJp3PgAmFlxK8dDsBopz4
XMCRmcB0OGdTegWzG6ueN/ZxC9hGxpBUUXw/TRk3RhLGQ9xj4eGeixP3c2dBfBvp29SZhGXtx8mM
ZbbpR/NvwCobLkBW3sEiwM4VFlrCT1Lujev7li0yUoEfu76ccUMoe1D18elBLM6gOkFNgDWpExje
jBYolejPkhC3qFLXgWb6mu8rwrHwJD9XE2lKeZStaLV47JF7dRC2zWK4GHoVNhHw3xPf+rzoZtGY
LaMXThsYytC52x5QQnoXtaUv3H5V57ERbQUMGZuQxVkzcQ3cWBB3Sh2ClOw2bjZPusfdgmv+WaEZ
rXK9PxaNBoGYTQ8uUKVPYUCNkTRPzLMqZCpjZzMOKZazGp6TiAWQ7Mdhao9jUrBhWpEjFTQoT5c9
po8HQHfemEhP3CpG+jvI62Vh5EfI/R4CUeIA8W9AgpM2HwlJCug7xI2pH6MZXP2FWVnEaAJDOIqd
B1vZr2tlNL+FAObji7YfkJxw+ewc6fWEjMQKVTwfNkpI6g+fmu/2TjUVau+vGRus/8tC2sFmxoaA
KxRcr0y061KDSDU4T20gNtk4dohncEIOJZ47atbaXd8J8WHNMGt5NrEnzlYCV1Po+Yb4SQtiBDnm
fJrAW/g4uyQ/sysZtuuFPgSDwLV7HC4hKWa7t6W2blNQ06+DYBluWG9llIp71e5Tm0UKblFnuTFF
R8dG+yWpVTXC+DKme2RVigt+6GIA2hnuQ687GgTvDTFOoRACWmzEUR0uiAP1uuuOvHhl1Ia/Bquj
SSkPBvfs3VKQv9kyJHG5rJq6uPN+0jS+DzHc0z6x1Ak0mNf3omjX70weAcaUqrXn77CDo1iva4yw
5fyAVi2ldGwZqndnJ8Rr7Je7sTZez4OM+1Hi4lOIv4dRoIIs5gC1mG8mCLNTPmt35Hw9oBBMqqJx
ycT5ykJoJrXkiYrzlNpQIuIp20iEYZArWvGPspv3BxR2Pjmf0SF6yBoyWhhwYRt2WWwLi6MfkCx5
OPg8woCgxdZtXSSTBPxlja9dYH7Q8GH0nvWDACI/8n2MQ5dhbbtLbvUaWO2wTwGe0LJH4CMvz1nN
Znk5yJKbdkv0Rb6k581C5Fn3CZxA2D0442kx/hSCcP++4IFV51qTmzA9G7acbgM7sbk+Z7nTjzR/
Cub43gzQmUAe8rlA8qqv6rMMWT8ZRPEaUbd+jkbdrHk7Rq5Pz/suCi9KRIk+xmyHr5b8k3OqCqRd
VXig8fnRnPe0SKa8azzVHOflcYd5NLFRxBbFaccjeKbt3iaevNn1OXjxTYmdBdl0KEdYCQKMpjfB
75lxwZ5tsDVbLkvQbZNgKoGK4OjMWyS9PR9hXPfrabm55JKK1F8HowzAAOv5DPk51dJ1wtdtffVi
ZKKatSKp6LAO9Uqv1TzmZdW26L+koLZHcJZWg7+1APesX7Qm7QesA5AGwsMzx3CIMhFAnPhN+fNO
WGkCLvLCfZNg9C4idOVZd9cL2VcdWsjMCF/IrAvRzW3dBEEr9LVJkxnzjtKoOfPGj9g0u6wXfB6r
GKxczMH1vGtfMe2MjjOi3vKuXS077luQAE2gKxrdl2G7j+akqCJ7+P0bbzQnZ1aKDr98sWblBe+C
GyJPduFbwpFhYyY3G8PZzVBstS67gv/cMEn6Bxmq+0JI5AxekeNQMic5moZLdUeQR0kGjGArU9uv
BdNIaOEJCvU03kwx0dgjHOJ1AJpxNqLf+7eW1TPCBcaa+GvCNUsSTDsaeIEKDqEVNTA8yh+/ihFZ
pZh5mXGu101cr3+zeQ4FBpAQzzurZtYe+uERUyX3CeVZ72cREhv/Qyp2TwXQ4rIJWCBoWRbnj+NO
QTKbpl9aSd22c0U2A3j+arkb/xI2k+txMt1SNUmamF+V/gnxPhrqJKdIau9IdiqftzLvkjEU3W9b
s/WvyL8Gx4uBTj5MJefyFjeD/Owu+ZAnegI/0k0PX5Nfbj5nkylTbQgB8+WCytFBHkMGiVbxq3QE
T3LxDQ2A2dg0ld+8652zByIdRQYNA+lfr5VPvyhPOmrYdX01zB/KHdWgY4DyQfLyykpkUkb+gtyc
2lRFWYZEXnTaX67CP+4Hdw9s+VJ07MSf5My/w6CmVA20jb7/UTlM3EaWH3+WOtNN8FFG75q18Jly
5upn2euoK/lbJu4gvtjgg1wi4ePQEr+72qPWbaNF4dUvdf1L33Knckxr/C8TbvApshAlXLbT6rtS
7E2RWfN4e6S7UrVrUdffJWwAik8l064vZ8dM6AohNtNIktmnrBG+6jpBi+s6eqroy0BZ78OIJiGw
EmgdzZtoQEWWKroDLKeiMCCfdrWdCWX9+4ReESeeD03ax9r3mnZ+Q7pcTcnOA65xJ997ZYHzQxII
4kHvWCOSAUGS6Bfvo3xUfmO+B7WoY7B9MI+26o6nz/gSoLBxdyuoNL4/K3AjJ9gdVCtaG+Di3/fu
dKmMupYXW1im7QipLk5MoKlhLpo45Abpay/2GmSyYuFBTC1KY1Hex577DW32pma8STA1U9p2W4Kc
kUC3mz5J5a7fTDrML2+Zls9JzUUBivQ+1HO6odhocAjzhCbNXl79xsw75NHNG/ArzP0MSqKemKRb
gjNJcuTzQWrQ0BR6Ura/ft/dTnXL0TcFAqPtwNj8Gc5Gy/JfkwagOpEcLLYB2qOm9hChOHTP6ChQ
ZXxMHSs77QI2aCIP2pRxNh4jdePw4dv6uEpthDBlXm8k9KuuUCjpe2OVfo0nrfa6KyMhSDB8E6z7
LUDzvG8PweWLOfpcNkM6DG4NE3w7zybaVEF69AVorKej7stUdcUvrDqTE7+ZjNEWeKXybxEcQLER
xpx5WCiHv4XvOKyTT15bG2fVBU2KtcIyX/kM8PFRG6tFstYSvNSdqGAZXumvquJPkmv4enESzNWs
NRYc6Ln/GcVbOuhUjEXDmGBN9dedCB/GVzbt8YmDgsWrrn50usXEzr1UW5oZP8AaB0n1qim5va0Z
jg63VdtHLjzvgswQKD0mdsRel5DWroTNHl8dLUDQzY9f6vaBcH29k8m8nUwQu5bcmD2IPrN4vq2j
PK5CxscIduUt7391GqrZV5WS4XqA9ABV/SKAZchIblXUtuQWWZrE5mZD7/I4mne58T6QNscthduX
AY76BYNOtpKHyu7PRRe74esnfizv9T9ZXRB5PdbqaPBsfFgZuX+G6Tjzpz/lKW0P8aitXd+gu7gf
4Cf8+jSw2ManPsG6yTvQq+BIiRUPNB7OGaq9WToUnrcwsO8uxWS+0nJABlFs2WqlcOvjlllhlMq6
HriCwkVXtseU+LJ32SkfSNaAWcLGMyYDZMYWKNhjiitICOuvpH3dfJ40b2YkQivjJ/t7ByPHvFfi
6pZRAdBzomkayvPCQTPb/ym/m5c0Kz36/msYs7ePb930SpF5/TV3fb3K8W1Jp4B/KAJLuZpuBAr/
ujWxjEhJIoPVEy6dEUuyzdWWUEw9PEXWDUtfp1MkFvqkM0eC1LLnB0+xeBDcbkzpDGlnTSbdp4V5
ydW0AAafWAQzgLDN1nWRdbOz1bZiCdXujb3x7O0qZb0RPXc+KqzDpNVWXZskfzqRETW1CV0FOmTQ
7oF039Shk7FLkEcEwUph0PiI97Yim4tNZ4KgzSN7SFE3OV7bc4sg9HF8PLm/2v4pBVcQ8TEaDgOq
jqlxbYoeHJ3BcSG1OMadOefJxaxoJSTuLKA1wq7QvzM1tfKzmz2m1Iy4FukSmv18iUfcw7U92qMO
eh+xnneZxjCBtq4hnUBk5p6un4emJIyiculfSDz6A9PyM3FFsOvMTLBkVjUG92hqRDz7apPp51ny
YMewXv/mgd0M3/G4wILteYCz3RqVj6gWDtfZCqO8oFNJyjjwUuFHjEM91UoXKIDonPA6X+ZpQIYI
bnhVTaXr4ZTL8WcISMJUydyOOTt77z+2EKSEWy+9wGMyKrHRx+pNEllk0DF5eaqjlNnj+0iXeYrr
GhfjCLsKJ3tc0d5UPB/de+CfFB3onuCzhbgfwecZT/cQCpxC0hGg6PQDbYk12Nc4PAv7RA+ivhAw
/e+KuLZ8x6Bq4mFGy2zIYcYve3pE2UNZadoMzPdQ8UdT4rCbvNEXPuOX+Dvlqy6XG2Hjsn3iBP1B
d/P6S2m401aKy5P+GRKPNcUjXav+N1h0554pSkn9XwdBiveYdOrGjg8Dia4Eh0gliN99Ipf7+G9f
oipJq2XgOLs6mk0U4VN1Vk09lHdjzMqcjCdItMJ80hVkXI/GB/IMkPpP4ikxiyKNqhjReER38lKa
6mLx/bfdkpjj1rASSdBAyqoB3lWhWgaIptfGXC0mT5l4JA9/s5H8dcgXd1t/o20wlTO2PEyxIOR8
Xb3qf3TwJf/FqGEhe5g+nxn1TqrVEHHJNGFwSHWFOKH+LfQrg4Bgb5WI5B6SB3DkRjwi0SsnCKLa
bJUR3gSTkR7XJfxQK17Il3hXFfDXz86aE0UTbHNLPg6yHocTn9pKSXhIfMoULhVF5vKspRAVhlf0
xaiHtXSrvOwIXqFwoC81Mr73QjUiEU4XChdIWgiv5R9OrehvCSG2lpdu+XAckbZcYPPAbn+nQoNu
dZe5pDgytMAP4Mg6JPTo/W7J9+yT5CIv+OG/bSNqrsp5xleebBZnPwrfe+SKPLjqCGcmqowPscpL
/LhwwbR1GvYiMRJrY0nvYD4n83PfiYfbPK4GSblVS2tRR4QzbWnIb4jp/YYyCu5MJuQSy8DSnDXj
+KohwOMPRlNvoZXR2BISjwUvvw7Lh8wFzSuyfbuLToIW8RZTtq9qraBihwotk7Vqbagz9GvQ3Ird
goBXstLkcfnZNmwgcfrsD5rnqBV0Y193jXuHMEnKHkeIFxqSZxfslKdNHxDScu4nAC/Vkhi34/A7
V+ZH8FB6i7HIWNeXLTyQYGlnXfMMckajXtIUlqaBrN3DZ5Tp3HhYztNQ39Ouw+2q2mVuwWLVqHco
zFMNa+y+WM5Q1vE6ygNsa25ssQVRRWMLdvtjYxR6Dyw/upy3DFfd4LTfwsZohe0c9FemaaNOWDdv
pDKf6Svgi6plCIw4p1T1TjaX56xLxAKn9A8tbOhn7Q1Cid8SaNBURewa62EWdETx2fYEkcUUXKzy
oMCiOgKfCKDFVUsPm69Tk2qNajM4e32BEEp+7TwQCAxiQ3Nr6UvifoF2RHF95xVWoZoJbhwgpTEq
eAc/iNJwEmtlkt2ME7oBC1IiF70NrSOpPnfoLlHUv/0DiO8N97oXcNRxThT2RH9lht7SxRwk9bne
cGUz+lvJFq0ltOhHFt1IxVBGlEi2xqhgBeIYgXckyFsSEyBgKYdkonio0TgsE0m8qSoEDMlhccAM
zCgpSOI2lwy7qNuoQEnq12BX02uQikwcdsef8q0q1mjYUfhA3DWLJ9CmLBVUsSMKmfzVxqLqolPh
pBULBf/RvtQIL8dpe1yC4GRL5j3F2l4KxAAI/ql2SkL4r+wxm1T0ftgDLm5sfT+dmwWz3O0yZbBR
Ub04iOh7yucVHiREmBFSCyBlulrearUL8E+rbxpX1iFKIrRj2osupw7XfMIFFfqoeVH7bpOITIc+
9A4pGTplhTjxg5f6C3JuIuizNT7KW46PeQD8YBAPEp5r0+rlhPN4aN5JXUS+1Y2crC4ClzQePpYp
6/+rloCShGEkI/5xlA/HKHz+PxVw8Mxfl1y7sLfb5XArdHhX1kTml73FcqTwYLgLT9MDgTzggdx+
6HbCTESBjCVvikXGgbusYJRIHNJAqhQktbdXFV30RtWCTD1FukGWndnUJavtW2VFbkE4OgFyUZ+3
ulX0ywsIQoTOTH4d9azsxgn36hKwk8hpvYugsZzhuPbD9kvA5HU61VDjADP/Hvo86A1bDqXDvQvj
Lfts16/4h71UnDoSdLG8z61mqOKoDHYIoRvpb/bvbwBGMxhg4yQC1SWG3oTRqI5LVWcDAphv7qS6
wRSCoRRb8k34yNfiYz28WxNW9wPqc81h3HdKM8LxkxabChzOv5mySbUK3JCbfjsXIjBmFiui8Gxr
w9z5YM54TgHn2tYbnhBMucgfp5zp4fluvtQ3Vuz5sjWumSCpNNyDkSBvaKNWiqXnZAdRDR8qtKfT
WJAnHIWUOeNrnX4XDiXQG2hOgYdzICb127EpsTuDe3J/COyQhBcdLNTYvWalJEItkmmapdomgCTt
/NRuqAbBVHv80TDkr/vGvAjq+uR/t58m1PkXYelEx0WHvgki478cO9inYvmwRZIrX+wsZIV2JV6g
KbeJIt73yYvmWV6TcLSF8tXZZeHgGspoNz//gVr72KzHahLh4OPa7j5VFx52KbKH8YV72PhSPVFG
l28bjXBCbGPkg4zStUJVUMoZ7Doge5u9plkgv5wuJ05vO1LcdsvhKFGBgnbA67tCt2zxBdWsxij8
iV2WyQcuW4c+DzEfxTMER3TmqM3ouJ+OTmT8rz4AjdhjQgOyk+1wna+TnHipSfyiZXf7fXkxhVKm
tbhKL0szr8vC2ytbuv0b4/XnuJUooeJuXWLc/tnH6QzzGB1L/DCYj0ROvwwl4wQd/72hKrEH6mz1
TCE4d3bi3WvBhD5X0z7+tYD0aASqDHyPk85JVL/2czvoAI+EhtmzE12+SYqcnbOkA9Gh6QwV7jOB
o3oGu+0Sb6JkcxTUoFEDNjyGmCg+diwI3sE9vQ/q/oqWB68sbQ1nuCYKQUEMiWqdncctUYvSRRxZ
M8FtPrfHZfZS3iiKBTLCcu7dj3Qb1Gdx7fnG30eDAjHYJCpzs1kIzsYruoj0lt5vjZkr8K5+6pc9
A8XDE6qe+MN0z9/0eqzH539obO6Tb+XLX0RcbgDzSkB5wPN6lt1497Y1xHDCgFaDTL2AJQHGl/CI
7QYNUIylU0ZAfPrQddSPbaLpthoWl/wyjzt4hi2m6GBgHFnmycLm00OG4+KcgNAHZICjim8+iu+B
/0ucbwesddddu+H7meqhacJGgBAv9AmQQHqcsX7wUPWn8kmS2NZOg5MMYOb+Yh/wCT8ms3vnOZGO
P8gl54lkiEBbwvfjFbd6YG5Ayt7dYeml7aSUIbaaxKjfgT526xKKQzFz06iwj0M0FzOyqRzHuM2X
zoX7JS3a9rSqR/OSZ1jEZ0a+KuoY9cCEFaHB4fNO1UczRLFLhQnL/i5nvgqDyI9S4qD6EOYMNd4i
ghAo4jMCrgFC0/1RRv2CTosEmLKaO21cHnMfiGnM7nOM6Vt9QUCmxWCzW16MBXPVxV79eBdN2Nor
rT4mZhXeQKyTDIn3CW9VgKOnVROdMrz4XgQS5V+7SVyaS4a9ImSJRuPYqDxic0MnfvJu/0oV5spp
UBD5CYou1E0dg5z/PJbdOEj/06IMaqxfLiF/36nYuFOFpHlPAM5T37qXSxtgBUNRXfmSda6bBV+Y
L87xH7rFI7HYyVozD6klD7jkxnWnaaaNVhk3du7+r60FlwCwYe4q/zlk5wIk0gc65AQ+TPN3oW6j
vz0s15QaHGKQlqrlVbuI3XfkApbGyKBSqwQ0M9E5QRDdM497XELcTYL+sQIfQvtUoTPJrqY4BpsF
9urmf6SBs0eP6MlMTq09zUMslisF1nfCQRtz1orogPgbXzGR9z3HJMc5vYkGFjGZsd1yntxfmF6L
Cw5XoxwR31XnvUgeA/N9DlkOIy1Eq0B96QU/UyDr+10f07fJaMfyZV81kuuKIsAQvZzXD224EBIO
mHarT4Cpt4+cFhte/PZ7qJPz7gPj2Xl/8oltU1h2PbwEdH1Tgi1Q1I+gnDRMS3BiFk+yKAvoDSyn
B5mzaFJpMi31WcwaYRHcpc4VMPv1b5QOofe/aaXSeuDCbrL+XxGgJhstPtTP7b9y6DqwIjbGQtuq
eOe8Q2QGTBVw0FGfSGXQqtYNZGXeez7FxOTVGO46rZo+j1KlP4fnWJp6ePvZd1rkxprxoQRyzmGW
IBUEkmRE17KRwMRak/jbTyWpaVhbyFxhPn4EFmWO8hNh6+CKYaY2YwVMDha1Wk17a365sbCxzZ/N
WhFAaYr9uTtIWikzjeh1PGtXbnHVPSZ6Yg7c1c9EKUgitxh29iF4NmEA67CT+ZFpceFOTb6250q0
5tji20Mn5QXi9/r0MSq1o+FXw4ki8tofUC/4t5dlx7fg3OdXETra5018E+4B56Kmwa4fhvN6sUdV
rXinrDD18WF+1vjerUFFxQJjzvJSRKkMSn34njK+48IVT4dUMMPlHjxecqaT95VeH7DzbAZFR1DD
CdLIrtIgGfx64s13TzYTjlZV7xKtA9xl2w1/n6ITyKgPbVRGAi/exqK6WbV6OsSpife4NPxvJALP
apIqf5pbKu/OhnBGDEqZ7OavUoZH4Aqtq5i294GacNSbYvkOBKD+mhndZiP/BFbSZwLODgLC21tI
AKKtTP5jGGYKQkeUddjSxiw1cnJGQmtchNNDAVKKUezMRUvURD4cQiZG4QCuBLnoU1G56oefJmh4
+JD2fZAx0N4rbvt3EiL/O30Yf6pu6k3N4G6Eem1mMzgffqJ3nnX+dXV3FJrpV52pmLJaGQ2eVbm8
OKRCV51UPd+mJmHli+DXcrnObwXfRYKLlaLFdcwk2/4Vr/Hdr5l5JmPXbzPGwCFgyqi0bVjQ20QP
oiWifVm+yBSsWEpFxosE3FUSWsHzLnjiEsl0J1s9ACywbo2An4BehwrA4YcCphgMicnukZ7zn0cn
aRM8/szZcTFMvd0gySY0Dco2SH/SN/l1tyytbUbp62yojxMK2X7ph96tJ0yoXpUy+dTfbzoyBYVz
+7UGja+vtNpTSYPRWBaVQ/AHF0WLR4ztLWu6aM0fFZoQbKv0Esp5No2lQfWFsRvTavdD3xE1DTJF
EJQFx+NhlUsEuoagcv4UeQRcB+sFZEzDGM8GIdogkcXIEClHPGnRMsHEoLlzIc/7s9/UZsWvxxyE
CNEpUmlscFYShaSjIC9pmBJpU6+2EzJUBtmjKeclgi8a3mdgLszgsSs3mpMW3iiWZgyPSRKXIFcB
GJaOsE8WyVZX5zTq38yF4U7sbFVq3qPxxVklop1s2CMuY7cP/MRp6j2im2V4yXg/cPofji0J3QTQ
/6PY0ESt3mYXCHmiXgRW83P9A3tpZxvWt6bR1KDQ3VfIDyDZjdzuapWQzrm3LlTkH1Qmz19SlRvn
O/Mc6CZbzvPZo4DRVRk7g/II8F2BJs8eSUTk7EC5sP1KhCMHPMCAV0su+ZUaHVrlItrilLSiVLxb
lBGoDN84sPXpZYdZ+vHFkYqYBo4yma/5N9I5y8Eirw06Fh0pJDHeTRolJLXMYdurysLYdo4LV05X
SsbRoyMV60joeWtrO2tbFm376a28aYCIVl9GoNBHt4ULwIx+Aj1WAk5ABVCAm+JuaLPDZ+f3YMSd
Yv0niHsfoCI/E63rL3l+XEmXoTcw74xENGu0R2gVoLij8PVEVffeP6METtsMzj6n98KE/dSlkkV2
2NAJ88r+gZLLqPKh2M+qi4/Q/O+w9pf0FA1GfM0sFZjEtm9/eNwtpxsA+NOKhHevaaly7qQFkNEr
hhQ6PS6zwIR/zaNgHKh2jp0AC1X+uU9pSn1aF8c/bT9wMVdSCdqe04ExPPE/oJVkLwfiCCpzy6/J
Q5BjTOoNgZMMHKmPIKklQ5YKgSq8HlUHTx7zY/zRUxzCnqjQGnZvORhps1S9izqer2N/5sgkf+V4
mJTfl+BLt/LJ17iwF4mgQ6lyqrP8HrQ3KyHC3PELxzo0XcLEV32TcPwfKt7f6Fv7wR5Uf0MSCB0y
c1+FBjfALjH9pLTl/2HCmC71JaBBf6JqfON4fI7hXBwcxPj+GuIDuz5Nu3N+BDwh4eSTSzXLv5Z+
fR/r0zijESwqteg2ElH5+Pbp6YVw7nDVzT8KsaF3OrLfTN/o+aL/HabekQMLrqsyAYasnteJpFq/
I8K9UfIjFWMsrqCRSrxRClPxHJmKaTIdA/IpzKcQ/k0ML5xGBvYbUH6lbctpVE4yqdECR102rf81
maoLFHPcnZ0xbTwKJVkmFkprkVlY36dRL036stpqnVpLxmvOV+H8pYF8TG6WgDTGOEsKKBnENjH8
yZ3SjN+hQ+N8yQEVudBoDV3cOqioygon1kfHYk/0xPZoE+n42dm3DDGSHLWUlCtBInvcQHNgwf5Z
Io8JhSdq1GUz6msyyuIma17Q6Hx7SHVMb7JZH9ZSj9TYTE1vadztrMLQfDTBlCF4D8Muoow/4Saf
fVdtUY72/2/vFPcRwzCptIbCs6aFcg9qWk7u+gXqVXGgn+H4PGV/6foXaz41ySg0M2g63pTLC245
W9rV8EYgFUSDZOaFsHPVbCcqPpS+mnSJ0BT2KSCrU80N82YJXKoGr4dKiwwViDH56ugLpf0Unyuq
8kn8MF7LXp/M91XpNKvMrsxwgrhyTOFozOho0+CQMpOHoTVN2KflswYKRk2ovniC55VDeAAsB97T
3POb9S+eCoaHhuiJtByJfOWFBjbOGCidTS+aozWNCy+HdrD0yOhYzylQ9z4UX/2VpEH4QawIM3HA
JFQMneh2kHm95NW+kLivRtDeGRTZhQL6ye+vbXaeCmFtlQyzHl/rga5EZ1EnTI75wnxKMrAGPM1z
NIpul18QTW8Md3/AE4GGIdLuvY3QzDpetAHSJPD4tDPNNJJmem7JrXBoZpFQLAR2bIpt1myKGLqU
8Glv8WE+AyM+wD+o5VF3+yQfkQ3aVlxt0X2TRXLxHrbOk3pwO2enkXWnXjpoyvg9hbGO9iLWafO7
SF08d64Q+uRbjEXeN91PQVKI8DrzMk7h0wMupQBPQAZT0UKwVHIzpPgJ0xVaL8vaimcDisTmqPZy
RHGzEeWj6WBDGthY1To8p8LhRR2Bo2E2wlhOO/buCQ5GDcu4hRtidKWTlozUN0+VnuTODpcAfU7d
gzbZqJjIlnbpOOsYn9vNlLNp+oJDUO6rZ1aMs6PJKTocVJNszBG0eoRhTMSEJ7XPvTeYRYt0UFqL
P5pzqhXREc+vouZOXEAcRrHrPMZiLv9IynKr1ggHNZjsB2sq4Bx1stqYDMeLET7wuKodU6L1z7sT
tQ09WWiHIAAV/8Cf4CxOYCXKNO+1r57PeA3+1jOo5JXu5oVS/FH6KBMYsnbxR+kq6V60idAiiBsx
dpfdJoFf5ILuvdXcVt1r9W92UCPHBlQHd2Y4HZiBFtzSAdr2fzh7TG8SVpWbnv9N0frB1K3IbtJZ
b/dbS0rxGkJaE1lK0hw4DifVl6pZUOXLEYVoAo2VFrXzHanxPk79r4zYbSAOGPzAuJbscwPXO5n+
XM/0nQZZNbUkoS0hlXHW9HPjclh0LpwXyMPE1HVadcxHrI0gDvNAWrFip9JnkPVmzYueADhoo6RS
Wxsu/HB0a8Np+sRlxv1LdU6ds6fRkphLucbPq3+fao23P3qAtwlnEjSbojP0dMZF/TigFlEDA1Cf
oihrjk1gnMwTVsP22MmNnFhGz/kQsuPnArsCj6mbzk8BtEIu+fR8P6TXvZEtG4yv+gSQjJM+z83A
6/oLBCC4pYlli7tckRbR72C1w464aKh2jVaFDDtjNJCssT7uE3OG+LfRs42Z13WEBr4r96uayIN5
hZ65SZ2VsUj1tpJ1Y3IKIwnS6x38zRTnEQT2ffNlEhczk8cdcK535CvkoudpFYynXzTilS9PU4yg
wGRyfZuCf3zHKmEL0hfu2t2v5bKH21ymmmOvsQiMUpZdx+Wcv65aSnpYEzIugZSR2hSGF4acIY9l
1BTbdLhV9LVpMXC0MRWZvZFkcsTGMH7DnONtsBHh1t3sNDErFmlTuqniem1kqpByHB1NmNKHrtSM
Qz4aRjRb5jkaOw/xbZivDeqHrJv8zHREzTi19cJV+yN6xbZeXef20xRe/PGMvVJqyCqUcYXjPoye
fcEGYAH3le2m6GVI6ZVNF06xaQGZ3b4o2PEXEHi5WypAUFsjgs9wOp1UzAq57cgJBNWuOFMWHMGX
nVVn3rHjk0vKVBU87UE2twG62uy4FydR0EE4rklbfNUrYPTc1WezSHN/2xutdiQ6h/JDFW4LCpi9
M1frEPmHzi4VGVH3YlkakwNXwFnIGbezqmG2Gij+kxpGVxKeXGIHOlF5jwmX9XwdYLG2pTLS5VUt
9ZFjaNcjFFATyk2Ky06tIDpUn3attEJeSZ3aPQc8wAgtn8aXyiprAQ5TN7KYYfPcQ4zN6Mj4OqeP
Fq1itjKq72OMo/X6hQju3OvCsS6AeHxGo3n0WIZfA4fmz/yitgDIujWLw5WK1ILt2tghs1hMeIWa
xHai6AW7ErDU2p5PrHvYZ+DBHUmZtThBOgd+ZI3zRCMWWWBJzlnRXG7DDVl+tVF13+rUDPU+jRp+
gRoa7WRzF3hGhzcNSJB7dR/btkGnSPEw5YpEvBF9FSM+WewnMPk85Tx0TfKY3xeOb45v4nu/gQml
wRL925oZHZatkO1WGj+rPg3Kic5V8V0I8A+iajWKyWNUfzIBJXIdtyU4t0ArgWcV0i2+I+Vc4LX2
3r6hUk6mwg9IwIkZM0bt0GtyyX25jAgJjY1cgYRBKw7B7c5e6KSjQ15zfZSWZs/5dSDRzjH6nn/c
KLmUKvq9j1Tsp8jAd3M1bhmFVocJA/c5gCc0FwZCUIOWOUwoNePXYvx94rvzyWkHWZEIs6a9GMRP
1PUxfWCzl+guIhnpnJnTLh5HkWyTfwSKr9fAmLUjSjzLxlkqw2UIvz807dIwyLGET/Z5GpPmhn/y
bugwyJcCWkFRcHy3yfbTiaUVRRPg6QY/TTWAscSp5nmiDYJGoB/TX7pVQK+hl/Y3A4DrO2uiwDPA
Mp1Pimivo3mqwXoGMmh5aRT1LGRImJScacHj7Bmoti2y8ClKeHO1DTvWkGMykx6b2Il03zAg/hUr
k7HQMf9mFDj+m2cJX9A45m+S8DKtaq4w3KZaup9OQ/wnOLEwdS8VlxkzwuijeFE3ME38TcS80FXu
UIJV3CJYTZOW8ksxIxVKEGZuzfhmY7jxqw4n3CM0ge+rMo3PKiIS3y/Wznw3OjGNZGivQpLbB9ya
6HFKp7qOSNWfmWctA4rFQGffKDDc5oGtkT5BALCePW3QNyvh3EKjpydadcOJh+wP/Dmp3wFUo+ha
obUBUlgQeFWCKoZNIQg0pXpFI+5q5Hkj4ejAXfddH5G0V39ddOADUvnbm7p93NC5TX+9wnTv9wO1
n5EOyA/Ajh2hTb/8jPsLWw5JtbeP3PZPMfSd70fFSAR+irpl7/s4WMYFJhWjIfyuIGMXkCt4yJm0
EPQRqvVgQpGdtzomsxze6TYecd8omD+qw5X/VIXq0HDwgfv2UaE/UZMlsF1EkE/5751V4Xk8sHo4
BLpzNk5RTmIbBN9tHN3HoRC31Q+DYjWNjBr+rl7WZpoAw7ECphIXjm8NbcJoeFGZtRnLgSM6tDV4
7R9BWljrGoBtAsf/QVKhuvf0/fqv5EsHsp1yT4kc41Wwh7yMMk81SCwVeUoNcWp+VltizdG/bejn
6t/yvCo9Im3BpsIQXxylURa2N5wwObAuVixWIlSwmG7H7TSd9Lh9TjrisuSZvOjCQa/9oA0TJcuA
vmxoWwpvVEA0iyNDMnAyqW8CkmQkEyE9djdwjxnC2D70gnFXgHRMAvbcfJH5VjV5Ji8z7QDt2SAZ
7FajeCpRvBxx7yKX1DtNTCf7myAuGfCeCRKXvX/rwuRj7Wql+3Lc4sKPNYs1iVTO5cioRPD/YkCk
HK0qqBVdYVbZwMaEEaCTQ/h3CZyR4+e/+ERWSth5CvxK4uWXlplnUwFStfzOkpp2hvn58dscXdQ4
BwfGXlNm06TSFRmYci12/au/UVuiFS2tfiMhSi48Fe8pro4KzxLgYv6vEr0QKFRH8tn3Nl+C+I4D
XrGh09CKgwX9Wy28ySoDdAzmfI2Rt9XnyFJ3JXTjUgRQvIde5fE8Vjz/+Uay3CVy28MyHM/NHHFs
Ovzo9fNZdUY42kxMjUFUicT4HJwtVwo5NbDO5smF2zleifWk8a8xeZbPtfjbLZ4XnqiosQL7EtTX
v1r48jqks5w6lPHQI165VTnzrt3vTtAlx9ij0SmlQeS59OztfEQJw0XSUCE6L8jQg+QQstNri/Mt
rUIrXZaTQrhMSduNpETYvjUJFCIxV+ZBqM7HgXexv0Bze2vwJWHTJ6C/1tJ40LWCGAzMsjXsdkXm
TcsVapbAPevG3sEE4lksxWxLpQ/Mk1FMGkRbxpoddPYRg8jprEDRB0kzK7CVgD1effJSZWpiVI0H
qmn3AVZ8V+cosumY2JOQzByAIfZFqtoP/LwkKb0fc/SL9vG97bU65A3XPw7rd+Af7COZRL1TrBPV
xvHk8ukkXH7/J4+LkJvZLSTWlK4anopYrrOM2inE4mOF/3k4KzSyU85QCGRr5NVuOXA+kLZa0nGc
x3riz5LJUf8xGTNcTzAvbFhBObth46KJ0J9F5t64r24aV7zXbXpxIEnMi8Z6+AroCAkTycFXEZg5
sfixV6LKF3dCnav+psknxzbYmujpqN8gZpAgvZ/O/9iUytaGuBBK9JejwZYnyyPraPRBf7J67Uh3
z3g4k07OHXVAlxavA+s6qmZUV0j0RVdB4YF95TE93fMwnY6g6+JilUDsr+lzVb2rKMuqVCcVwlNi
qF82XzUWfV8Yso/RmEatU+bHJaRbnH5iv12am8XWMjd17uAvPdS5bsPj0ZGI9MWdBTwO/8RReZoc
0tmgj1riqN7EiZnpsbZtTr7CQDdZwUdSCXWllYL6JZxicIAM1aJw9QXyuwpj4kkX1rMu2/6lp0XN
cs81GN1ly0eRyt4i3boyMj3bddxnWjWefOh/OuTv3nuF6u6b8IzTB0sFlczdZH9bzWcQNtM+4pmt
JRX+lAzPQWxflBtPAkwdW1sWxacsKEN+RiZE+2/nJK7JD4OUa4HSKFbnDTid7llTGJ718uX4Hbwq
W9y1XQ4IXFc2nK7XGpcBMqUAw47HwEMKQuaO1Pg1wvuDqcm9Y3k5ku1b/oXURjEYhL8+3A0PdTGn
nuiHeGdrrcEcuWQS3lgp+6ufCq7psEX3OT1HxPAsGf+AeY1QTWyBBJs65eXm0nGb4ojD6P60yETi
NSJ7ScEcz3QIYMgUMibqyQtetsvL5dhk6EgoHsRkSv2ggKWEgzHHybBQ0EIT02u3BZNPUbb0ORQR
BIQo1qvL5I1BuFMm7h2/kkD9C0Iv2xHZ8QTHGY9sGgnWWLZbZKuBSnUqHsPSzipKSxJWwltl2ynx
iPp8ad33l1NsEolCmavnGhuByFgWte2Y6kKMGjKHpbPrLr0VgMsxrprhPa4gyAj5bCvDcJEg6K93
uBzybcFkOwiVgmJ+0GWq6sEJuR/WEMormt7gQpYxlK8AlbxJ8laJJzIdFK60cRBcbMEPZTF11btZ
yfGB9n0qmzw+DINxXma2YVrrbtO5BVP4ANoDAOnmiNxqVyO9RoNVpYv1a52H91bVGqERgtjUKr/i
22BqCBxjw9NuuzRcXZ2MQPXSecM/DG2m2AuxG54gXA9HEeckL6Q5v9HyTQNF+mrOzoYXFgHHRJbZ
1737aY5V6hBhTFnp4D0A0xCDPcZLlCKkOJnuKG96iAnBFBqqTeXM1DXpPjt1ZIwopldFHrvme5fP
Vo95kqHDufL7DEW3VxcN99bZFK7kT6MpgmfhEw3go7+Fk3MhuPx6glGWTddfEA5ymKNH9m5JNCEn
hU4gI6HzTUwwreolLcCcyTP57bXeGdt9BN9nBvFMMLkMFHEsDDdqEgP+dIzzxnlUGB1xy8bQ7GYF
Oh7+s1ReT88AbU8nUcRi4G1rNnwR2zg0H8WV8/wcgL9A3Tz/8+WTwbWZQprqYrx/FsvAsYLLN193
Ik5MvHt8lI3eJh9mx1tSthpzQQuOXY3tyBmdnxAR2jMM2M4heamb5LY/VI7zb09A2n7VMbo6gIuL
2w4Mr4oV+WCaReCswFFdsDGboAk5ireGk/VfKvG6SJeqnwp3rpr3VepXpeOZSDrXttFwFYrWWc9/
4DGyhjc4Vq8VIWJWDpkmOOPhcZRyxrWcscE2Z1n7D7+gADBnaZjdcBOFnKBAXzm1JwVXLEtNGj3R
0ZlhByHfFQ7O4Q8bkZl+54YTohxJq6Q0dK2C/+J6Qr7sWUdMIkvoU5nLjoTOkKxLMSAgvouhiJCs
6E1N5KtduHlDftJj0Afxxd97HNpiGm1OuUeu16E04lVWODfH+uVL+SzwH1BahWBKKRQFOV9FcTtd
6z2dPw4pJUinqKrLNp9VCXmVOBR8PBeRG+kKnL27MPkd/kP9W8D4I8HcxZkFslD3/5u3QE7KU3mU
XuJaxhqY6OOkQKHw2OCdbU3XaOgmhBo2E3a/gsndHxvisEsSEWa1ErdZRHX/S2lhF+5dzY+3ON2e
5o4kIsQzx2WF81ZIlqGrDJdEXBjyeJc8fkTF5COEOD+U9EXItfMsBmyF2d7qWHsI+DZrWMKhq2B/
GpJiP0czXdP+QWfHNB9iOEUEJvQ6STPYNJnUQx3fBUIiPewUqbbTBhHb9cxaYv5QDlwfJcu+nFwQ
t7Cks2eDrxZvpU4gvmboRb6EvG5is2JoETjAZZOqeQxyqOHkxyu5ltuwurweXWk/tGu9uc/lwmSs
LhjsW0DplE37R0rgr7a3bi7YguytI0adYeehvZyYo2fz+VDraEr2dFOAuh8T8L7vLfrdDtK4TUXl
NK8QVCu9D/ILF9vNz/Vh2og6CzHQqfhsSdcKBN2AtQlSWCqJDHFms5rRqG4KVghG3cMfTurBLpq3
YWUwY+URU1M1euHjtHbVeIhL+wwTEHxKHjHtPzimC/lZl9+sbbHJ2jDiBZiQ9Ci2ZLv5Gi5HbIdX
sXSVe5NHOX3v82g/ZWxBzQlgUHqkKegHf55AyXfCWcxrCHfl1cN6luew1crqWbZKsl+M6hRpRUyV
zXCpTwJ+3tNWmnb9Ip6lJJ+qly+zvASnFBnXphVwnZEqIJMB35BikRRgDgFZ6HylhUDw3WqYoVT0
eIqVKs6NaWU4+ZGC00HjKEuvJakbYnfxo3G87Zlu8cQljd8UIAo+sBcHSbF+MLLcEs5rPaAbay9d
EWccMrDb2kddWsFtVeMv/7gh/K6ipyEXZCqxZyx6o192fDldD+G2rl/217YbAWY3mxMEgbh8dBXS
rHniZ5ZHKFXO7wkeCyZJW0eUD2ubgam105uO4BZpBkEmZ9p4n4CHP/agGVig33yMM4OKcupr+10G
2kgxMz2TImNivS6ARK4IRfCvnIjQF3Hm6/cgACUPWu0O2oZoTq+v8SayL9kd2C1ojTYtFeiPW11K
iXKA/ObhqHVSnLenI7xOVXgH+WtOcit15o+e2OZBm8VXZvNvc1axEGnolISsb29EeSqUcTUoN/fm
U8SeJc/YBYvah21Aro/ljyX3fuWIf0g1bGyDaUJO/5qSDrYByBhoP3+ZQ5OVGptrVo9DWuPEuzso
HV6FujrcVopVWaM1nep9muU4VAqNG8rZsWCtLOzpNTcUbp0VL8Qzn5EDhqTTQEreyKLycKCiGVvx
2CYDdWsAoFOAsrUhKar09uFWLM8XtjASmsCtR2hm1Iwe6+TagbIME2sfiBYtn8EjR0XXzy9KQV9k
uYCIdI2uGQAhF6HLnYuyA82MAvw/rM95Zm7eUhBWiXRE0QOdp5R1ksYspAqMbhENtXTJwxc13o0r
rG7nfizerxgz7i4cQIBnNm4HX9GJaZpghkWFCba1H4as31RvVxG5TvRugejWS6dNYJBBQt+wXdEb
47dIwNeFHdnR68JYEG2Bv3liVnAYRSirft0PgjY79/yHfdQ/VWG8R80HasCKKD74zVMVJSylV8oE
CoqZVsmcTE+1Mz/q82aVvhMnFO19rSS651jhUys8SjnzaRIKESIQB7dmfCDEhGkcMjLsDNGi6BTX
3dBsHCXWH12ZnsAP/tYUDi4hRA0PHsS1Y9nzOT27ikLFgDq36fc+ElqhS/5yK25vysM64vuXYm60
O/XYlLYVwDE+Jj1XjLgzItPM2129wX+DD6dnOcqQ8uaO7Bvk5UUb1WK7tOfti3T154CaY8lHuVf9
+4zNlysuuV+fKE7Z547Aiu5Ok3914QY17t0RA9JvBxxhezgPz2u/ICOr3WafOWpJwaQPybtCj6d+
cUF/48b7q4qziQDfrPjPI+mIzXt7wVyrlY1kIbi8BWd953zOK1/F97uKd/lzwEJQN0+0px22eQQ6
bPnnGsD6kViAezsBnQKkjQrhk/PzcVZE0CYfLfQvoY2iOOz3XiL3hMWJP1ecGv2lH3b7XODzWP95
sbHHmUaoygxyxH6R7d/BFUIHuQAQTO5su8qQ1tfHIjvVSawy/N0q6ZAR6exis0vTPi7b6eYUfGwe
FwUyV93oP+5010+fRowCoG81eKAmDz8rHqFQcIjgr6FHhJfzb4x0yMgUAG0ShA0/Lr+U3CdYBiHR
uxTmqkEzG9YBQOhaDBzPOKwNUrvTuz0iNkxHgJJqNze5yyXuwUAglXb7FZJPkRX1R7lLyWtP0lcw
tW5C/QQ+bvHsnGPEQZFHCP/iTf0il2bSG1xEY5+lgVHSA7dmGGoqbkVX+5EcUhu7CXGs2aMmO3HP
tQTPW/02PQHh7HyaaSa/+6azCrJznu6UbwihzooY7YQtkVBAahw4XqzX8ncdnSpQdfMrprsBN8QB
Y5xXfVmSPFdpYV9/22gWadEJVufLofPLdMejlUAj8jR4f3c1NZk2LGfgrMplQkjLIdw+IH7Rglaj
840YfRric57DbltDuS2paVVRKoNAmYpeyktDh4/Sgt9JHOcOrYiUAh6R3lo9GFuoWaZA6IF4weTH
ZqiJvkx31bepDfgag1ibA6X9T9nBfiqvYeLY8HrLc6QnYt7wyBbeIzqAfQC/L5OASEzbcGEw5lbj
D3yFsv9jVo8CWG6idxg8vgwGPadngeX1TBtG4pcs8bKeCLfxJBemXgXpapv9XuhCPRykozkteys/
VxDDnkKfD8O2m7fO7qqMDf8zPQq945A39pXBCHa7LrtTuJofs/tpc1na4PpFmbFbNTbHIn6yZ64w
kmp/cS0SRCIeSPMf42lHj2Fu4nypFSw+2jXSItQuUSFv1uStoM+CAriCt8KXT5KLZcNfA+h4QyXO
+j5HKt0Fl9nR/pIajOfeMg7pxxm6sUnrU8rcK6sEqp8TLaGaU/PuyrC/ZPo/eKtlHWLpuLe8JiSD
3OHWLq60x1v7QSFJFOKUpYFPVX/ZJUk6VtMBXnUN0hJ19gxuS/gFEsHwT8tEqMNUbpQlNo+/FVUo
gDNERRSd076hl3WOix3ZV/Meg9GPYLu4OeOvKPd2arp0Y+KAONzL0P/FFpsKYvOLYMjEu0OJGfQg
76WY1c0UMnik4IA+exwfrOV5Pc7DFUJ5d11OKYhPTR2ecGNYS0gNPKea+qa9WvRbfzFrEpjFOiGx
xJRhQMkoMM9VWyzJeHN+Y+FTDJ5K5mqImdBqAQ5Z2+w0X4fhWQBksv4NQgyn08xCLy5oENr9IGjr
1i1zQnIzEegyPKsYoHR4600yiTPtnaX/JZ7MXxk2E/YAM+3gPhmmjMYj0Q2djRXLOoXRul7OgHqp
nWkiMxqgANUjYreAwMicK0s3V8pX1Ua/cuVFpRy/Cdtw6irLzdb3TERUgnU4CsJmmaeq1vB145qD
y2Fkuujy5ebNvXMEOyJKT0LU3jpTvvAd/86fbfw6RBYMDcLd+85mr0sCG5rtm9ry/ZF7UJmHPPXS
CZpwdIE+QugGTF18t6d1BXoUkNhCdXGEdTH+kMUGXQIs6W8S0jBmp67pfpOuApGmMx1HaDvjo1mG
dmqnLCjMrw4SPbd6H6T5zM8lnlDSaMl6CAc4cHWrsS64HoWCY9b9KZ3U3rcOgq122e6co+R7ZY4E
mSTW3EgL1urRownVW0VHRO/t39Wl8+YSBGy/nOUo5NTbcly/aKczN1/KsYRZ3Rw5nrm87p68mmv0
Nm2qmJ27pRowoLN4EijbuX0Y/4Zxw1vxi4T5M4uUhUPcQXmwh2kXATFKtu+AaIcPeDyhsC1H4AuO
VIn0PTLEx8PoKToV7gDJ38bJMa7F5A8CTjda7TSMfNNVxhnGUUWW+E+dVdDMrHeKw6/ClVe3jTBR
sNtM2HInpCTRA4lpQQ1m4wM1HmAxQVFGsZpPsPKz7wN0j6bVChGuMMitPezvJ30cAlLeU/S6i9lk
rSfLTczxrbyFrG63P0vuJt4r/gblF2Hm/8IGadYDQZob72Xnwf8FG5IrfiJ1pmOxJ9sNtZLrhVGL
I0OfQDSuaxB6vj6jFIGH8iwFgPMUrdvCaNlJ0ns2XJDYpLGFhTFZxH7wD3yNaO/032yXqs8RGLRM
DcJ/estzCl43obR790gF1BMdVdJ+ts5P18Nu2hB3Z6V/Yk0WE5nWkmRMHdjOIPUWb/d7dCaqX+Hc
13NefNcI0BAkwmkirXPe6Z32YF8HtBmzdlx3xT4XfrJdrP2maCQDbvtXgBF7VNvp8b3jhiQ3VHSw
X3ftvz1v2H/E08heEV++NXaBn76O2zKKl9uuUilfz4zl86GDX3/J9jSKsCtC4KQ5J69i9SgCl+nw
ljerV1ixEBgH9TNtnkMor4Gsmh8yDirtGw46/vo0eUV3qJJFcgUu0Oo/V+aIb+06fn0pN98Wt2hS
/T4ShHTnhD3bbIcYz8KzEK4dhX9hx1g/CCL9ubVYFSBqEOvQNNzCGLJr1HWZD9WvpKCtTjNIFtLZ
Qon+6JemfWmjc8ZYsxCuoUdMw8aO1EwfkaPI8lMVHkY90ZPZdhyTz+tarc3x8seiV+wT7CFp/9IN
aex++SFRvONonHda3HV06C3sOkCX0WHGkiy/2kx8WDKYYb9e28gptK8666zEQDmSX2FFv641kltN
OmJYSdT9MnC5ps6SzmaoHVNy+ByXR03daG/2mMGj0RJGvq/Thu4BtAbtXKlK/mWcTLbJoNSUiTQa
7BUYyp7Ui0lHD0+ioX0InecvPORsCkr/f2rKMgUkNA1/8GYV5KMpBQ5GTAHm/YtriWZ7By/7D20r
ToYFI9K64jZU7U37ll0+lMiPJbRercAoaJzBZPI/cieS0z7ukZyjU2OqgHcClXfGXuM1ZUJKfUvv
54pOBQ2JaaPOdFw9TEV4/DnKff2tf9KbVPjXKK2iB3nOBg0eNFvjyC192mJbXPSZ+q7fLiKboari
++Yavghxskkl4L8bNP1GOItNk2ShVjHPH6U+OI7bY6o66HiIlFP95sVl8has3TIcDFUo7FW6Fbh6
4CQB9TWf8g7RBkl2ceIajgyRk6hERrZBL0tSvWpkkB82IszotVf7cVdEAs5QBDJzIk/QJaUUQKqQ
BWXvmpo2q3gAYB29deLBiSVOBLsOZTh6CktZ7MCtLejiXJvrvbv3AhzKyGSv4PCHFGtmcqxVZy7b
gGpLRdfdPs9+BpOV3QrsHyzdCsNTZ/PImsNCK694iBcKYQC9x0eJxDwm0jwtY39fLW6YKRHvtTMj
21ghOlOQolmkwd0c/ZzxyU324+Zr9QIuB+91PW2sYuMmhVmyxVp/t9XJKjWIuUVYFcRRuyU+n2pv
lROqrYaGoA1Vt8iGfhqdhAUntt5qjxeCOzKORAsi/C09PfBzYGlopuKxfZIG1306r65DcNu1pDoT
1o1TKHGw7aE50UZuowweiuYOSAhMWkPmmPMHQO8WaWFaU1vvrebII2X8gQCZyVqgVRXRQ2eo7BdE
fUZO0kPKmU2MOwZgH3ELiXAkXayUEvU5P2PsEUSFM4gpxeNObBcxrMfhrKFVFLtlExwmLef8EMmE
g35GaAIuCVuZ7LyeUivP5jnr+PlgTJtDBk7lFkSJS4hbv95w5lsYxWHDM6d1fb563kcP97lv7UJO
rqQgU3DN9RJVOFwAfNT9OXjOixnzU0j1LqZJBxA6Swy8GBnVnaInyOfqJLz6oj02Aoyfbu/42F1m
sFTv6aVyFjyzxgF7rP6DfXR79IL/rk4jJdEbr+36lJ0SLsBejaa8arrfISit3NaKqdCn9sccnXPB
xf5PRIXMpGR2HrNzcV9un3K6gckoTJq4d1Ls0K2qk2315afECoFxCF43drKvv7Yguss2zYgV0Ooc
FTjpoCR4mCp6x0+gnT2y9URomZ2iim1Sb/XgU6pqbanUmPO3N6munoCxckOhVul9hkB406uIM1kA
WTH148x8Y3ziq7txclegakz+e29Nj+WjZ2+VmYFsebu1uLy19ILRx9t7gyc870mk1OfcLNkW6uwW
pKlZlZrM5GAOgqRM2cdlRPTS/JDTPR5CPw9TSkA2rXY9goUubiiW7/djDtYgs68EgSn71p5yrFAR
GhaHP+hrQtaJa2IAkJt+C1DCcHoIpKaJuNQO3euNELSvjklXBdOWxdcRpqHHjlUpcc4mVm+VpIcu
bMAcQmbQI1fpLY9X/wZyJpdUUFGAx7IoO3KpJqpd/S5ET9Z1v692ux3QfVMBED9GrLIUgX0+HJ1f
1uwRcSRzOLS2QaZVUORMCxIZl9QKePqKinpFDNBqxn9vxqbdsHLlmHKhNtUxG2YVffSZwRCOX76X
lUxpMRpMdklrP0JCs4bved3h6FXTfGRZKcSS4wB/j26WsDp1Y3B3LP6bIHyEqokYWNvhoEXQhCVU
zOF6PvZiTM97qqLvrzAjPkxfdFX9dGnt8ItwWk1KITdP5bjxC2GWUg5oO22ZeNbSNhdKNLBuzqfu
Ba+oiH8GmySrj7bJ9rBXzlJMHUb0kumk5zpm1Ztyhw75Xr+0PDFCCLll4sB7ZBepsGm3MyYYbxk6
/SOZOiPWTu2yXSq5XPqzqNludSCOvc9F3cH1bGCvLBR5kxsDWZDTUaeftvTtij2O0VaMh/3vujNm
fu32+DeVt2j8yMZ+lciNDarCz9jd0085fqD2Ty+nWoMm5RvWIuJCxhQxX/QOEqxFniG5jyt2pA3L
skLtDBOBrl3ogTn9osG3IaCfGJYTWnvALjzBgYLkgroZRO0YJx/2kdcZsSwPMbpwCmX7d2UHGpW8
iNOuTUBIo1WkijxOwrkkda5BNp/XBNwOwXHlKRnOCsE+huZAbKdcKiYvcGqEPKW1lmstBFCw4b2x
CVf59DlaijAkKuxzK0cAYC3xVUlESfBYoenNrF6kKyOfU8Vhz9TpSoLSHiOHVw/JDRRdnbFqBIfW
ZmRXHXz7tuQFvhCeZ5g20f9qWkwfIjLnH9EsrcJaAP4XiHqCRl5JkJWhgE9/3kY2SPXF90kr9gHt
A81WXsExUT48/qr5Bv4HsAEn98CvIqpIqV31/gKItIdoIAeyoNaoSrj7sSIHL+XvopBkCga1Mml0
e4uhd1wH9Kvzb/CSk2hesF0wrE5IxnVkL26n4Zu4edFOPQJbvIEkFcaiUBLs916184rbMFr63qp6
mJ2oPJU8SAgEf+O7bIe+dnRlMOclutXX/QdR1mY/6oIZzlBT/k+r7F95aQgBvd2HR5gVa9uOnvir
EFx0GBvj/FYgXyofmvzm/XlBwS+t3xYc7P0wKlivEOkA16b0TB6Zii6aXftzWellqwO/wDREOxAS
92JWbBIhagFqlAP1DbF5uo+aD+Bt9/UrC7Cd8OORaVGl37XHthyqsxwhA3qCLjtcLocEEn8x9HHk
uB1vU2JeBKVXCEY6wqtV9wVeGkYuqR83qXBowofqEBU5zRUucQTbVCJL3yFUgHAm+ErtJh0Ls+xl
YO44xVSwF9QStbX2K/161xq9GEv1eknyf52Xaf3xb4v7BQHRWtidNCxCEaNXpR2RB9zpnb4JrvuT
H71CueQv9guSoNexJrevN+kW2qw63/74YqdUAVldoQnimYf6CKKFTR3bMyE9HXA9KE6y8eoqqcZK
dk2jkb1BxFTFLH+iSdysTxJ+JMDohJN6f5rjod//Y2YslsZb9etYXOWkXQYcz5a6ie8/946OxFbV
ZiZG9mMemebjjRpA+zp+3ibEpAVjKnLEg3iWUFzWYnf86o20JeeGxKYEZvpG1VAcn6w2wo1Hi8Nd
CJcCsDQ8Kj2ePZklNF+8VTkEilBb/bRbULT6Xtc6AgyCRrj4llvvUqWBnutYRG7b6Pwuv4SV0m5e
wUQF93JhpJF7NwRDGSLMTPfmRIWgRaBYLHEW1QzepBqqD/avWX7e9wdOUIMt/q3ixpnYJYfEJQCZ
nFlroPuQTEENQ7nfN8rly5tUjUp8Brc52UkscOPsANZueRdIV8pVa1d0KYNunFDqx+xsn52TohU5
EngxiOEplNRs8mMLBONYcE+aSy59VVa52yVzJXD3PdzyqTz3BF3w4NHo7QmZsDg2H0G/SMFGGdMx
YH+ix1QbTHti7q4Fu1zqSdjxbpdixU1KpRPZaqFvc8NCtUssAaax9VgH4lL7moJRr5Uwa2uHnWy1
U/lDMlmjoPcpnwO71evbHk4Cdz919yd+xTMc6fe8r3Y+nJp80Jirzm7+TUEOpm0kyUwVKEaJ3VqF
5b+ekAIvixDDwaIfe4vsc7vENTWYDUEvvhmLGMR2ZCESVMX4KaMyD/QX1w9PAhPmJFu0W/oLziSW
A+FgoxCjLte60u4BeIAgHEkP6bTCVSoL8qwzOo4688qtfrwSwZUipTwSbdTw2QXlGM1WzT+8mTan
3iwRB64iVgNLwYsGjirCSsx4Avxihwxf9b3oCsXBXNJBGQ6KmFCc+G3qxd4C5EUcv9sirCIEFdPp
98n9m/s9Dq53FzLl0fHWfwNnHkHBXl9toAJy2zz6Ztywh7HshREMNRW17FDD2YD8ZS0ZB+nFnvFc
WPnrGUuBKBuaAtn6mo1Qe5jc1a8WDhb9JzK7NtCXiuOZ2YkhJbZu+RJjXuhrwFcfTwbAtuL1VOA6
X6hPwcQLS3LD7n7T6F8AV4c9z3S9kx8U+fVugXnycLROufK0DWq4hcj7y/NFIVTj5WpCyyszsH6R
pX2fWDs9W60UZPkJHows+H6SEJOkth08/MAGjK1MNYn6/C5tw3oEo32NOkxp7lvpIMx+gt3/jFpI
0KF7rhEcjbwduZJd9VfE7+cDtpVPhDANJrlpyM5gYdx3IYVUIiFovIr14AuTUNOeXM6+4qEaetL4
FXWC50K9bNw1G/K1pz3ud6Zh7fxM25PR0n3go7l5LfvBDt3iTKCpQgDSD9Yggtj+wPjzXgfb2dS8
PsO9I4yDTiTrNhCrNtDHJar2Z2UahIHuCTfAnOCs9LI11FsBF21li9L6Q/bkIU4BCe8d7Wa/cwo6
bFa0SG141g9dt2DtjIXpr5wk1pWTKVIyGjiy3Ef+pu/vieoPioIa1Xn5GludtxOzrXrj3L9/3nxd
4i6vWitTH9qh2X3itfBfQbqvbphXlpUtJT3+c1w8tIjeOjTlMwdpqOFa51xWtbvh4oxR+qRIPLiU
aXZSOOLm9P/02UYgJ2RllVQCBgLjHa8QReNZ1b4HGgKyw7vAxhng1g+PtisQLwbKyHMrwMFI0skH
1ikUzADrE8c/RVu2B+UrHCYjfeTP1vooA+EqDz7d1hVoWYOc4R+TNXEF6yMCtnc7hDw6UlAk7oMJ
J/vTozvMph5ieXOd9KoQPOcXh51vMtVnayD9uajNvhluOCr6LtGHWnV+HhaJiVlWUx6hdTipNTQA
reyl865KKW89vB8yzWN6TAb/nm1Q7y7RU5w6Vtu/MB20rEtZNMYSTLBfWs7XqqyKwX6Jc/HWJZ0z
D/leFAjsOndTTjcjqPPRISJp8a7Z3mpFplc0Yrc74UbqGIHC1LI5/HtvZXRsyqgVhhFtAIC/o466
BNUg67ZCO0FQhuUHWyPEb2E4EwBDSJW7MQ4fYPeFTY69RAhj2EntK7SJiDMb7F588NizDkKgcuAs
7fhIOalDWXRYoPQGr8+Sr3dRzEI1t/CfSoeElWB9vXAll22xfr/eNB62Bjc+J7O+Pyv+W20IbjDy
WPj7sz197i5NrQMP7kaHka42BGjM/gHH9YDgz3sp0ASQ8xxlKBflYeH8I/eC/TL2KdD1/khQcKUt
LrKGBryxr7lPjsYZmfhK1bjuv+7EExcXr2NQFvfxpK9I09x4XTYKtJ2UCm/GzKBjeDn3gHOrGiqs
kG4ainvvo7cUk4mwoyn1eMLLV6RvBBv1fvHfmut/xD+a2AOef2oq1+LK4cpaTr44Jxc47A6aSVUX
Lpy1yvMVdf802z8AoFv+1iAw9yvSjk3uj267/3J28Lm+bufHiwqrIgjZvtHm/OvWPi8g58JzBcCl
ezmGtomsRRVMPfFhq9r5qYwj0oWHNLwx6XrX6n+3sn5C/qVpZKk1Xsq8WZpnbeedW+rYn/7+0gmm
Ygnv2bN/3HqcbGvSqM9osZB6B5jUY4TQAnKxqMy9cUw7gQIsIjH1biT5UeDa53BxdORd8hV6rWuL
3g7xi3FkRjkOB1pn+l3Cmzy0UtieIXaqAoL2Rg355b1ecWv2KRhD3Qd0lguPkjXlWIvnxEGzItPI
MU26ntF/XNI0uYrJi/yAvQ4vmadHD5skHT3GWsSPCNP5vfKyk8vQeLbB/Q+/KFzs2HwB+EZCekpY
fMTykA6DTaJyJkvVVbwAqaJQPls89IzCpXnQjiV8BYkhpwxSaGn5DJIdvABkN1iSobXp3byyHLwh
XyOSAQlzYXjw7oJf/hhHi6SA+dQH+hz4B7IHxz+7JEbFUT5N30LbPiEvCcTmVwVFCOAi1pXwRH49
2prLdv0h21uZqyXSu3oMjDz+GnV5S9lAa1B9XEdcxdd1O/Tq6rxrWu3lXTp0qjufi7Hn+K6yDNqa
+QFIrkQ9UDycDHoMOE3qZv/gerzVjr0+SoXU06f2CcAutkO3gEl4RNvWu1ZJqJDUmRDvZyZBud4k
6I/C7Wi+YwbJR1/oHFT3YG3xBZejzc2icfRlRRL9r/eQMeoVdkn0nHE7X8FwzrEUKOmaLEmjOJId
4vDzmLMInw79irl+9gfsNWUX0Wvo1xMm0+OZwetJD30NjaJg8thXcj69jJ+rYhp+SgdYINnFtQrX
WMpkHYf89klHrJoH2qME669YockCsBNIAgP6wevoxIn4LR0i5hWFmDB8t8gfvZD4fPXldz1gyZnh
sRtdMeNjeuIFYo1226QKivm8U4ONlUJU7i/9u8zoXy5pSS8D4YYRHyF4Mb464W/craTlrcTxWmA5
eicJHZZWoeWZaMAIkTm8wyZ0KDMDT72plxbQ+ef7ayXOudYuXFQpCFX5KxKSDwJX2P8sNgd7pDAn
vmzTngjndaxSbfCJCkzAgIq/21yC9x8ps+uRUoIpQ0yDQtYboclklRm0kyLeX726GSBeyd6EXa0h
+q4ccm6DlcC1RSjLbftGcpjMJdCqH+EKy/6tBdcy+EGOCK45TyZyF1v8RaFG18hNiwwaF4yG2vYV
ala0CA7y2dk3xNDu4LZIzvuQqYT4XKg+ygiOAJEdvwYlDbC1fQcxTMH7TD6SUU7qVIaMAXJm2IUy
1a91jsJugUwn7fH/GP/937l0n5oyXGZNpnJogTouHHgtY1LLHjv8/YbL5SKowm43C0YJT1bTGzk2
1LJaqRhsWWdKCsaRPMrSI6Fx7Lg+klO5go0/mN3auTTwt//Yvt/S041IMzyMV/+t7vM5HsLbzYAG
DfCgb8wL6oCRUa5OGE/r15Tr4FRrOAHws1VN8IH+37qz9vkKUwSrKiciO6/3869+hYcy3eieS36+
X/KyEvZ0z5G3mD85xKuJOm0h4yUSm3UfeUc3+y4Ys5NknA6RkpZj3A9kf6gdzyTyjrtfQlHvMnC9
weLDlZdxnUH7VoLZGgb8UJ/OX7BcafDY2OVNxq0e6r7mAzFpBWvIN+KD5BswLX7mgOu2yV4OnHBD
NLj6Qf4UttJEbfyODJzVPeuIE83kFFnhT9ZuFCurXDpx9L6d7lf0ayG1xzeSRhEQeFcrmEt2BNTB
YYUHBO+zCkXC6gtHcR5S0mRQzghm7Cgy+C1evXEjF8zp59gMXBQOUeXzj2WdoXAtJcguV9i+xMu3
/t4TIWvdOGwPO2iRzbSEPtObqRLurwqbro9nBW8FwXlZ5CqO788zOkWPP9qh8wir3E3u3cRDSyFu
ZYrdf4jMfjxKSX2Y3qoHKUhrjZ0nZmGprzzYGIwZI5pn4YWKnzRB3HCIzyjRoxVH5DTx0X4nS6ly
tDuIIsrHg/K2cXoSBr5u0ypRdKnzVkQcE+0P3C7tTsA6RRn3q/+T/sSQEhbv+44m0R7HeICdk50R
6qGN00xGTHmFHL/37gRVpITA08flzWUuCJOqv+LIGDUuVai/vydBW4uwdGmVEv1H3wkzmEj6opgt
c9uW54/GG70mMIZLZt/WdmREInzA3VSD7M4yh/wrWOuu4f9hf8K9/5lmcjP4YRe3UkmJDPtAz+S7
WA3/CqVgyJTtJnnH7PgVux/ppwTP+5fmbEv/uOV0+MjPzKt+2xPr+uufnVmdKf7HKZCeeAReCX07
50MGjrqrbh43eGFSUuLfIVjf/Rsadt2WyFcVaBEHWnvOunWsjZJBKSHt8WJ14JTZ0glI0SMltsK/
s2qfGPdmJ13oLci0MIJKxPK5xyabrQmT+DK70D9uYvpOfXTUdf40peDpJi6CaEbFo3LuOrtW/5Y1
kuY8+FTaOJFazSm94pBmaiZnAEfgyeRa5mlDty8PPxvqwyTCCVrWLgxu9qjQnN1sXHauhzL8Nepp
ErWgjbOFTfYAuhLe9sT/WM1ci+kl5EslC0sGYCMATfTOClqyvrQ7By95M3CJtuVHg24UkcFHiYcY
E69EE+SFksZwVB+TCzPkJFNxc/OYxMWamDHc9GRxFNbuT72Bw9PcKQW+aQ8AK3K+hME64yk/FCKW
VrZcC0WgkTnwue8tLK02NOo9C1NdvC3Hi+1IaWKvl6jigGXRqxI/wq2hyGFeMAAWGw35N137SLJo
CpalnMo+eF5NsrnRqzfdPPV9+01mZBN3x291CNu312jM4XhhI0akyigr0GtA4wSdpUP9ys4Xm10D
SCEXFs+QDcfw3dpelmE3+PD7CeuS3zSzCXx4lC3OuFV7hh0CXnsCdkELJ2kiUpwebcEo082e6qVa
WeyFSE754aFDjgoYgAywd5ZWOYE/OFoKRjfV78z5ILz9wUce9/7ZZPIUXbllO4uHbmESKmd+/BXT
zFjZ1h/5EbLoNxw5y+mCBAkXkEpI0P4EedDWajpxtqZthDe0xRj5Ga0I1pUp0AXAgoiT3LHmun2s
9xx6yRcSC8km0FE3pSG2CxDpCef0n9Uj5c5dlzQfGZHBUQ5eZ4qU/BvGcwwaO5OXZvCmlnNOR2O4
R595OXVf2L7pBxHXH5eFBiC+ea5RbPUdEO1d8C4uTJ5HzILcieIJkKmt6S9Q6eDjlx/xPv/DVSbJ
WI2eQufhsMbq1esCLR1z2lpU0JNBftCi9938oMuCaeg7/A7/I6dK7AorxE70GafLut9A8sNk1MHf
LUwUOraVAs3BdLWES0mbQnfznqFxUUMKZj7zFN1yrBHY2y7Wb1MMG33HaALB82l3D8TJAkYosQJn
KMhSFiu/lJVenVBgXq/0mwBCLD+YyXPqMiqGyV6wPUbOkrso+27KanhIPzoAYbigdxRr8Cgct4uI
vIVPEfaGFYsPdLP1BOR9dLyonH7h7vY1EyLJL5Yjj0q6Y/NTuKrkWu82OuphMjJrJie6e09ovN91
aYLBe++F4IpBGGNT0clba9ip7E1BrpILKuYhbKqMkkgf2pubW7tGmgb8DJp1Z2mK+ZindII5boOW
L3s9xcUJIKKNGIy9VkeKg2gfGfNTMbC7I746E86CRzyOrL1R/KbenfzafEmcsonA1ORgtAOxRlH6
YhaIL+N7fLEVboeRP3fHMkPJaBqLm2gu/2HcUmr47J5oaC8BlV8DVARFwUMntJXY+dHmxYsxZjtE
KTQxPoIIIbE/ZjQEwa6FQzvm8WnIjdQR/kZrEP20HsfXAflECnzzH9pR2762vMK7sIUmf9IdVDQr
1a8JD6MMYFwZWSqFRgRL1CJsB5rLznQl5EvDZCCSGB7xpXyxUwW3c6fOjVoiUPEm4fEA8g8B8AS/
waLwiTXhcIbPofHjK53afqfDWDJqTj6T7rbWrh0g2hT7SmMB4KqQkrkFf3AiyCM1RbqpIDI2oXQT
ztNrDGRDwYY46tzhVrGO9Av3y/ULI0qP09iImT2iejFUT5SscK9hHjOmQkEemSn0YDdYWPLJNilD
RA1tnPgyqAA/ivkwmTZAuwZnWeOGTq5U4hNyALc78pLa0898bbxj1j2bJEXLvxSkNQMbLvjsGKC6
hHRExovYPyN4a8KCKfZxMNFEUzZbTPij/+e7lx3HrFlD2PcoYGGwCWDE3vLjm65ikJ49Defe22xg
Yb+80fJHnfN/O3cr8pUovoqfdeerAI3xCCQaRadMnwuMrHGpQTfHP7Dclg1jZlZCoOtH6vFDLK6g
wT1y2X/h4bcWi4cNytDj+Gsu5S+OYi+PSh3XBeuJwcpPtRA0sWeXdClFJzSRjQITodfpwZ9ccAjs
Pflk1XXyBg6JwaVmzkPoJW0PqrVyjQOtQcdiDpYO+R5tSKHigcuBRt9MIT4YQD3vmhwcF0RT3g1Y
o84ZsPVMrunIvQm+FscDewv0swvAWcZNWns+XhT8kIfRdU8vtF6S8SkdRs3ti9jHnMqv44PO2exG
4NjVlCBAyCOrTxWtYnjMfezABqhRYAcSSNqNns1r9/urXrvfmplMaOyA4Y76pVkCpbQO3za7Txg8
yN/fKrIidWLXwt38/WIOO4qCF2HUF1fkVYoSb/fxJBJemkPkEF4TDBzfLinWrqEr7ah3Rgf6UiB5
ZjjYrN0K3mZDK2haB7hpE2Qsesl0VYRSkPt50Co2LSLD5c4A+Pqwga2544qZaTfG+zhG+aui3Ozg
62k12SW8mjz7PISzzwTEHY4Y+wWyGOzugX4nXmM9G1M7K217H5qVS9ecUGrOMuJ0y0hWLwoujATg
bhv6wjXPF7eXkfD5d6zZeE6zUnNnpWtqM4JXLxQsB53fA8+oqHN+iostuO/0/cWXLWiCxrYm4bp+
NxMS4KLM6GFHzAgwckVBP/rBIAs1REOuTEne5CXEKSbosmhnVX9xRutHNnsttiAqOSIVuqwWSjMv
3TkUmP8RefAddp4MOeRWZ/qGx/W2QFOT7qTrHcWHRs2MVG2/hmrmABFijolu2jYKaBBK+t13bVDy
+rEEnFc3wyOzNT9Vt44Aw810/Xm0pHnZJKmkTcGhylbn09A9/cFLrK1IHbP6p17hY5s4DJXihL/q
ePfPsk9j0dnQOZd1m+z63OGgIJFAIGVHTHLilQTIHh8pCIj91qGElWTmuDOxGqRPf1l0j8CoVFtN
nkoxPdkMAH7nb/Xx7i+W7QLP5laumE2GXahplNzV5rECUc+YdS1XFkrOCdTH0plSuWosIiTsgSDR
FgbZTz1IwGR3PEs5uycUswVWX05mUvq2uw0o5lSH6+pcEty5sFppHBqFuaq/HXYGWe2bgTLBmDMk
ZknHnU8qyCqCYCaVVlU0v4nqwWPY2RQQRhzNI9PpnT8LrR9QSzDvfbKycxQoFm+RKQJ0vmrZMJHn
bV84Nj8pFmF5x8Pv5UrryW2VOJgvVPjHVhi3Wtb5ut/0KhFtaqiYA0dQv3V9XvTswyetj4yah+L2
gMVnwtlmHFqDZI/PCf1ZnypomDKlqD6PkMzjSTV5c82WuZRozLlLzz3vx0aif1qI6WLHzloEXWaC
yyYdAZpet+1iAMU4d0DQfyZzQ5blwyJNfm54uHGyXIqESJSM7zh6BUXNDqP/jDSkD0MHJHz4c494
SEuJ6te8SweCT/ZORv92/sq7yItZtTMU52PCJNvce4Z3j4EBGD/fUKrQrocu/opsxPJxsgLNDLH7
mgRezTJJlHvwEsHzStGemyzNXIMOYDllVsQ8n3N12dGctLDIaFeqPNAhNFb68jgkixMRnKOgx99c
oMcKrNgFlAwA4NjgyTVApA2j+5cyeUYRS9suCafO8OqRKAYw3Cv7SaK2E/AYDGpqHqmE/08c5pIY
utirHvMzcKZHc8YRP+x3tyarw5twKwYJzp428tjbUQloStI++Lj9B2lCIa9xpDmEEodDIpMZ/WFy
utNkd3RIqU105CtK+9rVMIXRy8vLVs16X3LM+SjRVzwVlDB2Jt1O/bKsMa55sahpHNhlmK4Ol+22
RAwEPgFsZiPddckxSi2EHxT7FQPgx2xUfNzgNiieKwTEGvr9nIajLR8SrjRF2iyKwjQeiqVMptJg
MOPGmwDeoBCkn/vaIMb9d/OdmaZ90qSLTZzc+gvMgyhKqdSOd3YZ80QWW0pkDXLysT701WUTEuJR
1aD4UFUlexUvA4xvWanysCbP3tmiTFW8VGZi5kL3uRn3kaaQciwNeD0kDjbL7OhNzjhTUsfcOQjM
NRRbVxJOL6QYekBJcgLFOt/Qm2MQB1pjEJoRDDVZq4xmzq75aGfL5Z2pAL+2ijiNd0Xdy/PQq0yi
vxxrQrYw8TqtEZ1hoICyV5psSkqU1AKCrSYIdryqqISjwm9SGZ6lYTAzVHv+XgOtuaLX7Y7A+PrO
hvGQEHgarf42xQhQrx2r+BJoWhy/jQPfgyzk9FxX1m76BhHwV9ZsTOKKAC78cMhioi03abtELpmz
S0RbGIk4oHyw01DS6t83SMqXi5FQXAUf9BZsVU8UDacfscwJF2PuZ3ZLzMiEMFLF0LIJulpCdvT4
Q7BGW2CuJNvs5vKLA4rtqV6Wz7qnTmZaFHoYgPdbbC3OjFMOHE/Na/gHXEjg8Raiar5FgjALxfTK
M6zhvNU40ZSo1X00kyTMvEeP/qAVOeToniUDfFcIkWlAd7DYh/5vN9EfEUK9d25KrMBigT/QNwxM
MPxrsXIf3If5jFyOZcxIQ0Wx4omw4bzwLQJZXiECXXEGGJckUEZyLAZ0XN9T7s6+frj3xmemu6oC
vAwwJM+1Z+zb27cOcDZjljj8NWTDZB45IjqAAOK8Jiz20xPBqadS4gagqbJkeuz8Q4Bec1SN7ma9
T2ZXxbaInTnEX0G7rT08pBu6jIeZoazuXtQoS4uIZ4PCZzh6uuow/Wc6+e5ZkSAW1xXBcs6m+JC2
cXu/T28uRFTYcKVvqqlxrLI1APgLcevFx2uv5WTmOWcrfba9NvzgXGLJN9axmtDWdSnxbLOSWM7n
T2V2qH2SL6B19CsIgIox0Ygw/W7AVKt+2mO2EuZ3JutRyih2QnP5bg38VqLZ/TIHQJoeXu9pXRg9
DWpWjLldipVKJY+toSv1Y0E3oSSeLHtVesJFGUWjSBaXWyQ25+JHcErnPLC4ujPYDM/sRfRODmTy
dfvVKMVjccee6+2/nzbBgC8Hbjr+l+Hq375cKKsPr/pwrU9Mjq449Hl7VTQI3Tq0XoW+Lmp6aD6d
YdQtnMEg56S4PnkBvKx1ZQmZC0tc8eByTQkxB/F1Kj+AfDV/LT0L4GQiaEVLpQ7AX1UJ4mD6gF7y
ua+2QdnQ28bKnfvyF+GJAwsMG426Ex/S4x0nVLpv54vR36kvauBSWkwsHF+9xiBWtc8nYNXv0hq0
BanUcc9LRwHwKnxmUxWUkaEkTBOd+/EYrFzhKZl+48Hf9w0VQlKhI8LBpXGxra+YWziDZX8fKJ0u
wAIQpxKURQmJlUM8dS29nNbgNZ+DecDs/L08VHA3d+T2OS19/o1BVVKUMvkvAS8+4+c6QHeu8RB+
xoy1duPtC/pX3psXIi5jixa1SKnbiEXQcHtpuYQN0m0HqBp6nTOHNbEFaPkVnhrw+D7BYe8qv558
9E2xvVd3tlkcuZAd1qBmauY56Nf/eJycQUhCdL0lzmS6+4tYt+Th1Uvcvd5sr/qj4aRYXDsNIGru
xpedltHekl1ma42Iz8PfcukaRpBYCprck+CpjQ8j7qP9vA6hn1tY8N+Ei/AJkkGY817PA+jP7pzW
4Hlt1/X72+9Av5MpseZynldCamuCZTBwnBWNJZXsP0Q/BnP+xHzYzhkAdA9hgSreTWubM3z/OCdh
V4LggEdV1hwY5N/qqXhBj7lXhDjbo+QSfY7Sv4lax89C7gRY68QA6BdfBLlnivIqCN4f9PFezJTN
wdcWa9ephuv7C0o6cx9hwhk6BUdmLxQ3I75A6acZpAAlx72Ob4ITYHAcNClsYu0nwHElhoCZ2/ZP
2U5gZZyUAi/Kvp6hjN6MqVVAmL3lctRmclLsBo5TbuThZQw27jaBU0t73jvnKJstpYdNxaIliCJF
YAlbAxvj0bNgqDYwlt2x92wqk98hkwd4ZW00vA1zE6Iiq71gNBeJFWhjtYdUgcL7vdwyl7/VYfcG
0HTk+FREbhK84s14cjKgIcKGPratJWPpnUX4zsX3n2FzHP9vIcM4UxelHastBSfRk4+9y5QIihG7
ZvFc3RPfFomjIRlupmlX1/joBswYgtktD5RCMhwrNypPYQKtwapXwcOnZzygbCAg85vE0yOWFQsp
IYd813c3+9ti7f9ig3gU9lcZsFU4lh+OGaex1t8n4+/VjcVYLmeSokeAXKUoe8d4Ve4FSXiMriwF
WrsFZTbaHGaJsWCTUqkMDC1akpizFeHNzIxyGZmEKLCWHG9iInPDAA7yPE1WXmBmcoJ3GhrtSE5C
rgrd+AGO7qt4qBYin3DjOFlaZrbNsFB53lMiddWmkwXQsF15N+UnJ2DFuqpEbYhtFkKeNcqus86b
eDzEZG3rpVhBcBT/Y9yuv2hZCyscgKqm8tv8TIqhQjhVnTqXSYiNacmxxMhigoDelW7q9Y3lYTiP
KoHUp3sYvdZsGOk0pWBcCG/97qbFXYPth3w9F+61a24rPBPFN69WcCdzt4MjSuyIgRnUF9yOKCV/
LfHph2ZATazg+Aw8hq8x5gg6rv2ElvmBFW2hJ0jElB2AvGHT1AdGMGKPYD75Evu8vkvhqB7x5m9Q
NWUtm9AUq8H5l9MHPLNLaLmzKXVB9zGamZOV5mOP4KSQRgsYhVXwzFEuRoAsvtXYSjQrkH++1h43
MGpgbQ3BR7yRJlMFVOnUSrLVJxNCHFu517ArT3MRX3jHYHrH14tqD6Ym7kfbVf7/80O3+o4jJVvs
ESIKSePno4FOdShRQuTfF9mNy2S4S2e5of6m7ySNNcLs7upE1Jwp0wNcWnWdVsIUjeWutIBvtLXT
fUK8DWH7NVoAnIsf7Eye0K0vRwqUCLS5LUhe4mQ03BsmeXR/fHN0WcNxWgetXVm8rWzMLmKV8tkl
tfrCsD/LVekO0gsXLB4I9v8hFQ18S2wmqeiueupv5htTm5zPh5rW2GoKmZjDR+o2Nfn0IA0ghFis
zDYwYeqi8tu9miAM6M+Xf0SocDPD6oWfNHWBo22dRZiFpkHjCSuwcSb+02D3mVqMeerFbrbWbWEY
Rox1ZYhb25Zl+Gt7wDQY0HgbO0x9dk6PAONduHbnrz3auFdNfK9xwr4EWBxmRWDQ4w0UhD3k8jCM
NDx29txmqjLWZfhYO0mAg1D/jT8t2xpu7DTNLoCfKnLSeSmEQCs8D0EQNhIZjvXiuWJX0NP6W+q6
aGfbH6ghJKny5TAzeK6vh4SBrofqn++5Q5PGO3IhcT7iqJIQDA0kgfa/Rn3PAm2CFuEImlltKc+j
3C0eHSt61AhELvQNXS4RqyfrHNzOEIoKOi9LB5+kyPKbIbosIje67iWNrQ/XxqHlcScFfKeHKqwL
8Ffq/Bvn+Uh18mPO3ptXwmCEJP+fRAaWBgLq3YODtvfyYuQHSah1xrKup8VKNqjEMmXn1zvj1HZj
z6bgRJhg8wj4juBvcGFoEnIx+reoZz2SIO7LMapmuqINThL2oM5a18NH6VuytoOrWtEQ4CKxbvFV
TZAgYb+whO3LrRAComrF4OjGU8vhy2+/jhCEbdsELKbGKAXpDrmhnsCcTxqyekYrsV4s3xap8NbU
ZK0CE4QdJu2RzZ16AcG6EFc6YLQ6RI1Vr2o37/sZZlA5MJfmKJiQInEAZ6R/oVRqVdLM0UtnOxUQ
8TR9Yj3lrIktmByeHhyEmKbx1gVSnIYcRYWJ1zMEV1V+t2bVhmHhIwb5Iof7tU7eOrn4d+f/pQVN
9JBLCmzoEeM8WRMK+rs6vIDLZ/wm1wlpy6AvkQigUSjA2/1Z9MaPj/V3LY6YsUsD7hujPXcq7vNv
qZS4+0CbYsw1+9XphMbUCKnMPiVjs2dp9DbiXD+e9jwPvNK5I2G2M3mwF2iEa0KmIppNBwsZu4ES
TsCEvpQLDhSLq9rzRzI6sYoPWgXZQVKGvDRZhSadGqruaxubfon/SwKo878u/LnP8Tazhyb6nTdc
xcastXsP7h9qB+g5FIIy4hY4JEpJTT6/gS0K4GmlnQygl15Nyg2wWWEFy80OE0SBwXtCz7vwkpi7
MvWDjkTtUUJPUnkEmYEvPAiL8e0waudOXa2db1V79MbIDAv87VVFT38oyllOEZqHfiaX4Q/r57nT
7/jZlpN7U2w+7WMel20jV2xpcJUqd9Hs9+a6inXnK9DIbY16KwPax1sgaSsVq0RNBwMnzeyxSkzy
eGSzneX9cskE+mftKpWh+PiMUAOtjG2DIKGaWA/clwVhkuV4+aSpid5Pc9divNTEJTJCHOd9wW7A
5B1aVfMBefd4ZLKDN8AphPuMNH1ATyi/gqkmz7E42bVmfQ9D5bGjK+Upj4eDs4911Sg/MJZBICdv
d1Bsod/5LFZJn3pgdp6bzUpm/msbbgrwnDuJPHiVITBNC9IJ7uU5XjeYSKB2m3/biL4vrS/m/eCs
/b06zHzxlzfE0LkACcQk4XrsJ5TQYfZv87DED9olW8ohwBA25beHn1NBGaGgTIDZfM3PkzP3ECmk
LIKOJJ10OY2e8tDgipiWIfhtW2flFziwhyeYTg7AY6pVz7oME7+3u1Bjm5Es7yrRWm19SGxzYQsY
lbmjN21mIsk37pIMwad2Ast7HQmZqeJMmTABk1kiMMO6gAcQ+0UmSmkGzkN6HMtOY6unl/IqeJzm
C8PbXyqZppLm5YAJx2xX9jj7Hq+2MK311JwlJebp9FOFcarE7uqrXrGkLv6QrCdWHKJLjTWvJue7
o08dyNW65picCA4HRD3KNFwLE+ZJApXD22/pMoYbZkiytLC9CcTu76EyVHOMUF5ldvEHQyPS00rD
6m+wu2exyaPAay8es+JIdAnHhcUqY5dILdvOJ9LNzCW1nahFPwx4d43QB+sn+XQqvnkwrOlG8okg
PPRBYDXiuu6epo3EZ0BIqdjrIehqMtaZ2vZ9PIQcutj/b19cxOPgULophvUn2Td9yWIKq3tPxx+K
1RPSAqLb8zRt12AI4P+2JZR2XegSDsHF/BCO3P4Ov0jlMNkMsB2yp35NHD4jo76/63KJ5z82oRcX
19sxLLnji5PUExUcPizc7X6M974abSzEnwwAIz8HwnokhREU54RyMWTfVsjGj1PaOxyP/5SNnhCQ
SyJ8m5wr+FatoovDqbItLNPEJ1jAaz7mvAeMPYFvZSZgwjy90WBUbzNIoyDFzGGDgytA7qNYN09C
wrCY/T9P1mwLMxNNWWRHk+MMpCdirnYPROr3H9z5QVvxhUKishSsQ+VZqEFSRCkGsD551EqXxeKC
JndYu3jtGQQb/k6L3vDIEpm30gUL1xgrFkK6QdomrCqlW1PrWby0AKphkHThfctY5JssVQsHnrGk
IY4/wzqpllejJZCMpO/qTTbM5MJHGVmaz6+hlLqlgwRT65vTZm2aIKVhmIkmTgBsvjDLlDdiBVZb
QRSFLdT4iTBQIogo4bk6aDcosBx4oKGNuTeqqbkWcso3GpCGSCVMcDF4jBvewDaquObYImpEo2pQ
zjYlFNcfMNX4CbpzxmshOc4t8f7Hjbg2sM4CClvYTJ99RNKEHbt4jYdqdZz2MmHLN3JH988EvEzd
EsmTDjNrb0cKF7OdGs4YWq7nJISQLRCaY10R8DzMYUFt7KS/7okCHM7P5tSI0sLIyX2zt64EDYnm
dHoOWYPP8XHOPF+KBxfmrMDR/ZQhYYvkr3SPwca0c9xqhqTncyhUD/I+TUljWSZjUUOBdCFvNKHt
jSAEftqy0h9bGA902CrzGk4IrmpnQNTem8h0MoZH/SY4R6TXDuz/6oozqO5cwZc6/7zRzBKELqa/
gVz8mZsffzMxS3YAGMyn/YveOovDve38TeLgn4AnHArVyHNFdA8jKS5S3mkEGynfdAGEeijN+CkN
LQjY7zQ8+zbPyMrYFLbxsJ3PXapIC8BTrkG+XL7FoAY1Tqn10n991m9XjCoxOLVNDavuxO8w/V6Z
DqbDhF1sKkmhgAiszSuxSD8UQ+xoH6QdQg3uf4/IWlBMjXutxlqIjmiYVNLcdA3BkzXBWXpImg8X
A7571dB1d4p8qnjM/427W5h+WVygKUPSG11Uexo331OT/m7X4mmR+01N2JX0w3vkEzpHW8xgVlOZ
njbrjMRUNhv3aMsjvFcvuoBCAeBb3HGpdfuIDv7PO+28n4QOq/5Zc/4twjOpXg8hc8zF+Fyp/uOW
PAQ4kjDarMCz/ZIwDLfbpjuRY+1pDov4889zquZ3mjKdg4p6NSRvWbRn74x4y/8fJwvqzeEPCU5L
edxURP330KigzJJM5hyEQxeZLWioKk6wECstjBcbfZnWh9Sjp1g4WuHiBSaWcgPJ5BMjKoDZeddj
1mXLgKE5LF+5eEaYGl5LfySHAVaSUNolDAvvZ53GWxlBmdxbo+/CI05rgy6y5ItKxE+Nb0EEgfT8
8X6/0WFi+wARXBwZADkmn89BtkFPgDyK0CyVggpJZDFrl9sULVCkjbq/6/elDb87TmECai/eShKY
WXcUJHinIZJkp5BAmvsyFwOtqakR9qMQ6yc7uEO93qCOGiP6u7ZbfUEu645wpHGuLMdbbToM4l47
yNTgM91GwhbTmyt1WTs2dKg0eH/m2jsQQP7NbWBwba3yGmrsaKpNxQl710N00yJRQJKhEvSrQPL4
sy/tdoEi9YdgFVgSrmfaLFXSfgqmX8JolC9gaAXMhvFirWcDPFHK+ksU+eaXzKcBw5hCn5UWppfb
bp8rmccGBjz2ZIAtiIvciHvEBaNOHI9mINVwtxlBnUh6jdTgRBwlvPtV3onDrZA3uX6dDEePIoHF
+sON9NxXmy6yDgtes3Rep4ZRIgTrZpZiPT0tPXw/WGnzqbx2so64k0Vxy0gMsJcR6l685np+41b4
3I35Q3Mi7bzs1iaiuuw+GdytYDhGXqSlcjP0kbyWcbnoyAVPUwU8dRo/CKAxoxwGZx+XFEEs/RVP
PHerBCL8VYUVt3DCpQ4dBw7cmTTtPNtOJoaY4ynAw435wO9fsAC9ghrBqadIx4LzudeOszr71spg
lcbGv70jh7QxhYFgXvF/0e3yNsOI6oWhIhkIg3sjI2mLj2qBRsURYqC4vSabwkMhL2KrrLeMuMR/
XRUb+VKmON0aT3q/I1gZ1pfk/eisEmeU2PxV8+bOR+PE2ZGekJBb3hv9+ehloq2TCxuHps1Xg+ZP
EYuoUwBBowdNVR+HFX48IAgrvu5saJXaCn8EuvbG1gqJYkH8o/6dtyfFBJVe3fr8VmXKtUinr9DK
WhRRMqTMWkPAywDRA71vePFE+1wiO2zHsTSWcHFCZWkH5py14SrVBg3iTFDP6JiWtmA+cmJPDVpW
J50Y9YZLagcz5ZVqLzVqd47OKHiw8qciWnB4ZCtfHZouLr6lBMspr30zuu3s0u+/UkFE7NuWaeQP
t79pLG3pHwcPhisQpizUu9NI1cDm4CRYD/YBx80iN5WExK0BkQ1NF1QQUKspOd3O9zyNbbQyDTvL
bm6NbYOX4VhgtOZZ3YBkQBNkGx9ht+DKUJMz+xdC3u1v+XcgfRTSXeMdX5Gdwh357s6vbyILuFss
HAUJUYV8H9xX5aVvb4kBlR6obW4nE3oANrSnFq0Sy4j4iYTi/DAkDIW2flhT8/CJLMsCuYzuORhM
+V2ml4hzQx2vl12QQtE445sqUA3nPI48cK06LEPir9KuMeSgeez6VtskUeyZMFsmuzrJOoS+gf8y
K9sqmKjOdUr1V/RMtHTvqQ6c/4JwugPykn6UwjfAcXrJvx4l9mfeEjTHUi5i3cADhwl989bgHWbT
KQ75JHV3Sn/QG6ZAAuQAFrx7QFxd6wwsgSix5jj5ITg3kyDPktIqzlDGak4THJycAtPZNLdbJk6w
JOQrjn53qgcTrNiiqVKWwmZglcsdk7wwCYVHurA5GsXuIruGor/Yar9l1cowN+V/8ZM7pdLt+qtc
ave6o3WIPUZ9DYYm5UwaOx9vdDvOyd5JiSg27cj87vuVZNgjd5nMuXf2ww65xYuIYDsZYrGG1+7X
r66++5ekvgH1hlEdjzrf8lmqkWfW3usZL1YqZW60gaAf0Tc/w1rlAXgxNjU4BYPMM1PwXKKYCiIP
I2tPHvLccaWDUBmiemtR7aoAG+FEJp39XQGmpLIO95ZyU4sKYY1adbmmFoZRDquXddWDrXZqKYzM
ukbi2oY30LZWqswI0kQdPqF7eWCEvKExblV02vvI1UFPv7Qs/gGQLvM1d2IQQJXg46UvLb6Y1tzk
cfPePKNfL9jDJ4Lbwiq9ysAKc/yL25QpgUnOE/ZQRurzLZyI2E43GkVvh0ZPP0JCiYG78P5txjFi
tNnxdO05u6KVQsQjwO/ldUCVXunJJ9ZKf1HoZdfmajQg+IBGlguiUyONFBnfiOFz++0kBi5Wvibu
qepWZu6I7LmjkTn4bA+M9CqPjcbO1tcTNCTdJTv9ioXqS/iI8YveOCFtsyYP7xf9U+EnopywIltt
6b41LRwaen0HbU7nAdU5c9sfHF5HeOLxYLHm27afBlijJuYeRWjlk5u/1vwyM0Oe98qOnUwdBxic
l1+Vng3cYzqRvjTAKkK+pUt5bQ94L4xAKjq4f+s8yea5tthcLcKY8mowOs7SVcchhbzn6kTDepGV
qzXDIAORmCrHZGmvuch0zq/e+N7Ptlkg6QIPOgFprRZIMp3FP/1KxpzXbe6Dyw9rlPLLLClgoLyK
awOUB8bjTxn6V3MYG0p0Cp4+EyEkvpzneP1+/xqytSFGHn0SxpcCyUsmujBCrY4AvVsvLoQW2MiZ
eXhqP7sX5iHXkLU7ychR8CGTPoGKGWbChbXiF6jbp9Yi3hQNbD6LECB8NF+kmgcyydbqY5c50baj
e7uGve683tfe7JabCWetBXPmOrcLPsTXA4txOiBBdMamUGLcmQ1kSe5qJJ76IbKpZF+WMuwoptMk
txg+VBwgbSPFxbKxq/q5fyqoAihwJuBLqqkNwIiXtwXTiszOEFvMaoUMGCHCudu7eb7Epi9ztKIA
c6t80vzJMi5dxNCTDTdyNl36J6u6FubR6MOuiRNar37K6tJ24dFAJKn/zVaa9TiBsVWhbiccaU63
OYY8wHrTm3x2l0OM/4z59AZyXkbNE/sUQwfBFWv4a8eHtYYDhXd7e4IPg5pXUPKFw4644+qDOdgu
kJ42Sbiw0NYIeWEy2Ppa/m7PtSGgn6J2ywK6cXb7SU87aRrl38/8ygB+dYKqJtzz+ff6lc4hKXf8
uRHKcu5QEfJNEQyP4LfinMfMXMKUzCPje6ht7VsCwdqgrNTbioepYPJHlIwLPp4HeSg0a/N1q72M
yp89dryEb+Uigam7ucQrl/xCqXssQ6BL1JgbxR3CzI799SPxEPHHq50O6Vq8dgzFUD1IlhrbqkHH
fB+LZq/8gUPJmaIyNXWRWUns3HQqZ2noaJSaZLi1fNLG/1VXIQz7h6FYcGX5qxjZROySuUtGy5k9
dlmBCknx5uUVkt1pfLxMTU7UuBBnoFoBtg5reXBnM55MTMmhyqC6PH7ejup+sn+LyB2Ykqz5tViF
jQp6V8l9IvK+nqCHYUjUAam1PKuUBEapVPLw1Tzbfm49Wn0zNCXWeTrCCXK/N8sMLaVXgVVmppTi
Y76RnblBrYHSEKl/WIgIWLji6qlw1Zf7a+059pTJA/4d8EROVoto7BvwsJv7vG1o1UOCjALwQHyi
JaTz4SG5UC+sTlDD58thioqJu4c09C+U7H0fYPm6SarA2HAILUtoKQj1CJ23rmPcobhJRCD59z3P
juKrCV226R7mBcfYJe4hUTqqnWDsQ8L0AIpsLJw5pN+CMDW2hulygFBV2MXiGSpPSZYgcRXMSoky
73ECbvaaaMmuj9/sCAho5EWk/fhiTj7UbGTSk60BHHMCjwKW6j5nw6rRPf/7TNhDKljC1bFL1UDU
mrZAkJtHhXc3WVnRhRBkwuZDRoOwGzCKG9iLsY+ZG6tOakA9WxaE13V9PI+dHvWa86N0U3YyPhOB
LnvM2dbwNWhRrj8Degrj0MAHUkyjy6eHkk0cxC2LnhuVM3IwAQenzYWC880oMgKYaZelwoL6zN3t
rN7Ec6BspN106/a2HBC5qW0/1PBn7hKCtkPM56pCx1/u3D6SuU99et11zj9riWx3ju/iJe4RFeeL
WBBpJ3kTsNpUZJX+yrv6OeoVXdVwokc11sfRy3W9TrQUSuRF3yrq41TCkXLey46WaRjxJxJhJZj2
Z+oR6O5Cc4YfqbBGulAGDOFlXqlQse4Q4dTOTe/MTI/rOFZMRuTJShgrpsarc+KL/QEmn78r+XvO
UpuaYtDLDhOVgdFhlPmd/GZEkp2Vx6Gq9DJY4XatD9RlN3bwUVOtY4X09P69Od/oGM9G9Y5NDqOJ
Ps+WySoJggQkPE5elKFBEsTIFMvlTo2yHSO37HblYvb66XabpEMHi3OrZtuYk3d+GXmxHBPA4qo2
9BT9Grj7hJElhwVZ967ulDdpC3ylzF71ZOPow0M4QO0xf+9bXcgm9u7ywBPdAm1ee+l4GGv74RqL
3OBKthur16bvM9f7hWAnTp5pzYaN8nxArCNf0JDiFjtYa+4ivRgUv88h6FsRElTClPK1c4NiE5ep
MiB9zVGw+9s1X8HHm8eaVcetBrcyqSE4b9vOuUkP7Hbzb3H8hV795f3I6gmJebBYgJqP05kIRA/x
jd4uoW3jhgpgvirOi+5PfvK+gprOWd2kBRP3RHx60iFZ9RWbklgZmwcxSMcmuZKL5WGxWLY8erdz
4YnUkoyHWSBPU6RTB4TfuMMNKoqqsOft55iZnBndoJ4bq5zju/22Hzze/Ptwxq8KPUPpontdtETM
njBNq/vqRt+splSsLiqztAVo23rt2YWemoNvsT51WxNv5JRhfzgdkGExPqwSiYaIW3AusTEj6ctU
A4kq/ETyg1MCPihGznUzxm831/iP/ry6lI+XJ3B6rg0afLwikJPrlFPumef7dazmIritcnNjQMnI
o7sU0q/hry3QYwIsHqyl6GhHuC3DX5XMjO8i96knpEGcLlXaZHQ8WWiEPKJWYttH7r0ns8xhbK+i
8gNHqnkvA+yaxt8ONhBRdB0eCB488Y8uZtsEl5WQ6j+ulhhB4Cv4VCfMrZdQ4k7wHkc6QWIMvjpR
WtJYPuJUjuSNEFKGwNFV1PkYk2Mvvp9wHYlEqyMcsmhK1rusWkerFVkhfe7+ubP57r8Arb1661di
Cs3ZPlP0oYrc9B/rHzObb+VVsBTz5sgoV85AlnR7FZme02ad2ZV1Gh2xUjTMo8Fv4y/2LjMFN4iQ
fBq+PG51T4mtWt2QRx0i03JIxtsWWqrqNvAvAPdW75HXclThzPVVUKUxj7Liv/JQKLnrctbDNczh
hMR+zkXMCvqvhjwyG2oue1V5dnY8cLjMI5+WIJB2pRVevPQfOYBhqLxm55a1+7jqAQGeoUAEt6S/
3F5lsgOUskNd8+2zB9qXCTZWZT/uFDMji8VY4kvNVJsxsvkiCQuh3D0j9lFV0PuM+asGJxzSlOxn
vX/SfqvPJBC1tSlcg9EfmpLOHqKGx3XYcuQH/YJUKx8wkeQEG2EqOTHi7v/mTMsxu/EKmBTZNgpd
mkswSYc4Ra6ix46qyd9j0ARy1wicjUyHHFDmI+r4s2LNzo7Vq64wVnO4ITBT90/TN3bvQf3cbllK
Se5RPK2WWFy0sHFSApdg4ME4N2QUJoAeHRHN8og3jGsYx0RiG/Zj/stlopk7a4QwZorfW6ITroY6
RbLmRYXsGGUWt62DqaklXbb1ytUq1pPN9p+v0ySjgnL/pPszbZv1WeO3fQbNIOACmm0jt2DMWQTW
AJFlifFpnd3l326P6T+mO1092MSdT53oqjP+agtEYNDPmuJD/oYbnRVkLjpP0Y6XYVy9oDAHJigB
iCORL0XP5CyLWu7haTVdOFqqV3x1z4LHVwAfqVdKRn4DeYmusZfENOdebOOjHlhVsNSDVEdWo6zo
91K9Z8Yfy7Ak6vBrLTpMgqLgpsD7ZsrC5lYBDpJufUvOtJGDf9o7YIXKDjPy3THIOifrxLMEAom4
ycMk6dawkaNtnpzqpl1Bx5vTTMSA0gKJCtN368brsdykE+g55YH3hmLrqoxQ1hLu/vf5yjCVhIF+
xfoTMsjJpyKJhSaNAVGeexYFm284F+5g5atjt1yqF58bjBD2a1pq2WoBxlTlE2S7qmhWF1BPZNGm
uNn/7HC3YWOQXo6Y1gTmyURtDfndxzaJrtjcPy9+I3LXXdckFzP9UiNL3aYiDtqkFabDcfzgk7b4
qv3i4xtcbRriJmk5/iOhZ+I0j9HgaNMh7mlNcjoCK68T0q0TF5H7Usvcknuh+ZV7n5uw+dA0Gxo8
fXmUN9TKmQkHo0R4nLimY0X1uX70QUU2yp0Xz5oo0AHDE7iE6wEgXThiR3Hx8eHGcmVeOFLeWHiS
XRZEOAznGJqVquKvMgx/Wxq17FpptE1rbr4o7wpUFG+ZZSLKeUdcfogUvBAyltdYr4HF81xJjgwd
OVGV6KWiObbFlSkequikO5DBR0ECQvquL7ApPtcqc1EeDU1wdn6gvEEfkS/9XAWhOZIddvaTV15s
fsTjCVU0eFTa3VcQ3GUPM6L0osLRb5AdkFD3m4/ucKt1rAMgUcxUR+Ohdvl8vA+Wsu/x3iHPPTmr
SEN+Bt3TaNDjQa+424BYNgYIhcxkFFtRIkez9fRMyptyvTwsj614IoUBaqqR0xc4W9YzY4QIMKSt
t4/Iz2lpCERbHfJeOsaHuOMPDIh/fDoI/FWHRFGM8e9UjCeb8ho92U9ygiBUUO9Fi3clLLbBriRf
vbpVdG6JCtY/ZY3B+sJcB/mky8iMm7Q6QFOInYGr4bE2vniRVPErYsz3j3/xPyxp3sx2B1VPyCRg
Ooe8xIPgF/mhO+Iy85szGOqj9ciLFjC8D6UTDYWbh9Q6BhfxkLNyzZ18LKuZ14vDHlsdXkLE6YA/
dNtaOZz7R1Cr5J+65FmAE3gncMyx6M15lKC/qDW8+FDqmCVTVv0FW5uVWSwyz81iCaB6CFiZElGb
PA70SN3SQfGsUQBYcu4RazFU4jRCx8bn5eRaFnDB7ArwbkV1RkUqq6sy/A8SyWvBK22iE8z4tpvB
luK2rzdkgOyDpaETKXdHEO82GQCLoghCmM7f8XQUGnCC1TRBPExr2w2D9VtldJv4KTBUAQFpkmCr
JS1Oc/2RfVICvXoy23Xp7Cdcm52auFJE45mk0ydD56Vr5OzEmCA3UPoEXqlXoVn0rVf4Pwr3MAR0
WkYOCRdaJqh0qt3MePl+APq7MheoiLjKt0WbJKbSzC/Y/LM/E5G+6BZraehASraj2ER4CGsVf+9g
SKsUlq3C4vNjdfqhos7PTVe2VNTvgP9rOJFT8qS4WnqWvwheNhmx+KjtJrFwnfVAgGTSw+pTLJZg
snah8mOyXg7QqMxwPwp8eSGA/PEyv9+rEbcfPhqGBQ9cS0DlJgHGleBE7Pm14zl7paYGzDCljqVK
wH8jYlOJwW8aLPhloVzJLN45nKVkvjPwR7W2IkuhkM2A3BuwP5VOZpnqu4uD/FZRJy7RuJj0iPTn
PzTNtyGnm8xzi3cUV70e0x5cGOy1RPYqYa655s47BYv+dl3rPwO31aDhzPc/b+/3gGt89cyJgDUs
55NN9sBPcOqL6nRfr3TVi5KS6PQKifLHJsS2QcSzfGncmnSiNqh7v7O6SUYnd5k424teyOSAskyf
yv2PB45WiFf9E3Vnl5mNxsqYm3ANR1FQnWVUigbgyGTf7ZoC4OWeeKHW7qkLchw0otIYThukahcz
DFEAMcfiM6CnINRUitwglSnSrXfOo4Yj3vDYLhVJEohZugRN6u9J+u7QDgaXC/5r0ywaEbvBVE+U
M2okAqtcEkCYtdVL9rs/0tAbApWbavGWrT3LVt/1yCGecYbfyWON4j6s4NUAGydJhSu436HaBMkL
qJPNlCsUZD7H7z5n2BkADJkDlIKhzzEAte5U4RFa1NFy+9V+KbdznEvh7VUajtI/vqQTFptdgZhZ
ha1ZKqzLNpkjQgs1w9WxZwAqafxuj4tH547zPpu+sUdTevCABVn8CWub+YGQ/hH3zm3I7PpeVYWp
ImAg7Ot4PU88y0FFE6fYMM9PXnw5AlZyNNGf6na9SfSQpXCLZMoppD5w99HMNHAVDsnxB9HYc2UA
xprP3kLuGX1HxE9WbcSO5WbaduqAiuZtGketFtn/7ycwT01hgZSnWnsnM3kWlCZIkPJhVB3KxSAb
Vhy9Z2cmOmJOiCfYVrUAs+CLcJ4IbNWwvTx/PxOa6aB7IuGuKDW4zVF7168FKCLB+ImzzUMTZNh+
Tyg2r/IXcaLCzUg+c0JLL4BsT6Uh+2GLlCCtr+Hj0KqM8rHA0oqDL3H5pO7VOq8qpDaUZgXIDE4l
yjTrcOEOxfI3WSPNj0GwOJetElbGmGZMiktmS38JmlhH1ddu336/o5CQ95ob8Sc/UAdWcNhMsvNV
krtp6pIjnaj5iUTBTTcn0NzVsV1chGFiVdaUikvQdb7mkXobix+R93n+ywPjgzx9pAcOEYorh4Y7
KNh1iDHXt+6lYIbHjI62p1EbM728xjTqtGrQKanxLinyM2JsS7HfeJ+vaJ3sgMIHIFWs9zrs2dLw
16YtpFz+S3yL/zka7oquugDz9FzbNY78Ua2AZqnnT4/Wb6G+vV2/9e4yWln/hA/NIzpOloe3Wo5Q
sQ3ZdDwPf2JPc40GTrLAJgN+Dv4oyDLFHDuPDJn5ll0d2bDjHlO3lOlx8/zqsBWUjaeuQJMn3dNZ
BUA0f9aKYhliAhXpwjHNltMy/bMHW9k5gKUvB/dX7FZwyFuEZot0Y/gg9bHdzbUxEaFdTIOi7sUV
8Ea4gpdjF2KWC2MJNeVNj5rpzNJh8I3eYEG4j3W2IdkYDY4QhJw+B1SPbenTIlhNsS1yIKUmXw1c
0ptOgI5R7ap9bsS/cMlPnehqG7YVxof+HEZABAHCG/1pTPzOQBBd2w6cjSqH0dvwOI74b7uy5A5T
P4Yjhq+IXtgDJMedQIT0PI8NhkfVdHG6byM2GMzFdLPrtQRBFpbNUQEeJsF0F8RuaPSu+Cgc38Rf
FYNq+YogNkdWKEorEQrApN/V/BfsINiBnY0Rijim+ZSweEMttTt9/twtEfX9mQRuV69O0M5z0dnY
+JVRAlwfr25N/wxxOzXtWHqKjf0te2zlnU4rc0Lamb2h5Juj9kcKHD3sp6s1jdxE75mJyP6e4+0I
nbVvwl/qvYbXZKo7VCBi5OyEOhAPRlKexeVXm4p7gB0RF6MDJF48J+R6MOMZaqA/L7xGBbesYzC4
0Lvghs5b9HJwAgmCSt95AqfzJIjRTnmmv/HwaVEftl80uDQ2L2MSCdojyo6kGYq2ekwPdOQzPPFp
OcerwhReMPGvF/Gkdgk1f36IdXl/L1H89rsiyFZ+lLv157Wq2OtEcM4AxWOcaSBR6fTuN9AxLqyR
9/ywpeeSIQSV6gowm9PksdCMakMw3CfWdTAWf/xJwW3CYOm16nzfL03eiEeEc6OyCWBiYoWhCUqh
FCd1AhaNsUOvvuPeNdKhpi+e6/Hl95ai0QkZsL6gFOlEV1Cefppn683Hvdi1PnqVYX4Zbkk7HROx
qr31qLrjccQfrstq6hexGVQ4UjzAzw9/GCgfCZIFG+eveakDLEv6gJ/ngvi0Zjn7CEcJWTEXXOE0
9SgXaTVZkSQmYW/XFlLM6UfBXVaBvfjhI9NjpUrEPExJ3+hrxvO5vf1vB9S52hgEG9U13N8yd8nc
qTbZHWR1i6y6wPtmB08LFLbeGhXILdjT9kpsa4x+D9UBuSSLuvqYnWnkGjaA4VJZXy21cazoiNhE
YLNgEXGv2oAFB2sRq11ND+od2iSTKygEag2l1qVMLxe/HvphSMyx+D/RlyBZ/IBYz1L78aFlCwfo
34vpOY8UIOkMRP7lxQbPg29xgoqA4Hn3TbSHIhlpyxVEipbD/CxyEC3MMBNg3iDrPxpbQvLWRRdG
/YsMybAjkpuMr0sozyAWl6UWgyvYRX3Pmu1IWoWFXdYfncxGAhWY4mTZP9RjS/mQudfUHwsnRNTc
0a51r5565qn4B+sWBaCVulnPch7LRR5KroG1yzvCKW4YMoLAswZBP9h62yF4HChWtkWemKiSIdxX
ECQzT5lsTnTLPlX4JnBUyfPUsCptEYH8xaFYEJBfg7+Je/Mi8WQGdq1cU6SFauaYmESOrmsewrBD
H09I+3WVyiRTrkf0Mb2aGldfF9plkbUma0FoPXW8jwZcfLuA++VHWmV+SLJLj7ER6iUQ4hQR+254
KSmA9pstaI+FF0oDayWTQgi2U3H008pEOXUnAZzPImdH/Zt5FIpOk4KXObTDX+T3G97UA4LCwU3i
buuKpyKvydooJGpM3O2FjfX5MaKCmbZ94AdZl50pqe+U2as0YShj9WJgGiTGVDgyijXQes7cjtTn
hC2XXUJvvKvl5uIRNfDgnM1VjYTuFit5JQqzVFFRG6gP7B7T/HfHhQ6N1Dqx8arUJMGaaOUKllgP
X7nhsdas9jhhWpZVHzrBwM+NSLGWwADHcfr5cggWOPsCtsBaeVKy5U7k7SQqAIOhHodzslQsDWow
GwDg4Mado/WQLRS8r6gemWkVgY+WGZ/gGTFZ9ekXyIooY4cBYlu0ilgQsef625D2yPNf1XiSYdce
kG+OxoKQC1GwaYP+Ff/dB7zxa9YvwRqH7USHzM8bjqNBVpPIa1BskTjg7lV06YNrjq5+LYVHpFK2
+ERDWjjzsZNsu7IF6U+ULRcwI5Oy+ysshah+Y4qAr82q2PCzwelBbe7CzBLpyZWktPOBOa57Gwzt
auvKpErxV5rXfgfPjKvLd54tF1QmtZTEDtc4k7SDuQPw3FLrIQWm9GjUmeqo6rvNdFinVSsggB2H
MqkZPFv/dBE3rCl+LNzzWACF6Ds78bkdyWulW3G8kCg34W4PxrgSKj50A9TYdG0xTHRs4dN1lWxf
gnkivwXq5fEq81L0JcnmK2EhJta3X8wLqEvHP9PLJ/hkR7bpVfMGT1I1NuQSh/y2S76MhbP40p3Q
cHjT1W+Cd8yHZfTXr3J1OhPl86S+Cxznr1j1Fe3FzcyAbWlNOB44W6rmY52S4YUzxZez3F0KNtT4
cBkrCO6alf9D6WFZRDPrKnMYBFzUEd86UwUixaOGJLJ6kg92l2p5yg4yCodrMwpl9v6uzHuKztlw
XEkxYOtdnbD5HqYXxyFpcuYUL/qGno+/Ig9iZExk+mQsudDWgBm/iH1X4/j7tUwGVCCx9XxclDW6
vh3lnp37ChIqjvfJSGTmPu/nLMZ8sJYzQ9r0xxxuFQyGdcU+oBodgLPH5A8YKpBsvgBNebUMWiT+
epgToKMNoEXu0ZqoqvZB7wfgcUQQ9UPhOPvjqN1g4oACba6X0EH3Ki44lSh77X6Bx7bmAW+BjZ2G
zpizSLybjdqSuMiJCl84WFd/gMVIEYHB4irFJcjF0Selg5dDG6UgT4JqJB9cqozoQq5qoQ1CoKNH
ctZqkyP5f3A5mfT0BKMdVrI/yWwM3u5amQIWtV7xGs2nJHIKmwfy/T1DozTOaQu9mpuEuHB9IWPW
NCLeLSoGFWqArkrrTWd5vGES9WyFdsa3x8FppI9Yv6wwkyR+8BfcOE/JlJx0jlG77EpnPHKXO+TM
Z/uq4oaSLuJYUgxIENlSig8a+NPZ9WQtxse0elA6C110YW8KaP85R/DQOLGSznmVB9i5gDA2O2iz
hpMhR8zKvsKPGB3efXDWKntoQV6oegHTYo+y6hSBomfqvLa3x5uxcgq5j3lwTy1aY0DHXbh3r2ZU
KH31cFYPCLKixoAp7HOHsCks6KLsAx0cuqJPkypDkk9GyjMiwAAXa5xz176Uo1+ACgduBBP+ZoAZ
Vidhux/mOYS1UaGJPzKorswfI61EDRGc0NkxZVEB84zSZh1XeH55miIiId0uDNlaWVPhGscUBEzb
84+HI0wLk6llobX2DXH0Ccn/fOa+wSbYpiZ7klpqlryStX4bynmsBEsKtYmtQJfairiVv8Osi3fH
PtkqHQoNX+4A4fyjoDYmyC9iFoMiOIIK9MLsh7G1BDcMaAaPgcYbjDUH9E3Y4YJq5PJ11AAN/tPk
aeE2jhHvd+GlHZpakRtRIeXlQDoMZjIVUxEsEgPqcTlcqVnRtfwpEcMPtA9IbadwBNQHb2M7uFuF
0JpSD3QVT2z/jBj2Zw6JbhINNG3k3xXBtCystMyMCQ+7EZqyJF9TsTkzwG5iEfpKq5AYwno4pzCv
Z+gF+8e+UJngdlQhWPC+YoTGwn9GnVIy9CKa6+aRb2DcrXWq+Jk5NOewTdKOviV2RzARNiDlezPs
8aD9xPcP24hOU++OPnjGLt+uLtaEsrYAePn4RfOTwzI90rswsPpibnt/183CA8aRrngfVEwRzj+9
f+v/MwoOOIqw9VVlsvu12kWOPNEOA57rAX/AmUXOVMfW8lr8l6JRPpWIfutb3zVUoZCURH3RYQWu
oH0Mf5YCoxIEtHXqikS+NwsJhyfQrBjkLa2MnCYI7DVk75duGq530bfGB/8/NIXZ8Xrt5HqrPIYZ
0Y9mEojDSBl9PPPHoCg6y3JMb6zp9hl7z5uJMzD5KTr9TgXYBKd0rKhkmKskSiMJSjtQzD4YRtEd
3VbLDRe2cdTgvWw4fFlBlsRpNticEtmHfnSVWqVdMXRe1CrLcoXlnnCZyjZsQp2f0p1v0VhDHaYO
9X2+7y+XKTAt7ESE5aC6QERJ1BrK5+vDkSaW501AMBOytZLkNwXXxcjxQe5jhp2TyQjG23SgWX2l
oB/2tYxR0X7TqSFxt72oOJayUy2EPqhANDNf6c40ZBRrCcaMJJqJLS11etABu43D2x3IZpuwodSg
HXqGJGeDt51k+LyJRsFx/Ap3iGnGW/U09sT3b3Am1PQljg7W0WrNpjw4D3P2PM4tco0kH2zuDwBl
+BjJeopF7Uk/YkkEj5z2eKKitMNuNDmNagMKrsh2yC6P3RL50Xb+bOU3lOHYMUSOYTsSLCX3KHIn
A9jHmXZFUGnPWxyBGqHXklP/mPc6ZpsulU7PhTCJbjeVW8Ro8EnDL7MALNcb5JfXtrMJk6tOWWFy
kAz0RxRxh4K0v/Dl5lxl3bidEV2SOAHZ4jqZAW+rsuluv7iP7O6QOKIYWtnP9igCTbjUCNYE7Rqp
WQdg1yyPVn175WGx6Embps/tAsaiyly0BlY0XlpZfvF1mH2yO9o1sjxcG1QPeFvlZVIIrmabb7a2
HXZ8X08E8//wxIoFS6srdLvhMmJB263TkzlzLS3hOsLVz5jTl4TP1k/8Bo/9ZZitbC8xQvaPbAvK
02jMBd5lKLnz3OI/8Vt9yK/SJGDStIaZQbZ5lU7lAnLJhMUMflLzkWK8NEj/X67+YJVFK1cLJB9O
JcaD/Y7I1bYbLsvRcTsnG1rNNS+4nvRpSCnS0y/UpZAHvhZ2+heY4jCvBHIOGrEnfRLVPLZHBwCP
vZHFi06x+Kce463m6iTvg/DNteVyxv7g368JRl7wM1hjyGzFW4nvQWW+ceA4lZuxKaTBr3It2km/
dvTIsuD4U/G0pxJ2XuziGzR3ViE8M6zK8DSLCN13qb0DryeuToyxUv9QJBxFCFuB6oj2nzAx9D6h
81y7RqRgshjM3DvyLPX+KLp0MHBom6ti1f3B4GvNT4xAJS2Jl6KY+560Oza/aX7NtrPewAlMNY9g
rTEd7M3WsehVzBdB4C4+wQvvp8rVUQ5bALyyMz7EVmYcwVsmJJ/hBdACjptP8/yiFE18D0vEHaZx
H61Uypxgip1mvuiPtI8bISA+ADoufadpNf68qeYwCgCSZJIa+wNjdr3xoO5chgCedBtfIp3o5zVZ
u4/Id6QPSOceLGW9xCXdSmhme3CZaTBoDbfVZsxR6qoDcwlRMXk5xF9NK2g7LqU0UadrAmN1E+X5
1Jsaor4V8MYGe16ngTccKh3aZ08KR1pnBGSjIzyRRMbfUzSaVUOxcV6oUHSCVB8qQa9tKBhDd2e4
B5nWhm9b1B9h6Nep1sxaznxW6h24heo17popRX3vyRTqETGMlN31JqHolFIf3qE2DN5Lfjg09snn
ZkFne7pImQp5BkWYb3QO6FwYhLWrAtMcSZFbLIqyv1dE1Zgv7UB2lSbkapQS6qBOelRbeOposgdW
XojEeHYv4yXGIVytM154or5wGmXeAwrcdqyPJsggMGQknykkKA6fWV/01YYsilTec0OIFTnTQbUo
je+R/m23vNMGJfyeXhGDz6G+jvevx+mlTdrvbb4/kiJThk9BaP/WaoFPdc/rbf1XX5iGBL6ZAB2Q
8D8u2gxR3XJsSOI1QnH/sSJ9ZBnzaZcx9D2unqZKmcZvAbXZW6hJcbUcgvnphVxgRz2pndl3BJDm
cq9aNeNoMpOnl9iv8RUrB02uQcW4BU2KnKT+Qb2XmnlQ0Z7pdR8SxfiPsK0kLeftLyY8mKLyyE59
Cgm9tFWQIntj8Z1uIX/RrvPDOy0bVaavBao1dNZ+2iMzmwuLHhcGY4X9rc+rEZX2+ZVBH1kaSXgS
j/nUuV/9/PCz2H5v1oVKwzhacT3ThotTE0Yz7S20a3fExX19IAALLsWbgxJAUKajsM5xykLpFix6
3YvxlKIUqtlBlOkXxTKgeTfzl+ksMGIdhToUCIP2ZJkc+rOP4hmZ/d7jVC6og79p7c8cy6hxMqFv
PSLyIFurzaX+H8Vg+UiTCCYaYAd/qdTWBr/ePo9Qjph/T+7mUkvukslHklSEwrkp1LDObvry3wU1
kDYmwvUNP1aQI6hjz3c8TWjGAaPvDBlHd48KG8tDM+DwlWo/KjN7YCl1V/OmH2xHxpLenOMM9vdF
cw4Yi4bk0XFGYt2fYx/HK9wqQtOe//ycFhjq0JRFzPLvN9R94O51wkDXxI7oosma7QU0xeR7NRf4
x7yVWsJMsCzGAaSeqQo64owhW0h9dH+rQq8xcQNtOKgcT4YgDxjqBaB1DgAAV2+fTY05K4dHt6Ku
WQ0q7BVSCr0HC6YV2zWwHYoy2CuvpHRtDVSwvqr3InZqcYynxF5aupe042FfLWmsQnXXFPW7y0h8
b5N+/3Yf7Txy1VADMNf39v5jFfck0x35/KzpFyz5YFdmq5KFuXGX2sgFOcbYHx+GLgRPRmDJMA4y
ekHnVdJASc7FNHQ8h7iC28VaLbbxf5E9eyYmMv5p0/3Q2AqgWqxrkMcWaEHhLnTH3SAZgDxtUxiZ
51c6mq28tzX9eg0g29wOl00YysSMkSM1Vfgf/clJji3RfiDqAkO7+aQmbNTICRZ4LMO9e9qKc+W5
MMZVd/x6WKktBaY6ho8gTlsuY+0W0Dp7idwz3VqP+AdORGS6f3nNFaSVeaNKOy9UiEzZ/Xba4gGQ
7fBbOF2wn/vsVJhb9gHzesPk+cpOPJDrdr0xCYv6n3BfKIoDhMIPLBB8GBwZE3nMcCu5Tpv318jp
atWPJsRmEO+tf4G24OJH4zGA6HxC1CSwR8v/aBb9yS+K2lp2GhXUXq3JAJTCo7xlhnFCwAMGa81i
PJR5PLMcXmucad8P/l0GpKkjnE7+I9SJqaOq1OixnsIQDjLkQQ5uSk8wUdo7hudsRGEwRKkAcmAN
bXmETO3iu8sawpL6aVS09TmdsrIPOJjksxErewpof/jlWzRdeRqVw1ThmOegvUDpsn5AVDtdGLHF
z9dDpWLGh+EIWoASPMTDbAavM2YmiIaWevG8FcwWUiJeC4lmHF8iDlbgvJ0TGbI60cDX1MvD4AuU
tMCDyDmpDEC+UnTX3OevDlILWCVy4qdWn0HgAGfj/QEzGX5yWVtDShzBNvIgY8FpIq2v4zo0mfdj
UpJSrQTziyFEfEGB9c7W6P6vxT2wFkT9H9guvQO4gSgu66PK5l2KIwVpHSuLmEBSHFksSXm+5MAv
g+jRx9OrZLIrsjZ1mFDKqVctZdS3SdahmZnboNcH+Zv8Bxrn5RJLSsEqNUXQAFaaMoNuvQoHfpQd
3GzRsB/IYZiC3eeWiPz8mP4EVQUDQTw0epnjCtguyJSW02s/HrFFKv4gketxnonD7tEg9ISaALxh
loy3wNWFL+k3wMd/xNO1hoMCh/zQCR308gdx3RXOJrfHz/jmOMBWc4+ITDpeeSWXKnTkH66fq/A7
ztOUIK/jD53waQUFed8lMkkpf4Zka35gfBEgd1TCtSE/OZSs/BALMaui/Z5UH4QtJ+HR9lZAedpV
JBelL26PUCm4OKGhnd7lXtZmVHXJ1GaunNJP93nFfSTmAXTNiLa5/L/0lXdAXSuq/f2KTmoflBa1
vaVg2x8vNR54baI/ULA/Hr+aY+mTl/WLEuwmlV+ZqO+qGUl+fpT9uH7C0sI9x1I8WilVtbjgY+We
bJxS+b9xLo1cyzUojO/oGp6yAp51E2KCEo/bd7EA8BddsMYMpgVExGDrTY5cupSM8tDKjfPq3dkw
QcvGGvVC/Fkbcvr98mAIYReKUa3G5C62S4d3AabWZI08H3u29FSZogqFrw1+43df4Cn9rXTwO6kI
DCgoUtiDCFEPeiehbeJrrlvOnAC0ihbobwAeqA41P5yinu2PyTwlBlVv/shma7ovNXcv/ATJc0Gu
P9f3MreziBTGf2pql1yKhk6tAa7xBRWzGFbLrv+DWUUF1V1DpDnC+CwFS6s7fy++oGEsXO0RYerM
7ukzbcuQPZiCpuRy5OPwGKYpKaGjSIDpSnri3aSGYP4Gg3pVeCn8B9qUOCi2X2p0rc7XTsjHakYh
opQjLJ1ph5plzNqXPKVCCAbPLzeLP6whijjOtmGjIu3UJlWlEYuqbLgljLMjPfFldkG66bCFHEnN
vTW8FMoDgnpJs5r5pY2b/C18vfRmkWmpML0E9JPMM37S4/+usJdpO8MlPr5QQUDrhWyDpPu38Why
/vKWN+mDFqkd6fgCnt0s+F22oP9JPRQMjk+WLg6AJ9GZG7LTs0DjohD7iHAgv73cuFPQgUUgt7ba
5ka92kTGldZqsIMbO4knDry/spG0xSR8BG76jXdzgvEGz422sr8CofzURDllWkkyTGVHyHSDcZYp
q8CEB2HKdosbub3uEvJ0ZHO86tE6H+i6Z4Br6+sB/Xn033tgHQLuUbr8SSdzI/ZGJ5bYYNVOpQHf
6uV4NAjZbapWoJ5qyEvovAI7aw+RicsGG5lezvXqi1w9dn1mP7tLh/Hh/iptniwTCqGZ7W/WjG2h
yoRjtrqBNfijhhRI9QBacC7JgSS+8E2Jv8PlvnkdyI8CY+/WWS+pzN3UqMY79pnABT0+TKw5BGDI
RJnxxEIw5biF7+w7AD8grJ8IrBRNe0FK6zYg80I/E1ivywkBZcTFfvAeRVsUXHAqpxY092SGF8Hp
Q0bHIXPsYkHcu36S+XYpSE131DjkGrx25OH9V77bmrBfY8PlqTP7QXZQcAD3A0I6p3dxjWKGADMO
KkY8qT5GV0unG+crMNnxHJKlpSv1i7kqandzldHMQmgT324NecaNkuGJ8yMDy02Qlq/Dl+mdWx1V
NhVGvRDNVrbRJBugk+9dZXFvS2D7NzmNYrZy+94zcgY/S3qJ8adYGkN7m3CPlif4Smc1uPpiMKQc
eGzoK5LAcKbMcWnsqRmWVXEldJJo2MgPsfAIOq9Mwt+LMarHtg0Ck4gh3wlZllUo6fAbMVyASrWz
Ibbi4tciNr18gviletiNtP6amJW+zBzNjlEMpZ4JSTxzeABksZCd/Q3JIdb6Vi0BEg6GT7kAhGEn
9KMGEnQpZsQQuVnd8L6lTRI/f2xe5t5qLE3bRfLfAeaCwOERGR82tSsPIoy8nDSvbPgIhJEwtNlk
KWxJoOjr8PaqRz8zE1GELp6YKS6o297RosSL3OPRFKnWza4CEN4gtf8ngZymmcAA5wlM5E+G42eu
bHHq9VMEDiiqyAhsaLu2nA1ExYkMNMtSsduL+iAw0UX9tdy/PWtSuONr0AIUv36Gj93dmyucT19N
fZisAfI7SDP/iyI8atQdbnKLhjJdHeEyB3cAEIsnSb3629FT/k6/ua1Gg0K39JbJfN0G+N6DyszU
XZ5CkaXJJIfpF24Y/ni3IsFB2hrUJQhYDHxw+NhWjgjMC0mjgOHO84m+do2rkf5yPGzNrDkH5czO
XTwG/6zK9j7eMbCnfprSie/AT+sKoD/fQQr0Or6TnI7Q7l7IQeRqp2jRfcAggKdIwvQCWQysy5Z2
4kBfjxIB/fXLTZHFrRgCmx50QjvkIFZqVXkKZgZfcABKc17L1O5pOT+yhA6L9R7NgrP6sSw8sD0g
79eTCEp28zgEXPn+iXeKD/lyMjz6xFae5FnptjyRASQNcpicHeb7Iq3XvQxGZeUjbJ585DaSYx+D
NXdunNVAH7/IuHaF48hr0ScrdXkI78KgOxyeW1JlNcWe6BBTX7M+jek+zf3KnRc6tY9C0q1AgqPk
RM2+RN/BYpYTEAN8bb+RmzN6qN+p78ICwQ70cfhkXXUFLkV5rkRyNr3GvyokZFdv8cBLVo2FSex4
jd3zZWLIkohTO9NvhV8RmSMdtAk7hbNye4+GNmws03OEktWpeaihfegv6aqWlNN3eSVt4yMCxaCG
O8prtzC+GARcTyz5OTwT9AV0vs0O52EQ0XxUWwWfHQCAEItY3PLEADzFTBLUex1RUM0CYBjK/Ke2
q4Ccyv/PrUhmP/vxDEAcFUCArNAvUoIsl7HL1RKwNCOk/NNF9ez+i2koNBzwBXMXXSlfK3wtft+M
7wSp0h76rp3O1AQ0wXmvEOqQcizq9JwVSBqFBlWQNRatjp+NTscW1kx1nFbpfhn/U0TRYXOL806l
fb+RS8oQHdFpds7Rfh3E5BvTjHp/vW/IxD6kHfvvP4WRi/4gPk9Ds/ez7zXira+eGa+DbpwmAAIe
sSM9XhrrsG5xPZ3tPGiDQSJvM8nhUcC7pIdixRunBd8yWwuNwnpG7KOiwY4ChieaEZs2edYShQVS
OQsOS9Rk8EvvAJJW8EsgKSEWKYl4vK0walBKyST5B+gMcv/r6uTHhbgzWpblJIJK8rljkVv425i5
+M0NpiDQHIQJC7lmFhmU1JpOWQ7doBWAAqD3r15dxgO06FrAPNjkG27QEPOsR47HJlr4v1Y+VRAm
IBe0iX91POW9onlOb0VH2SmQrFFn3S+5qMrVV7grE29AhRx8Do+Sto1/Oph1EEWMr0lgESWwK6MM
5D8DZctD9TIAq9zvz/wZv5N9hHGCPSse0bt1MP28L4RuoXEXk/CZVJPZrj3MIF7o4fdGdDXSChZH
Z+3edM6YwcSmm/aDlcCe9PKRAFPcCdbAr29n8peW2EAl+xIWdjUMK2ymzJzewa2oGedtT2s1ebqY
PovB1DXIVRqLdPYjHScielTvwanHFb9AqWlM3yS+mRLPWU60Hp2xtCV9NXdxEqe3VDoMzrlptuN+
q0XF4fuOUgoZUCozoJdD0IN8uALym2Q/oeMN8+R1RA5uXsWtgEkPVZGfL/V+yliaHyIX91rubpQQ
e7iEslipZuU1G5/65RAYqTNQz5saxipmEye6PkEfeBPuTEojSgny/dgQ4AMfbkA3daVtc9iUssRT
iZ9G5wNodEjRzUsbZYKIdfNfXB9KzTFxZY8p3WZlD7Eq/LPRr2f9wTrVzbLR94INJDY9tfTH1sfK
GLuGpB04JQarNP4LW2qojmTaygk8Ck4MyyWmwkjgLsjpS8m688vS1QYS9/AIMBIhdpPU5pSnpd80
ooSr58iQGs+w9WEY11bJdlIKxOPzIBCNCC5B/ImpjcmG6nZchyOWtOSsn7v99WcPIV8A9UFB5RU5
TEmmfVxa8GdmxVvGQz/xtMDxxAqXZAECXqkJ2cxFAcN0n51VAwr+o944KxUfwgdOMvqGkg3edR4v
C0/h96RPxKpqpxVGNVU/yAg/wsEBO1/DJub2H0dULdrhzwcvjjP9XlImdizLsbdfklttuFWT2vIi
MkkQAJaZ26szk6VOm+mMw3BzUdfArY5XdCblT3tAA9S8A/XdzD9CMVp/L2RRvPVFoTA0uM/4RKLe
HAhLMN3c7BcaUNP8kMr7EeO78JAw4sYtRCBZSmKFswSAgWzb4JmX5/n7lgpTBl0Zr/C1fnPetaPv
HxX23bbI4sRBfeXQiK3JSTtF50PwEZ0cYPOuzlSRc8bP0ANOKcjIDGE5F24jr1vlu1hY+oSz7F9R
MRWMbt+YOKtd+3cmf11BTEum+5K9sUVYt39hPGTg+A8GfqJ7wwdVAOkfWFdVcg4KM1jsEs25Mwd8
sddS4vxKuLI7Wbu9j1Nv1paNd06nh7d8vwZzMhtRW3cJd/pTlzcooXT3azv22bhtvzf+3LSlb5GJ
Ubm/0fmyA9cMCSl2DuVPJL7/nGszm24dG8h0RrRutb8+NEVmqwicYsE11TfaKG+YVGud6HtoAFxd
c30nW+ZIYO6mWblF5WpeIiaXNWy98Yetn349DSUOJS89UGAibVYZX5Lap/XOalHFYAIcNwQHSXEY
vxfxfJmW4hAys/9cyIqT2jvfb7IAJlXtsOCYcMNSjB8tsZuB8JQN6X8AFsPvOt4j9Y22Y1xUeFRG
Sa17D19S+Mt3ej7BpKib1FpkvppWbyVXOLpJ+Qe9VCHyBtbXqnzXvBe1Grc+JE9d2i0Dfbgoylm7
VJEDS1IoWJ4TAYTqCConB2N/fzsVe4gMUnyPdajxnMH5N8THXWKr8iZwBMm9mf5mF8JDU//zAEP5
zbJpuPC3bHb1TKgNrW8yFp3NY2OocsedaTIFKtdMjGHIIFDmSD8t9uB/Vi4yxoXBJlNa0JtxUl9u
ZYF685x4EucEZhTOfGcg9g90x3DtRs2Y6UcdEtZcRdxwoK3ZoN7DQEwrnVHtjDV7JTD0SfJphaMP
RzBIKwjCrkmW83tABdhqI+qUn12D5/hzz5C5qqVv7cb5tZIRy8O4/0fuN7u3WuDTPwFRMWhCJJAi
h6V1uEgXF3RJ49ONcAwvSZaHEHMMEEIv4fAzxkyudYdgjj5yC7jm1imDPjpK+sbWWtR0d2eAJFho
CtolMJYBAWU5sded7p7y5RzpImHA+HGWWotVAwl6HVndXGYRPMmV58RiG/aSeNgsCdVBvD5Zc1pd
bxS55s3KuySnT+RLPM69VXGbn0NBfXdNDDlsI6XcfFM3f7MktaYbKsoJGX7ta95+nrMnAQU2wcnx
k/hqAOSqXiBKWz1aDDdBnedxEhuCvOCuPY8gVve0MUAjhqT5ucpd/55xirLuZAZqIpThhJB25Yhk
/eSF+rziM5vXQhmEpF/h1XpnJt1CxGCMwxYU0b/6Cy2KvaAXv7smlRN0bMf2QMRmAyaJtEkiArgD
76LrK2+rhf6l4A2lWSR7Ql3KV4jpFO6fDQhrI32ZcSFkMSWHdfJy5iUVhnnde/4Lfpm5MWEdYtwB
0XOIjSXqbPF368ZNxFmihOYx1VHT1Pnw8xFShUVR64P28nvIvY0tE2oLzmpSDUNrg0ZjL646UulO
H0KhXZaQiw3ssIrjm+G0U812DFUKOJfLMxCbfthhZqfHHiuBwGm25on88haQH8fALTv/53sgSs+u
dWV+HywX2Tnx1Yue0z7jsThLtB2TZhUvAZAVv/zqWjZRzwy1JpQDq5zmB/RgKtpnmZFiLe76ruaq
a7QkQCbzZK+Ot0/aMjKcjS41ICkvOCIc+2jDTvXYeE63EsCrLElkx+FaMic6LJpeOE2kiZyh8WLZ
u3DPs1k8L7BShn+OKWYow95Z9TU8seNoMsj85sWBr0pLl1+fq2BwETCyDFEYzKCakp8RNfsiX33U
YzSwl/tHDryTJYsWFVIAGZWNEC24K3jjC1l2Pp35UCU4gnFsRFA8yfmOpsTV4JtNxxsI7qyYzYRs
IcejKxjFO/NHgX+0dMNNpRqutFKnsM4r9jkv7F64RlH89WVnWWZ4g5MQ1v2nDjhpKFUweNVx88U/
W94TpRZFopHm3k9zJDdMMHiEjblGHBMrVQ5BVN41Rz1D70zXyzauO6riL7B1v3coNAyWko3M5XYW
raYyE84a03LmGNm6Oer1rkZQ8NUJcnljzPyfKlTh/7sNOc43tShHifR5x5khcJ4qei2EiPGWmu1V
tkAAv2+YVNfQzn+e1oBGY5jkBQrO7Ls3iow26L2x2GHcbFK7mXeChAt7BEfdUqOOUQq9/jzGAYrI
0em+gDgWX4O8YdtBQPtB29Mb+Wegumo3SdEIJPGl0l9xrQKNONK4fV8TJwhEF6SVZ3HyoLd5GtW3
RpGXXutnSARbWzY7WgNL/C8sePmmRFDmailV7zuZAqah9mZ5mDrL01Cv0mPl0L+WviKKKBX2TxhJ
APx1GdeWA06azfyIfxG+h7YdiPpRH/1xxWPvwE6gtXgSn02ve6kic3X60E+zskpLrzVxsHJQGlQb
duA2K5UmZ6pP7UO/PU4hKKF6i6YAAktenekNdiVUK6LqHMJiBU4ZK/WK8MRHAKTxXZknkzXkizAV
DTTEuOI/WTnfzfyRh+cXgA9bJpjGsujL4R/t8NpBn7UdmBIDTxC1KUmNPJWrrh9JBXIPXlZ7owLl
laoxlTd7q4wKidyC+9aGKm0exkgZVX3vqoR6y5kk7j07x8+kwxuMUaMhQ60ywKtzl2d4VnC80mD8
ms8tHO6UgRm3OP7vnWFfOqOCD8y2Zm0XcxbaoUWPQ+VYo5qVIkr1r1bVi/+jdsdABtEm9rSD8MU8
zq96covDTDIk+GKwzT8MfVbuGFVoEcd1iCAPCN0XYAbeUcZbPYMpqsWfKmpzpVL++BCKwydoYtfJ
BmxM0l/jlEGqYeMvljToYbRIBm1kBUiFORza+M3aRw1YK4Xe6aY1o2FGm87CMYjBwXccDs45RMA+
ZrRESc29QdxrWoMYLuOOgxK1F37KT8IrJgzBn2/yPZvatwqH61yHI/AwhpsdrHwAHvMm3se6hIxf
+CkN2TldzijIfVTZbLEMxFg+PYw7E4nBGGChANJYS8AYtl7elx9XnroSA5O2uxSZKMYkVR3Himrd
1RfxxzP+KElfqKOIbLFnCQYsNRIT+yNxxDkDxKdnOE4Ma2oguokX34mdL/hocFHDIxK5VWm4ykce
gIq50IfdeS8tRGqiaXlCmUJNdNGq5GvCE9WwnS5XqmG5SLdpQ2zT8s9HjPugM1rFFve3Xqk24N13
jt6wsDaE1xz2lbhaoTzc83qd83fE8Ng+YcLp1IKor0n1BtQgMVX3T4li8aPf+oCgKRy0C6FPiTnm
SSySQHCeo5F+omjGOYkvj50lT8Exdgm0Ue2SqJUu/Zvy7GX4YE/a14sT9I9+5ir0O9kekciHbiUj
NmQb5Z1UXvZU/9r4IcMlS+gJV986AJ48Z/fLYZg1JxQkqQdb2aV9mn+MjXU/uImArEuHyAuZME0t
fUpKqNgbpX46OtlwTGbHp/lATeaoRtK8XpQ5EoN+rTlY2CuAiera/I+znPR3dS6BhWOrZlw82BpU
qbx7F6eXTSQxSmftb8BJ5ZNqitQlCQn3VNhFHq/v5kka7P1CcufQ5MBUgSjD4rfL0oC2pmX6dU/4
6ohNfHOWwDkB1WeIvEWBnq5qCGWVFidQODm3dihHxHMfKPKyFNHKxQlYVHzizYeumblGk0Cxpc75
aR/zNvC3IwMh3ZWGLuNKWXY8MoNiSMrNuIlQVXlXjSe5ur1rB4bmOlwrExsCsty6MQCY+0GCGmkt
GhGP54IZpn+JWLlm1LI6xaOgZY3gItQO31vNcbgAKE7ATZoybY8hqCMhpmPLQzSL7+axcKUAQYxG
40lEyBe8w4/TcoGF31Wz+4TXqMBwAIzB9zahISG6IM+TY8tvzTJXOHDpdo8A5xaw/eklcICT1GqQ
OdusUBLnWCQWW65ovWOjVjElNYGolDiwPzg+pghm3QTi5KtQ9PF7RGOKw8LMjRkJuOydidiCjHqw
nk9j0EhJ80ES3ahGGmkh5bi4y9PwzglcVAMUhah8hsrxTHqMZj22bjvGfzZFQjd3eHow/YcOAQgp
XstZylFqOywP1rEHbHJ/OcSc0KFgfPMJVyjhSQfPxB7PMl0QaUF/qVvVFmV943F8e/qvuEq10ibr
fp/1kylN71UBDYu/18NEJuQ8iF0ZIFFE8yFGGJRu0piMacdwKD1QXPWzvpmLRo6xWBZkJPwJGeW/
Jk6LE/hlN34Kl6b8C32TWmbXyOS92ZqFDHOIc2lN7HhuGw9hboxTEhX1Vw/upSuJE2idSldcp702
Yi1TnII++SgdsL+8HyNEDIIOWz2CKnOkWdZYzCCFOAZairck50NQ8cU3oT7QiYZeFJ2AcxstvkAu
S0H4ZUZsOLb7Mrdr8ULm4LuFEbJW6QmrOsUiBEbORKjJ2j+rznNJpkl4kQ+hlw1CsHQjZJJbymcE
FUbYEqtfVZMyFS1Eg7jSxi68O9uuvodaw/86CqJlBrPO+1s9pQ1IxdrtE7ulWNkoX3pYcv0+M3D7
DARYrDhvnh1H6kd3utff2Ii6bDnvPk0qPmnjDbP9echelcPM/xSX6iObXuwMfHHbB1/q3RFxCrwz
Z6VtFHDZS+yBIdgbfzDp57elsTXXdsB+l7kVq7XbzaBD+nDy4LIODZcZ5kBucqOi2qSwrb0DCBRe
C+drY2lDaCTLtFpXmppKZjEDnLqNXW6gjVKx15WsbA+DcRxYb1oRk0VncFkrdcLUz0UA48fK+al2
nxkLxEETZ9UpT3e/BC1Hiyo4lRhtBa1J4eqVQqr+9NN4A/pCeu3w/PEzJdE18GARpf2vfloKiiQD
6ddZRxxT4wpoJqalvV0eOFURiQGVtL25A09VJqQso7yELnumfx1RUfWGW/MQQGkMFw3Uhdy3zis5
5Zq8W6y1H7wZgG6S9zSd5Xlj8yorM3A5AopM8SSeoVeUgQ42R84upBhG02wbyGttxId4Lr1GxIj+
WAQMEJFMTWnxiZsFcGhoazN4dg0OKZp9OQghsXKgU1eRW95INa7blwoxT9EAdPSQReJyG8fiDv/Q
HUui5OXOMdaFZX52LbutaIais9FWNrtXJVmtorGAqik9dOGn2+KofmF+3g0Bm4guROetsfIi+uXB
NmCDSBvVoLYGbEhae/qQ0m7trD8kvkFUwfXF7SAPJpEo24q/1SsMPwshaVpGzQ3YaC2c3QJ8LMy2
MYy2eyoQDoOKuZ1J6T1nsWbIoEzZ5Jz9GbUzIROlrHsThqSxHu3myCyqbyhkI4D9Oqi+99/7Qeom
vtZdos80ZJTxAy34qRfwBHl6K90jr/bMh+agBal2DGO69uFYEWA0tmLFPIjsgRabavwHXBsS5Fj1
zP6/OnCtka8QcjRFvoJYgxDV1whoZq/aH2i1Zh044bEFsX73CcLG5lbz77PVyTOK0XdW4XJ4lPaM
ZZryfmCplXxxZtFmg8IQF6gsKL7xRr+D6ntqQaIlkrWZ7G4N9Vu/v0xLVt9c0VGvDhzEmpAL5WaG
zDxEiX9NiqUehgqMi6IACSguAvPb6uppmh9K8Mid4pRVZYSjclWnXxLA6gK8EQA0w7bkAMoEB92M
PuvSwRohtW3VWagL1JVuy5QjJjn+mQ4LWD3EUFlMaz7QU3/GVRC4Ut9/YpnONGsBSPIcB9a9o5Ki
tbaTvzDLrouWB+ex1UI907WheiUEifdKsMcCxihgIw+tSuy8Pur5IjfXjz1RHD9GVK/7ApsLnN40
SosqYwyom7hTCijw24wEfApfPGzzl5oafwiXf/5QOdH9LH3jv2uKB882AK41KMfKuT1mRaf+dxet
AD7OPgTBoBtSMGYtOihWtAHffpiOtfesryi4DZQYNTvab9ci2H4nDZZruPzyjVhg5UAgt2l55dcD
jbxxB1aVlsIEtn/HiWhD8ka6igwzJgTDA/GWjoff6ieWEWBsrWTDBo3ttolvB9Xl1iUqI743AdfV
lG88wO48J1Xzu/NcLrmiuBs/fpkUtBbnkRUDweABEJV3JpAxt+wYcX0TaDUSzq7LVDkRe6Ilb+U6
5zJzaCQZHbshrwVMnNnsyvjeFEKN62IRv0AhdBGuqTyFhN+XTPtU5pvQVgVlhu6XAwJYy0mPeLHw
azkHBo9nimSNPNnevyEEtEv2ezKbmIkcvzohqyyWyHQV68ir6U2W+Aag97BC7yrX1zu4h3OCl7b8
qNTLzHalwEazA/BTsXwE3h+qN+ZCrDHZfd1zX1kMNTKavuxhnhgBaJNNGYwGeCZz4nvtwTSEK9LW
+zmdVe6qqwCVJVFWhT+pblPJ09VM17DgrywcznonBIXnNfseSdMOkjpGGj/NefTZrZeOD16rBIWs
pC0ppybu3fKQWKuGBOa3hIm0pnsAQAEy7PfXBZsgGd2hnG8zFaa4Mpb/xSAhApbekKC4xWNKoXhl
LnYXiRvdG0GZAnYkuJs9u0Loni+xcB0GWqYAJplzhWzaR1ennKIk2MRVgTbiORJCEfcfuaFkKAP1
qA/RxqkuqRk7MseqBB8VbJL6Rg4t69YiIAiDePnNt3VRwgD5g9QE5OztMBk4/bCkYXcDuXooCFJZ
Zsyyo591IWcTugqU2KxqqBszCsuFk7hsoTxHqOT1Z7C0GoSAgx9S3zQ6TUs1mfp0jOD8aXrUCWDB
z0rW5XK7dq35nCWt2fo0Z8wFavN9trNaqoYS268r3WpBogxdXY+xRTMf4TMq9k5V946p7TOKY9w9
Vw3Cd1guDOfHioLd+i9ISOvHDKnJHsRCAtnC7b5Ibrpc3HpzptXZwnhmG1BjUaSKsnHPICR7mYb0
9t4VPPBuMg0O+ajKwIBfNMpF4RFluk2a9VYg9jCxcur9a6n0F/j5aYQMYKPmyfW6DQc7QtemJNmG
SYPOXHSwlveB6zP/7YntOm6ypi1pgC2yqUGU+msivvpZkDCoqkCXeXZargwyr3zTNKvH3leWifKT
SJUhvuOVcWVkklxbv3VN1hq1E0Ejcqi4zRy6/DARKE4JZUCdoD1s8X1gsYPw3xNncJ1+BsUH1XAz
lvqDjXn2tGDoIXrIYCmpQjr/zxE8tt1IXs4ltOikt3lgPLHmmWoVB2wAVn99OEQGOQ0ah6JY4gH2
SeHdNm1hcug6WALGr3oPdLS7x/ofwkGHN4+dNAjhTmGXDKe/uFsFXwwYQZQj/zeM4yQWf5GkcZ6/
gxe3bSM4gsKrEQbwltd71nsv1MUMfUuSdF+DQ3n/jh2xaZd1PRFRXpoWP5lFwcBxtDw3WszwXRsI
SkRgzlycoVuITyJgABKXrkY4FDB3H8LuRj5zz3a8ckWUA2C7Mun9Wps5xYJ+dNxjWwkhFHAT0gz0
3xQ4TGfOqKJmMfgqwm+LsIsoP0VRnF78noCyDJ+Fg+rMNbrso9K/0pmKOxjZ2LOHZMEA+pex/Ccj
ugLG0WPm+nrp9og2DDOCc/FqeSxa6YKbYacl58CMzre9mGiTsg7pGzIi6JAx/1WyBq/ryeVgJpBD
b+2dWn2/wvxNSnF7LGhZhzeE+qY647iI/vT4v0FcP/MsCU/NsqDksG/b2yrWBWsSm8bY+HQyKqwt
FBb5CSObHZXm74hpL8zMpRf/mH8Eyk0WntfYUijg/Ht431YblrRXz1rASOFMdOFFfQUbNxCPCQYX
jHzGOXL46Tc/d+vootmlcBrecbG8L4SoYvqepi9TCWNcLOvBKTYd7WMftgl2n6RsdvExBLFLjdk5
q8V//NGTzlwSbHHHi+NCfB6w0H6Vv0DsldhwgbelHw3i3Oud03sueLEF++dCTc/LoPov9R80Y7bg
Oz+2HSrQbLZvbBRgqV505ajnRdmnvj4C9PG3+goFpzEJY9FuwpH2/8TsZJbUS0DR/I5nq5tL0MQM
9SDIL6rLkbNMdx5Rrehit+hNWmyLqfO418UHHrGoubDDmXc6levNtJVUM/8QuroicwMWYvN2QwX3
65cgD9vF9uI9B45/ZY0LdYT9NsTNk861kaSEFnOg/+doD6jvdEoOQtIauT63CWLGqdZX/K9XFSpM
dCTNYBGJz3/FBCe5khTmmjhYy0IZwoRk+a3/VmmxqvAd5MTT9t7D8jz/z6flnY1tAqdhScffblJ/
zjAIFGK4kf7i9OqYw8cJoSDln0Ew0Br+jkFpw205cA91/+Yok5Z3VFjbJXjeIV5KEk/z6OU4Pak9
cmkXgeNAwt1teZmFb1fzD+nzy2nhJxWTihgicHp9525lxssuJZgqle6djEboLrfeyBHwpus3DQ7C
wru1pGIJoj1qvMvpuveh8ZdjR1yRi7lvC6P718W7i/Nikx8RaDTJZ4w68GiTky9me3R769wxIHhK
+ojv5NvgppZNeIyHYM8DvPbYUZrEXO1V/fFxVq2PKW6MpNIDjCeDu1FSNDO92SaGsSMFMxZxuNbx
HfyhU0Gk6Xt7dLSa2mVDlKZob19jY0DJt4muVN+zLv97vLcvmsGV2Qx6ScGWHNSwCB8NQXT0gdp+
80uyWs7HvQBxfMPYXGw0B084+Q07W129GoLj7QWi5BxJOGTxVTbY/7Zyp9uOV3EXVSkt1wjTZkfI
BJrgm0zVfRq2397Kk+VCoNKBPgZ1T49ue8fCJxO4emuB5TyWf19cv4T9IWq340UbPiSl2QEqYRn8
CngA8R8n63fspTYmh5vdLWzVKmaUkL62zkWjINDsUNm6KZ3ouCgLMt6nLX0Z6xst5xVLbvULMB0P
MzbjOD9lHyC76uqauh///2p9YbJ3RgY5VQ+OQnDwnmuhoHKqCAl4uVMYZYPi0gduiaiIb9Ea6bp/
nQoxMPf7BpFttehWzod56cNadivXN5rdXHpDMuPOeHtqfUozksuQZLOq48GnhdTDUPaPUy4d7JUE
+4kJ5fnjxX7G5dL8B18u3rEVSQxkG30OhLy7rYqwaJUT+2ni8GLacf3++W9AX4hz0qLcwUz7hBg+
4u4FrbS7qwQ9MIwCw0+x2jtHPrVekTAjS1lQDhQuMeQhBBRtw0CYE+l8gko+GygaR3X35zeu/wxO
nw/8ah5a0LZbd4Tuf2WfkIc3aCvcQULgnflfWRqTCgpZ4591U1sRBQysq98jThITU9rnlwQyvPse
FdDvErQ9Jpo5av0FrCBoiCV886SJzV0RNG18L7Ik7zFFrxNqdNU1WvEvqDN3fy5o8+e0Rz8oIcxp
tsS7tpgrF2wSfEO+pWb9XxiOi7K4bnOobt3CAavMKuA+LWZEevC52d/EUFfl5i/pNrVDlEmR1Etq
GTd+z+wC5LzFmIKjLPWaZAi4TfLoQhqfj1whmnOzHEpLsIOkiHAUOU+hXdORBv5yGpGjzYuZABjK
KNx6YgqX1cX2iAhSGzOC4pb960kVhm+4luuwRzdj1LRf9Q6IO5gGsRNFzLx44zg+ADbDS0Our2R3
1z2y0iW2ZV3yMjRh7//nBLH1y7e8zk04kHKBDpYgv6n3vPdA/IzIyCijK0T5v6zYO90LDly/Nvpc
NG3kc7Vkj3ZZy+umkliNNWeEJJl4CuqqOw6Y6aCDSpS3ledINz0DAYh5mUh1roToFAa6FmafXZaI
PAC9e7LzqYKBvRSJN5sHhFEx1/nMFLlGFHrlDu+4q5/HTwWuJz+HZC1mw5zdr2/szGSMDnEZ1UfB
sic2UZZuGR7Aot88OwK88XHss5l4wGtmOxTcKR52TPX6/B4mktiiV0yVPATkGiQSpYu2vzFaylNp
+IveKQJye7UppZdMN61Mbbzx1XVcZEFn16r5UjUA21RPB5rANPpWKj1WhuVi8OnhG6ARiDPGXIKz
ceY1KSXshnOhgHohHknU81eu6jLzzbUBuqF3LKXFjObQtzC15ztVHBA4XVJtMLSNQZxu2nbik0zc
1CrHltIVz33uWEP4TMe9QWB2G095KGgH22jGRCwLOu9c+1eslby0eQycCwQRCszS3ISp/qFlgzxt
eDpYfvoU8octdRz4Cvc3ntJgCjIEdymam3XU+dQbC9eMmDUDxf9P/qvabfLHAsX3hkILeTZz8SIh
8qZU2M0TOq9Rtw1IOwsBliVzk436Am7reqg6qlLM/reyVHMKWfaooTAlUOz0BylD9tYNzGcJS6A2
jpctmzA7lE//huPBqxFeOGJnzOLFA9DzPSpoinY3XHA1kNcluWH8bKNS4zs1YtEB+468tpCucKbJ
UyhBRUDcatNFQyBKBVTc5PyrT8Xb059kIXMn0eddfBxIoJVEo0jYSXm6+KQfgPepJdx1pKGpeGPH
dQ2Yrm0VrSZtXQuHOSwCZN0RbDRqP5ZXHuWh7iuNiKZV7XeL5BpihL6gEbsJKnbCw3cjnFYodrcX
9aXiY/wBxJUc1YVfxMqYHISqVfRQQXJJ9ntF7QBEEMP4tRqL5PVW6irxD6E8ysDxwGKw+yQERXPh
8Wuf9fJVtzoh/Ck+CGPp+CP5KiC0owhGtxHhhJVEBxsuDhGXVIhYoR3JSb9/vekMYUR1FWI++qQf
5gXleQ3oxDyIo1n/tjLqW8t9cs3ulk9ayjepbA3d8+cOOQ84aGkpqdOFUZO9XZTC5Uoqriv9KkX+
2vlhLeclFWEspM2rTT/zWeXK1fT14VE96grkV6H8g2YSmS3jPEdBB0LxjQ94kD61587ZeW+2esT9
qAZq/79ZH1VBVttUaD2N/ho2wmH0JmMFfF5HQcuo5XSUt6HNHVUrjhouXEUeo59cqpMjmEBphbTd
Iwj+iXM2wPtO6Qay9gkutD04YX9DCIKgW9QoSQMYNtIk5Bgoqh6r3OW/Okna2CzWE/bALEI1t+1J
3RLBzD6ftq6cpfIVAPT7y1KO0EhhUaYnitzXPrCX4lDpKJzmlmhAgazBQPDqACZSpMuR7YZSTiyQ
H76BDpNpsrc9goFiVSNYqJkMJegt3nT8HadiOFzTtJGxjl9v5BICR/cXN/7+7qQt5Ci17E4CT9QP
oASzpXfvNa21XgNo/Urs8Hs2mu8eZ6i/2+/0Rzbu7vo3xynYpYyO5XM5zZfnE1nRKqSaFR42vosZ
Pt9yhVIEhLrZaxxVn4Nr4oxRHt1IWpRBmTna1Iam2+5h8PlWyW8KSsB7Q118BeJZn+MDq1KilZfn
fzj/+51nE411N8DiJdEzZd5R5G6Q4CEfKMUx7e1TmKCqQfw5YODU9KwyH+x3xdFBxT0SrgXZPHYq
P7BsjkGnEbwzEQPZu7EY68cBuqSQ/Pw2i5cwDqjxJOGWoPZh6U6NYnQs2cCWq6g/7YPVy5lmFyK4
iCvy65G0E8rA3nTba0/mSGuEAHRyvl4nZ3H4TkwhmZjMy2dGbZpdU8dA7vjZmTv/2POX2omy2mJb
SbziLQ+Vo2l4cf7F0dn4ElppxCnRrTOyjb6PdCAoGxo1vBYR6ixj6hmP9pib3VJU5KX7kUXf6JJ5
rZEHxLxPLnhUHEv/sihNtG6AHg+CxufwI1WWHnfTdVUn+CObc7Os31KnScadr8pVG/KwAYFVuJyF
+3AidkIWNzG0TbzCI4n1xvDGWAHLyqJfCSx74g9vPH5pxn2B3QEMV2kYVMlQrpsoJ3uUZcgA/35P
D5ckS1ZoqWWdvw8ptoGaVJ0BS32rl9s5hM3i5vXjRUa23l93Pp0iICzEO84mdwHAvO4c92EC0SDK
MShuz1RkSx3/OU5Q5FGIKaBv5ASu637bSyY/ZfuqFb6GcUkFvAQfbkc8b5dNVXcKlF/1IY+8jvQ1
PvPdTCtPffyAyfBrlFwsYWMV/m7VLOzKyhVram8GqLrdwPbiPVybydAflBr+JZ5E5xW6lr/dbmCn
SWl8XRMJBFBa6Yv4sxBNIfVsNsz+SZ68iAVD5fDRPNDNShTOrhInf5iw634+08Kwj09CDyRGEj3y
K9yZkTH6ZRpkPMWZCtSLDRbxp/V5cmcoPVtBlpMnKwJfs6JyKJXEAGUKKasDsF3QSjxvZYNu8+D7
BLUDOWHFmCO8b3Pkf5SJK4Y8Mlqo2v66Nu5ykPC44KO1JMSkpZMbZw27P3zkdS5rMmGDepuWr8Q4
J6UnNBMSowx5RO9LXsblrxEq5ntoT+KGEppWAHo5N7QNQ58of9tA9MSzv4NlvTuGJIe21IHt2wu7
xtH54m6Ut9sJH3i4upe1DB1KR3+YC2xhLTg59AoeDC5wkDHkLmy5CSsncOsiQtoy38qvpUwIOvko
pBUGXX1sjEqhK/NV6NfcCjPvcMVOUCZ220u/tyuiApZCirEWGTtuI9ex1IWNm66YJTF6SD0lwW2k
IbJRbssvP2txsBxDXwPNGk/eyNXDUQEdtRWRlZA89zSLcJYv0J+7olRasSA/tF3kP+G0nidaj3IG
A7+WXMhHV/1ES2apQXHnajM/1pHmx3Lnm04P5lF8wFDvXfXVEu5yWCYWy0NOxp4sDU7H/rfJDJKE
+n8jKHciljQ9HSx/gbg0XNKfyQJ/3n0aGk6vdl5lBOCtcTQUKBG3Fo44JI1TAsZwggvKLi8aDF5a
9Q7xb1ezVuZZSZad7QGyvVrdQzQoDbP927ruE31ALMlJ72Prxh4WRkpOhYFKhxscBcrVS9OR+dZ/
knDFb5Wliy8JGZErJUbNy2TGP9wvIMR4TCNy2cs+GtOqGG5cYQ/vu+Is+hE9d/CkRte9R//gG4Ij
7U155NCZhQSs0GqDM6pQOaF1PWrb37u+z0Py3DkGxLx88Jr7R5Yl4g+Jxs1bd4xFcXwGB53jspeZ
GL4dj+W5VNWcXIeA1xpyHHSywV++H7xmiH/xzWlLkZ26Ll3nugxxVId1s5ckEWeTkjXBNTo5gvtR
AlJU4MmZxiYUCoEeFRRRGTG7vg/gbHFGa2cfMvufvmSy/9i1lVPp4RzyjBkKJwbA5cn0pXNck2/D
rA/EJutYcn3LdgGIWPJkZUy0B7YC4/gf4Ea45/QY9ijGLeQ2MCj1yCiiTPl2VbJ6Y2R1icsK47PI
1hc3LqApPYH+wFPk7rAL3dbIe2AcoirpEcbuhuOB8gHCVt6yRDumHbWMHJh2HnPJcZgIjoq9gMFy
qkHB9IlTjlUol+APDy4Zn3Dr+UY1eQaSge0izMlG2PZht3K1eIJpSChMgu8P7oNMuUYyoBD0oeRK
AeOWEbgO79juMOLUXh+mybvlfWnp2jIuxpuhYSpqfxc4qUONCl7zyWkW4L0jZFZD5YUhpCfWEnV5
g+oQZTTuZqFSLJnfECYrc9pIPMAMB8JlUNJAECdf8uiCZ5opIfCxAPHkLOTthNLmc1YwXrMkcles
UGUPG3qIZ4s1HnJHEujd6QdFJ+UIn8BifNS5D3/iAIp89CePKgMGzf/ihItU8xZjPnEmyXMQUomh
08TAPWaT939T7zfE0qKflkyB2g99bQhTvDIL+qYiPd+7J3uDHj8VpiGAmafRpepTyWZ4lfznLJtX
qE/HrwQjP3Yy1LveurkN9oeL3ByWNXad6aRVqM9NFF1YZoeHO0/SuGc9r7GyrWnKTHOzsDz/hCUZ
W7/CJpwNki0odhJ6ipgvTTDE1bqx85xUwL4IpGYN/yaC/iKiRaI5CLuda9T+Conqbb5bH2IAr3yO
NZubokpLUtUz1HTkNWZq7y2JMTaVZfpUUF3N8AWFMf2IJzk2DM7ar3FxHQseCpKyLQyJm5bP2+Y/
kenI1IfeX5OOZlMDIJGTsWBAcluzs2Pug599cVW0ms2IrwU3Brrrrqr3RZ5fkGNRaB35LDtSvHhN
DPJlAXr15AovW82CIr5Oagnl+DfjdrUggqD0XitsvBVbUY3akd18yUtw8+kyQAP7qO6AVi3pTBRr
TvGxjorsi5toQZIFcwyiJPlrj4HfJPKgy4v10f8XoSKs6megU74GbZjal7pYUW/DzjWAZUAnIVZN
SIPtueYjjDmvnFla7bsNNr+xdTw0SYfcYBuG50OOBCSGGYsl10kTiLelfdtU1MJkT/XtMrQfE9zr
sOTHYvhLIJr7HNRJbaTG1L/0na+nHh5TxcP944oB8wJj/cgOBPmFz2U2istyUAfK1ncMtCOiEhPI
OQg2kvB4x9K81tMYpRYS6Qt48695eI8QrbFng8xnPCYWT6FAsaQ2H3c/hCEmR1VkR9IXqMHYGCCP
stf1GREu+9BPHaK3OSqu65LB8JeXhIW/OTW7vZG0BWpoNObP1ffhlwYISx0ZWsZfgWeFV6BU3EoP
Z5rHkYrHdePNBwVvY2k6lQ66Byiq1UhjMKq2Ce8W1FKYlE1sEiOzuE3TDElJE2QdWACCQB5fkw+4
ehlVeBymCuMW5iuf7K6682TeFuELLK/u5w8hAP0dzp44OWcsqfXGcuQuFlQg3Gm8vqcO2fG0KX+4
8YGa5WPBTb0bUd/yvy3pb/DCl3ecyQPR7Zhwc86+uzLHyhCGTzLKZsEdrsVNGal2pXyCyTci2c+Q
1L/Qc9SNYvVngBGjl1sfdoljCPuN0LUB8Ndb1RamREbV8pg8JUIrhOA8ma5J8zfJBbm6YsJ8uxRs
3V6HwTvw4QnMWRO4qBCJOE6b5zVuY6GO8gYW6EiLCM0+cy36zeY9jkjeSqzBTw8kOPwywuCtwqgd
VR3Wcqjk4HWKJuuP9ME2J/A4Hye2kZJ6crbCQbP3U4gp7OadcCQxCm3pmTGE2Wshod5BS6L/CYdf
bpwd2pVaTUF3WenTKj4tdUoqm5KqM6AuXzO9ZU1vCIZPPEHA2fmEXCScc3omKoHDHJN3fwiXpqdO
J+0M9IQtYwCzCvWaH+cd2Jrlj4Zh2jgmqboTYMrBbeyIvEij+zj/zYBLg5tZNYqTwiBetwFm7n1b
+wphdbr8ctzw3Z3gEkvE7ZT0Cag2pf5vVZ5V/BlfxISlBss5FSsS/8vXg8v2Xj1o0Rq4zSubo8P0
RInNY/U9F2XHOUK7CtSE4Egpyyjh5zw/fnkXUTRp6nqI0P5IQG7FG1b65bMxN73trcmQe35x2xbw
zh3ySUmwzvNANhpCh9hWY2NYK/ybksLENQsaXT/LO+DLw84ZMgHXyGPr4/GM80YJiuYL6nCfMvXC
QBipGpaakQeT1PN9CyHG7jnDO0gJafBnutmaThYB6y727PKoVBBglsdLRAbh0Zk8p83SpczS+dHT
+Hjum67WqdgcUSEuJg7l31SW38Otr2Zlr2Dlj4iCiLt5cvYM7HTKIQPxgM1B18Dx36VKy4W7vkvv
iASnQG43hfDCFkdw8C1GuJI97UxgfNz3HV/xo5641AkgL+oSuipy1X/PlwWIqb13Xjt4Hu30Zw3E
QaBiwkNynhQjuGzwz4zkvh5t1fypm9Eq710OiXHhx5wqDV/8tMP8Mdi+VMWWI3wf9py1j7gfCYeR
86b9lQgcF5K2m41V4eJdYM5YYlxbia5+iDlFnymJXvnLeGiuhbbA9A6tHpzLWE8iEfCFIGrDelQ9
Oi0gR7uVsYtxAtLl2Rlr5W3gyebWOKkgZzy69qffQvaUuZgLnQh71Byt91Cx9DHfXuZ+IVntaHrn
02IhJ7mAz5EhbNoU5A7Wd6uV41h7bGlhS7VIto6yjAiQrA43yW+MbwHHsqdUe64eeBL82DuRn63o
LqCxaJTsHtvUGKbTufQlg/+WtQBRtFq84hFUkHs4fIUHzrmzQ5wR4tYlEWdUTXB/wHc/EoxPxUDM
rB5CElPyxvL5V0IJDN4KoujjAhnDgLmbn0IY/FYvm5AF4HSOaG10nBbe6UmxQq64MctDIwkV7sbk
2ayjdPfO2936abtkkkqBJfSMPTYXI3q4QjgPB7HKJesB+pvkjEdGYy0XS2dTP4bQ6aVqN3ItBYVn
Q5D5aVQ+WhS8WjTfvpuPCvun47JkRZm/+bYFMQEuC1Z5w6PvSrA8giVQKRpFW5Nr62FfHqxFSIv5
0So2uvZfvyZMacSHXV8jWPq7aj1Cx9tNmjP4Jm4OOt88EQQv4IHfyNZFd1JLiDgejcCeXavspZkR
Xd6fSwZmDpYp+FEr65OH9LSwwX7KiHJvik0y0OTahVhTmgH2tEo8bN5GLYjsZa0+UozH2+3NfS5Y
+tbUjC/IWokkN3hcAhi19VuR+b1P/qE65Va6u6RqpvY2igkkTHOTV9NMGkbGCePqOBXuCG8hp7dp
wcPxCCukx6W4NlQj8UNBEiQkbsUXbyZCsTQDjLfrBeu4zPS+vwYp5XdTDxz1J7TpZ68thOB9iLsQ
eh2QHCRVXEEZ/cAQhLpttuACBPX0/BoiA9y5uyZxCKA7yE51ocU+8YKjCW/nR6lhXL5Vg/S4uqG/
U7ZZfE7vtL09EWO9bdwfbiVg1208PLbn1SzhAp4xIBowqfOmAgLBdWu/mNhCJZJayLHDx2EpHoJH
vPkI3p1Ii23xF5kZ69KqtgO7ghMvngyLARAOwIGr5YdI9igJ+gd97vZN6ldTUJ4r3HMrlwGEPqwk
Wm+AILcJTd0T6tT2VB0ic+wlXyS7cqB9VPZDq6oQowj9WSrL/pBpIKEDxqhNG0cwWEamUv/QRdut
GWpW8JSaJpe5O+DwY4Y/GyW5qu+RksIKPJzXdCA7OnVAfnKvEdCeae8C5vkY/gXuei0v3Y+y6Zv2
OrjwzD9RBMIhnaqgA+EHM03veUm8D1S/YEqhy8Sq1J/M9+JPKupwVmyee8FGLvv+L5Ou/Zp9wvD7
O3FVuhUN6KGEdMJet/DLZyHircwFr3vxZQt8RkQj6rkhAxv8eszKN0EZ8Ddb2GmR9y+bLSlr4JE7
jGFUWn/33tOIH/NHpGVXRAGOU8Vlycqy88WrjkaOTmO8iXyD0lMxw80tuF/TgGzdipKfRUTayaRT
OEaYQnL8cTNmbLDGjEodGu2hXqMMVSowJ016RDss4NBVlOtEWu9tBVs6Rw9Tx2+rawSNQaig28RL
nW0faDt+vBFMupRfXJGJcuKvhJPbwk4AeBxT2If3qjkgxviy+6htyV4RLlfr4u11fR/AThOFBjPs
pcznwfqM/QoMHaklKH0fMNHKtH57L9BzF47hcYHyZ99jY0Y9/m1yRf3n2oeqspj36CypH/rkrYlY
EShl0Lyi2y4px0H1P0zODzLdaxrB1yEw4kdHCVvoOnr12WUeaHL3FBarp/+unBNzVG7z5goc6XKy
YdFn/aybX3hQEJwTW7xhpXjnL0FNin39zy1orH34NpLDX1wEuitZrVjkUSP8xDHyz/qMsvwopOHS
1GVHEL9fS5ufytcInFE3sAaQ6muLGWe5qZeSWhYgFEIo9QyjvbRScdpc692xY+jWBlcCqhrcAL5m
SNcKKMbDQDyob+FQCeWEF+eLkkWYkz2dqfgNxElNAw+5uOU7HHJJbnnf+jpWWuJjIwEVhu0UkTcH
1bw++2ppzwyGqXW6DT/JcOuC4o8YLyWiSaQDDffKAuzguI8YiBwUbAQK3RJ1+R5Lp+qvq7EiSZTo
JALNSUynnwLf8hSDj0rnohHiw0IPzK8Wixh6c7jqj5RW1oiR0Wv5i7DflmpRrMLtcYnTzrNORUyq
Vqj5+ijId+rq1Wl9Fd3/iGetdk+bgiCOmV5nR6uJGHqmKWGjmj5cWsuf1xwZl/R1rts2jJxgt5tt
/e8Zr5c5YUVKRjayDg+2V9yTRNhncuTQlhO4dzoG9gvuKNybd2GPrnvvr5IXK+18UNHj8c8Sgut9
F0yQJRJwia1iOMqTaSq27nouXHZFAXxlhW0MMuByGfpDO4C+KRggR8eslAwwzxdPc3z00iMaIDAP
AygrIvIsriQgYDzgnLnq0rpasBFt6PqRT+h7bM5G33R6/wXGc5qZHUw6OliowYQtdCANGw5s9g8c
NLLNJiBNulErG0P2XA/lKl8HqFdh6XwAfwNSWARgxdvhvvmMj0qHlih/4g1bYiRKb6da7qwnvwjr
6H4lqitLAeHji2IZqJyKO67BV9Dv8puC5aenP687OGC1rrTzhaoXKiHY9CPEABT9k3zo6jQ9yMTG
0Bmatlp8F0n+w7Wt+UMaRdokNbdBFCDh0gQ0qOKW/Ah5QrV1xa/gkCyXOr7b4Q8Y5r6RK6bhHrJ8
Eejy8R4r+E6gGmLgstbB0Jvmg5w4Z+PWt+hwtL/F/GenbJbEpfAxPvjIDHNNGxQc+jG0oMhzNVBl
dhWUSWqzbxb2CCj/7lE0da2PzG0xotPE8NstOcZiPpW1ywdrKkiDU75HyzR1xJ8KZY+eSM9c5jrH
u9+aKcxaPYc8P+e4QYERYpRoLc5QgRR80LPdP19unVDWGbICLWozuMMgOWVitO8ZPwQLQGpFd5jy
Nd3m3BaBKw9jstbfZ7YvmzSpaOIzO47SPvgFrDWOSsDOWW5O6RrRISzReUQ2579f4QUTQRaxeIST
Q8B+J5G90eXeaQrjGWK+y2Ue3A3Ic0NgzMC7Ip7znACuKI6dEJVvUJ/Ecr792cqrusoElVTxVp/M
FB7a+zLv4BYx736wdZwgWmtfFXRxEiOnMu77OMILzpI9DtSYdGq11zjyQ/QuAGic1cUg04IWN/IW
pu3MDqrSzb3fHsPWcFNDrIjbeRMajBxi+/WXqNgThITSFRe6KlLvU1Jtpyv9EGHQhEztMj+x1zhl
uA07wsHtqqMQsu0yB2favLk83wqHVmVwATFdcIKPwoJhCEBlh09Rv1WQAjn6sYahz9kpXVBEA8gJ
FWsp+Hj0nuoq6JcYsodhFJT7+kSA3MGUVZTvdIWNc0/2UeDJPd7Jz/NXxYxdbq962TOYfiwUXe7y
e4hNB7IVxhE9A98Hn3/mYxlcTjbVzp+olzoFHUPyvYiP9FeX33hQRdqVW6qqJO98BKVSOBUjdA2u
qUFw9sME6RliQt+fO/yZUj5D3RtchdY2pxlTRi16t6SBeklvbfZqODUhZzJrB1nN9aEPXXktjYQa
fPUwAaDGdCznqLqlVym0GE8WkwNBA4t/008VxRbD2d117jXltPtQWcUCqHMRPCtu9k6v472q3NTp
jublxxerF7kklzf8ixuAEz5J6neYqd1LFQ4r8dlW7GsqChHB8F6+J5jW4PKhmV4i/HH4KPEdrkFu
gqr8CvMFmK5b1bv22b4uh580MfeUpEUcto1NuZpzQOG5gbjl6Q/tambecxBFUYmbg1g3abJMkhXH
ZIPFrbQS6lhDx1xYw/HROtpPJww7tXu9GKzbRQJo6dNpOxoKrJ/3ToT04vcNWA918eeOt8TM/4lo
cFQ2Y99g9ybkyhSYFPdnewpOdXfnriHdZ5YflYfWZPNxn/64D1eiXH2DZyRT1I2h/0ugXemzUPvS
ksuwAbTS81tBfShct2S+tiwrmJ/TkFE6+n5A/feeOSg/zh1xVezfUaUHch+eqZvNBv7ztUIwwwXQ
P6HZHRdw+X+lqFAzexL/jUPcDeV7x1zpqwryDTDgEG+DFy+9orOTAQoh4vDFRL0YiZFzwQcDrynp
FIHbOoK03cmFCFmvUA9dlVrvfH559AVA+o+4xRvRy0cfXk7Yn/V+Izh/LcNAgmw0zlkkUqjohu+F
HbHlVltKljEl9ELHVuPoUX8rMEePOfITSylkw3zDZ4LBqAjcw+UnSyZ59Dob6aKRAaTX+zlc9i7w
BA/QGiwBgCZsgt7uqNvgsW5VhV5fzCOXStgIp7Gi6ejpTK2UFIh5olRjFD0BFmet9SwafbYvpd/Q
1Qz0epnWLNschRl9Mbxa2S3MHAUeD+XtSk4hUt+wa2EJyoA67inFrRQzxQ6+JdnNy34QVWH/T9tu
sWyz+y5YUfuigMo1H2ZysfCALOyPGtnaUV/BRGhPE8Jy8ZxV+pskjtF+5cFkeCUeYoZOrTgRFQii
372ajrVZLkvSRkX2V5pwZppHvv48c5ZkWCHS1MwNtgSErSvsyOTTzpY7RYczo/hHYJ84a/VKriqO
72DJ+hcCCLJNGd97R5Coa+3Cijn+5xVgfyL8LdDk+HQdcAVTiXktmzU4yddGO1teDJig1vkfUohT
6Dwe4swWezupNcGRJA4DZVeVaf31M70Z7o/34mnjMoepkaBDCk7F8Ts6GX1dHt2YvBJh3t/alAu+
Q0k4Mxbcsmqs5QDWWea3a14497QHN01KWwZhCszR7bGNI4Z/u+ym85tE5sJkz/pRINwuPA61XVR+
3ytbmpPm28OYO+RPu9Lv7rINb4Is6Z2PYbU8dM1I69ySMvyg4XAmqWXO1d1DUPlF43IGe9paEYfp
U/OTagZsRho5C896CXzWCS+PKOVajHSd+MAD6hlfak+nQk0c0mRrXdL33e2JVY5MmWBxvyrAsOTY
Ii+9h9NbS+yu0APos1GIlIXcw/GWjEHkwmz1YKuXf/4NLTAf/tnyw63VNJCp/TIGrehmfREh1gmU
zwbL+6rCs8Aj1AUucFsGoBEdo0vllCYWDGiqbLHCq/YXwNIflCs71OpXPo3WstOXz+EmIGDkJY5S
0hzfSKWfZY77+2Y2BY2JjRrlbAIWpdBFa73xHLYS6wqAROBJhZzkrMGMEY1o9o2MLgR3QVkyoAjp
UfXinxZ1HRx8pRPPOqxHhLF+x0TB1tGAHNrnajsuVkGsh34ks8+p8U9uHqs20dqEnKaehlFDvhEy
qHBPpiEYTO98BuAphq2n6kk6sawGDnm68KuAaGzsIYsdH0gc1KN41UXANVWcJhWm4+2wW73DXv59
UN+EP71J8GjlOMK2legvu33IYT8K2G7iOKTE5q4o9ETPC9zFDFzO+0NQH9VcKwu9BKvrLSwnYlG9
UjjXjZsYw3D4nRdRRaXiBfUPTs/eRbkJQAdZM4h0rPUkXs5JQhF5477dxgYX2URu8ah+MEKpibPc
4Ip+mVLXbgZuKW4+RAMwsT0kRCGxUucyLeCg3cIWC6mdhOX9XtjuF55v9/UFXhocjVA9XxSb1tLJ
+T0QxtbCyIV3D5eNI0PJL/T5AKLe6bi6yCtoD+QjUVY+sWH+DvbgKylU3gUAnYYflowgCpbs5Xjg
uymLM7T0jYRFvKFW57rjoQVcBA2X/8sD2bVrs17bG3RwwzhDzu/xnvy0CukVmLP1Zwm2p+g7Jyiu
2nyU9TX3O1FGGArXFjmx86IONHnuoO8ZOTwHhSOqEBY7gu+naRuBNmPoosec/DFTmY7CvucBPEPm
z7/UASUNQeiUhYN90Q9WD/DTXTbflWrUdXy7pydgqD6JySe8JE2ScGu26wUIDel6zUR2ARfaY8MV
GqXNr5vbEmusUkqh6JQy3Ir4ck9SyVuAQcghr9iqDw+mqj+Gq0234fdXNUvWksXbC+xMx4eDEB4v
VugHXaj8wJygnhiQemImIZM2JmpLjEAJxoQJJB3E5xj1XYymfYQVi1vWluszZo+viXqsvPxUXJwQ
zGy6mqyDODouVvwTxLJqlIdFPPIJN+rC7lErV1iCEYadL+s44ovy0R+rgwOviZaj3Xwe+gMacEEb
9puLcQfofOe1QabFnoW4G/W9eO6yzFzF5D2tYetCJVqBtu32j8F+M+cRKN+T+PjbvUEQJW7cQ0Q7
KYXMVrcRyVSDa0DgS72lrW3xD/OaVjNl0oiCu6ftWCBOEtA3IYjVBnUfXYQb1mSn5VBYuaj3CRTz
TyjlV7Cq2GE1Y6O+yZfmn62hTKhBmk3zcpORylB+bAiNmKQHyZz20TzBMzk7Xbubh7OHlipcbzIn
+InAq5xxJNtA1infLoMgD9p9ikccJA0bcRQjs12vjmbaYHZSpEwvLypz+H14iZoBwI1fuJQrhC9l
Z2ymZh6sCVMIlaGg+FLMhnC6+ZfJ4rVFQiTrlER1DX1QIkbgzgd2EfAZcUp4jLUMblVkwDx3lD6h
LnW6MoXwzxSZxrntG4XJXMzr2k6l6Tcwyjtr9+M7n0WJWIqhVINgpH18iSOjRCzuD5QZnUEVGwVI
zf1emEswbsrxgRqT2Isw7KgFBWiKLckd6eCYCwhXJNYIdvAzIzrCy7WiOB/CLEVM/p80cJl53hhu
NOj24oQF263uVzahqTpIv3oJKK64NtJQoSJx0jNMJSwedNhNomGV7OQ1zIWsbme5p/zrOZBC5El3
wgJ4CNYlN+APx+BuveCODZ3sHABi7thahDsu5u6PG9F/TjhYdp/GmCF8sSIWNK6O64Htwt3BJE9e
jHTmWquIDroUtT8u8tcDrEeREhlTV1lIlE/X9G6k/YRDwEK0cl914fCLuYK++Zo7PTdVuzwK4LCT
uz0Sb1+h3SKcBRdXEaJJC31nWTL9gr7woTKw2abisZaou3UYNbBtp/A9dJh3IMJtF5lZWRmERlme
s13vAsBGVnRtjE3o9C9RIX9Iw/Dq+ob/FnshHmCEdK8C7pYf5wmkHbwZfmaM/lsmi8Q3HzNuK4lx
IKiOE2RF5l4kX4n9w/nSvDM5r5AJZ6syWyD6qZivw8i9LHaT4EbHBnBTS1dG+bJQYR/2VrOMxPVe
2AF9X7dwRYVWH69TdybTzFwpd63gJfTC25siLfNCKlIyIXFC99h5CNbSChdyGKQ8RX/B1SGTLq6J
bBReIEb5mCU70I3jxCmCaTWTl3WXFMkAxxzf1TyDfplFCCw9U+o+R3ec3R3Ip38VufkvZZc1Qy2f
l0p9W7jCvjVJSk761w8wazAwAsu/PCknAKBd44unnN3M7XU7iVMznByoHcnTAzvHL89FgYRuDG35
IdPra5A77JJ+3q1AKXiUBEhoa3mRxwAYDHD+dBCi6IKYIXNWy2c6gSwUHP7oQDr0FXDc4tg68J+T
+zk3rx49IQFJai2RRY5QzcDS8ur+vT/FlFa1+jD2WBnqTi8UPZrbEidyyno69BcitL47K3I5NUVA
89sktJUQnBQB5ZD+bs+sA2JyLg+tlR5NKZydPRweLQPAiuGlB66uaLJFKx1cez3mhb69/GqBXMl3
BHIgTtSO+hyf0eWAcDp3j7SzeZSX0NMsGtW2YxhnipFGGPjtEmC6Xc+kuW27ITpvgDwj9eHV0f0/
4+xOHNhsBsfZ6CQkGVA8uLsfpTDpRWdHUyAf32fole2v/UX8g3kLtNaYC3hoi8MaNJe000WwvgF+
QfcI/nK1X9brj7q4KrwPUGMGz9Wjz2jTYxlcz8iWQ1OAhmKYDU1PQgYdTz+QOpC/PmMve2Xh275M
YLl/2j+ObGsPF72VAqhEq9R6n39J+D8cXJvOOq117eHgHkLjM9Nv7jDfC65hOtqIDmaPumvGocVq
nqpAWdLI990L/8SHAbS3CUzCD2EszWgUgpqJwKySqT+CaTilgxQaTDtzBaSYMAgLYud7G9ktToCr
umkC/cEpnK2D8HHjTwnhSdBwnBH2v+iy5LkUaIeMzDVpwMOzzDDd8TwX/OQKYGDV3/OBY7TlrZO7
v3lMZcRqRlASLmWMpau6mjmeZ819TzPaiQ/SF9/PyOQ+dzH58XVR7yAF/mFDlf9bQVduzhqK2aIW
n1nxaUMIqDHLkx6FSoOKhSUONK15ziWzn7HQW0mtD7OCQofKGKAC/2sqDFw9IMfjGnjOGM90hMOI
jUT9ySLOOzNSiSOiZs+NoDiipUtiMZ3UekcBBB1/2DtdEnrC60QN71Q0Dk+YBYDHp29xfMcxrILn
Go43fk9YwJWeYLiejYD7nOCl/nTrm/HdMyZAVdYDveYBedtaBAIN8YHRBD9bgc+Z8SHIa6zhl+jO
jPkTMPELmdDy+UxrEpWqXIoVPUlzeQUebHV5mgff3WMc8szMIpq6UyYMvUFHwli9L6/QFwrIuonb
4hkKTVzeV9P3JfGFirUKxrJFICieZZaif50CBwfo33Kmj6c8PBRDT469Ys5sDG3eprCG2jVl3fHt
S9dGU8rPmcpY3DcPkXbzLs+TMM8JJhYaurts48KxpPYashh+T11+nRI0j1NYOVLMiOCCxBQI32mx
NeMeADIawvJ/KhI6k+WqXVbVIQeWIlB70dAKv7Y+9M4e1PHMiihDegfI/N46kyNbO6Jn9i4QEJoF
+jdXwsWToKT63cjk/IjeyDnQGlp+NypqrdGVe/gXLxV6LTfQuRsxOe8eoyBz6wfCx0uAiBYjcGOl
pbWYHJcmwrXvalUN5y72RobM3uO5EgxSrU7yDXLEWh1E4LiBOOt67DVN7tWWjwnDSj0jQGIa8h39
pwG2ThEa0L9u/iFKB/kBFoYbj1L37WJAYVMEhjcnDI2h2LP/V6rri8pYkDQab1w0WYV5/8t2zzX5
mn2yptWdvv7HE94t/L6N2ekHY6ohKLYcihr231x3yJQ+TzNQy/xMY5MpUqgEjj/aHN/Q1pxy/nZJ
U2bQdmqLiqtHMwSkGAOTpLYUYolIXbAbT4yjSTfNeTqZRHY4KQR7JApUAMUMgSTBdCJi2MAEBXJE
eQjFUNVTFsnclZdLKOOtqBOPe5AK8l4G/w6ynQM4hcB7O3gjccF+BgxJW0DXQkb1HFk9FhYriYnC
sUp+tYDtZDGIDF2po3wVfLa7WX+XQUIymU/c+j5AlP7L5SxcrezKViCn2HuDRjHh9cnQCSP6ihxR
9rDdz3+1nZ8mwolIp5t5p1iGt32aXbdLSJUMVTz+YJ/gU7SBpFRN7jI+P/E+AiCDnT7dfY7czE7S
TTr+ljgaIBtU1BPrQ3b/QM5ijq8820LBGxwVBssVYZ9ZJBXFU4cia6QwauWLAu3hxFlU+HyKHrkP
mSZPlaGjlhFJbtftUyaf6vHPvkMoeJQT9KRZDo7MHoUagYTULaH1JsZpPeNCiei62jrWuvSPr8LL
PUZHEqSQNxS9CLMDPEp9w2cI9omlC1Ap1MyY4yPrzRucY7joJv8oQCDD1hHP9YXJQS3iEJhYb10v
qU6EZx5OJZDagmbf4wSmM5H7ZeMw+zyliWi2+TVJTGOk2OmkWlUZLQdb6u2TnsKuWtr//UyTQqB6
GPcjFW6PNSFzt7hS3Utk+aa4HVz9Zt+3lgyC4eSinNSRDFi/T9Q8aoW+umdYjNXKrI8lPXQSgwbY
xPIbMMNZm7+YyUIE3AcedRpwivI4Aopbuj27dYgGl8xVt3SlPPIbG8g9BbgAwWmdjD4mqB89Mk8W
uv5vPlNiZfUeV1F9xONrHjKFvSeQnyBpyOo0GeNmpkfPo+xTm1kbtkbH5bVDTbm/t9vvXN52zriJ
Q005JX6CT1Q1w+KcTqte5kgvGqjbbGSXg01a1+swlIsfQwTrttOa2SOHnsXqHA0O2KO5x/BAHS5m
ZCyxcsI5jA0Ab8nrWrCtVLwvzLOvaxPLJn6IgUyTcrMP1ycUYg1S9M0PMwvtcC57yrH4SgKDy43y
GG5AXI1VyMaC1tCbSL8AT+hrPLDYTMVHsrWlPcopEnmEAIChRnf92SFahfnBDSko3SY9vlgnEQc0
ktJIG0N0G4HzUJDRsEU7NuV9G2NnhVnVipeQtSidPbjtTCfmMotSFgAn0NCB5y/XFVjTNXOr7r8K
3xG5FH6HRnsLfLWqTAZ1o9IerXZIycz3XzGonFi1HRsjyq+4oytZn2RAQX25x5Um3hI4Kbf7GMTs
q+1rbFOfurRqxAaJxrBGzRK5wStSy6RlPKWZe7aOdxqiqsqf87tM16f1zig6AUvTxVoi1Bu8yVVB
LWyKeeiygrsv0ldFhWDEnOFy+wHTrOZ/jEB/TWs7id3uR06RZ1dyuJIWSo3SD0iwHEZRpLDS0Lgz
R0l0LWJxBi1Vr/ifpwO+WZxdoluy2pdwo93a8DDvOiaqVnZ9Sqy3x/VKC8PGxLLPJP/3Q9XY3EIu
X78mew+3ltschhqdzeIIC9iFswUxmRFmWqIwkbnjut6pdFr4btVZJODAA0S8i/3wdjbpPkjgSWs0
OmyQi9uIKNA1JBAs9Bduk5oM8lij93woMPOFS8KuvuMKvwOPeFRiiQkuHURhI6nYMWezUrB+JUzz
j76amx8sebItghYH7jOLBfbhiVaNqoxuP5qJpAbaHl0yqghED9sJROwmFIE7c7smYG2020Fu/MBI
WQb8IBXrsS6gz4aev7Ef4lHH0L91UFNawGiGpdztIncBeKG0u1U1qqt/8CI5N99ZvYzx84O1mFbW
EJSnuMCISoouYFchJcYlxnXwD/ioja3E4uebGxLSNa68fM1dan/FWNFYly+zW2rKsRVniUCdD5ox
XCs9r8wffWjXK8SfoKMU0D40hpJl85TpxgHXdQRfw/LgKbZKD/1srGUfC3FfJuykvxc87UybiYqp
yVVxbY7Fqh9Nq40y76Sibgg/+h5VUS1xULh5TK5CNfeMVd9E7jpsBlt9GRjUSkYDnGCiptDIjG/Q
Tj9iqexlFHNMygNZZ7jXaSewCKpmiNJuWT0EsxtzsTRGCQjK64Rz2b8nEhLZ7iLpd3A9JPZwPb0T
2MzYi7nQZol4JdMZq7a3XoiAnSt/82J8HPUMY7Ycr12QTKSI3yewyj/K2QnIQSvz4u60DFfKrZSV
KwYR4cdKYRfSyCbT1D0HpJSEs1qSGc3iEm6QgYBd7RLXMfzcbbat2DVnnRd1UMuYhoCpOZomfX+c
Hxg6qcgiQRvsKH4BpMH4cxBzdxfQm9+YNkBHu90JBoe6yZGgEzfZUAK7KX0/xmNwhPCVtkacFeZr
iK9Mi2KM/Wc8BMFJm8BtNNWhdbY5N57KFG5Sjjp7edx3nYO3NujxqQFuhYrxcO/TycI5Efmgcaok
Omws1dn811H83z9YvxbuwTnP0HAfwTs+gB9jiJka3mhlRS1rhYFc28o1ZgDO2gBEpDgmUmVtBfua
yarKpYrF7TLyj9343a5hd55bOsT+SndjTz1dH1NgUdp398o+avttY/Hh2Ck5ZP89WGJyecEXXa/s
VUG2MPiq4vL5+gdWUlFyiciXK3hlkoOV7iSy+5/EX/CwC0if7kT1oAOcLi1p7fCiYq9rZcSkMmyI
jSBwweLtpUGWVEMG9H12tthVSFBNAo7C6PNCOXMZTTa39vXwbvcL/CRe+tsjTxmOr6SsmmoVfHUP
GWaB7cybol/WOE/zjc+Y9uDGdSFg58vDS6B4QQSoWQU6a6VuWgQa8VTICFPaAXE56rerwBYx8n2W
LwT9IMVqx2XSL5QC9GKkWdlzXTUmTW/tULTAM2hbAYISUNxavJqzOSl85KfbX8PADd+pXXEZJztl
UqR8m1DPgOLEXOqjGn21qJ5/ST+zNNSlV+kH4wPlXRSUAnD6DhoCOHi9UX3rDRRi+YpT9KeLF/GK
IIt8q9REFMvKr8sxRjR57xD+4qfxDKHJ13Gl1IYk+RjsMiLeeu2A6hDWu9Hos6vl3r2bevUHA/kZ
qQyqD2iIh5JaztgQejRDuOngQ5EcmergJzy6uKEkK1VE6JQMZo+ajgOwd4zLyhwGKVXp3eK6kYTa
T/FhFmozBg8oqdWagxTuzGFjWb03oUTuGAAnFLNLZDObr9PypCySmyi7ZWVwNLX8TFFO3o/O0tZT
EDQ8/vNAW6by8JrvXXb8PvI/jYXmxugPKlpAuq8xocMGB+wJsXWRyaeXxgMbNslq3auCLt8jLxbI
dn8zsX7A7V7Y8a6/S4yGEnhlmVZl7S329rHckZhHfAZvuKEXu8/Lz+hYzkAoOwff5TwbP+BOkfZl
PbYRQySR72WufG7QnLOmkQkpIHq7wcYl0uYkhoUIf+cYv75bP6sHeDyVqNgFEON6Z6SRZWaD8heD
1gQB3YxfsaZAYerlt0DKc1y3pvHp2IxjFwGZBVlXAunC78JJXKr49Qkpc/Re13JDUdxKJy/sSKZh
4eUs65XV2L2+hcz6SsNK7vx7pWY8VYPHIlUM2bM71v5DjP38UWSMYLn+elD6BtBtSFof8ZoQdFc0
YXffW3wXz4Nvgnfq4T3urXLH+x5Twwnh33K6dKxFNaMseIGkjv75aepmgm1eTn9YygXwF+9YEXW6
TidM4xU88u5VfVTzqFBC9kjwrFBW3ZBY8IUXnE7q36JzniNfSXeaCQxSQX6G9FrPuBw/WfRJAUi6
rfp8GEvpdo6fDZWrKUDppTWNDuI9+iak6lhg4Qcg9EZP5jUhU9oRJhWhcfUhwSCHPF2FPk2Kj4kf
3LvFrI2CB4P4JzvgeZLp3w3dTtAsuH9tlDQO7emVl6LdTkjuZ7w1hvu3adXA4L8uVJ+rE9xFmx2j
iCqGYnOVjKVgS9y+q6icHj7wOEQZMRH1jwvwiSL0odytHmNhvbhPpcCStRRokHGV2td3x0xrb8xY
Ah5kLMVQ9IzVtTE609ATvH8JQYLoz0srVYXGoyb9G7QBsYcgkaEdAL2ZApq5VzoI0Cb4hSLKq+IX
YWMc+yO0TpTuveG7UbkFdS1kD8xRNAm1sbZ+xye490h9rkBcmYB6uyX3tWpOSDUZZdNLmDSdpvRC
f7M2zkNRATJw0/eRziSQm+mNgzt2nleAaCGSAYEImkv3vGs1n09i+U1J/XVRXpWRTv3ZdWakwjAE
VnGyPrwCR1fWV+hsJV7bUwMFSEFm8ZHyy20ZwqOfWIDYBPY8T3uEvgyJbPH2Wx0giym++5lAOMfo
TYO9YCrzp4i7OIAuJLnXDl57jM84bQe3/n6qgAV6qTy4sUrjSaqMigEEVwzo3CHM08cHWoKlLX2j
j5OKAd9aGFgvQO9BJBSQVHhPsm+nZofNps2ga+JgpYMNm3FkyO48evYxlLv8U2BpD1m9fXvbhQO1
jkeXWJlL7a6yVNGzvnV/CcaTDiPmhaawoUmmCpTqdxTfT/sb2jrMALlUYSHVS3Cn7Y3SYU32RE1V
XYpOp3WCcmbv9YcDxpM92iYdYYxLAoozuMlzYhpoUvwyLI7zaS4aShEvrlx2BlBNKXZElT1hhzUW
yz0gw6dYfw5WLLKizJySP9nd8FTTe2iGH4brSGaujDPPpzq2KbAHdJ5nwcf9fz+LMKcrKgkVMKyK
4qrHJXvhiUkTAuhu0YVgCXjo+tfmF1Mu8RfM/UCWfjLd/DuzyfuTsvA1HWWpDW3vxQU4SpGrIWWv
WfAemDxX7xnxXNgQpL6nRvtPvNJi2bdPOS8g7iyMDZmNid60/xWoRZ/P7KQcYiZVYtu+ndHTUQbc
9OCJvQ8GqnqD0da+vzLrnUew0ogsTkLKbjNiN/Juz/NRnb0K+aj5TynaBVHIl3csQ3klHLa6HFos
/GjPwmjLTVoLwH/1wVmg29xLa95zI67d/9hvKNiiSDOgMukwjC8DRs4vy7Km2j33pAVYsSNK3qgG
/F91yWM1vyddTOE2H8col0qcKExFGA0wM7YqGC8IPteExXvvicbUCHyB/Eq5Dq9z6zWo8J5K0IPZ
fjW7JNjRF5kZ+wdRLq/c3IfISw+r6F1CaXU+nBlpZhHaeVjg5JffPkxot3TS9m/k3kP1Ie39nuTE
gz5M17fHie3avwRSV7PPa5k78RNwbFr3WeMp+OyS4FvDl6Aimm9elMbkFnACjTO45ITndUuO5o8A
6dVgINAIgb8t21dqj899eCGBggHPXS5MIJCxEf8Ha/HfvQyflI8J8svKoeGxkYW2x3TuRp5lzvsM
ul8t6EFKI/L3L+xGZL4ZTGUCSwxWItiZ1+D0fyl0DHZkdC4kpKUq4xfSfyooSOK2YwPstqTd23vq
1C55Ncyp2qj3oE748Qs2/T4uOwV7y8OjcenxcXO7HLyeocPCK2MPDzU7ghSjEEVPHLM0A6LoqJsG
b8Y6//PS4nHC5ZVh0Hq/VKwXcuGFJVhVmKue69T+Bj3Xxl4J+m33Ccnbz1Q0f8zjolEUGPMTswZ2
j1SfxAfWm+EZ+mcIDC8jTu/tISaoFFUCd2Q+K7kblpdRdc1zNSwPPWWjyp+7vJokWnFkNodyLpKf
2PAXGLpeXeTAvZ/EJpbjNYEcci7J35Cg1Uz7S+JyVoXh3t6WB4GgwwBpQjjuOn0qPR2q0jsenzBU
ZpbTVYhSfAXMpo6uzm/0xKn8f4fNKmhhjq3iWJdumcvjaIuf1tbEBu5sRpvDEOaprxsa8OhpGYxc
yI5ZSlLC8/DEi04OYj8SpWmBzlJH95tAMOYZcMro16cVvm3ZrFxK+Ib1Zgu9rwGngqG7f9O4CQcD
Gj/DBpXi1epBvOjq3xLVFWQxdKbAuoInZb7vI0zneE456m9bT55BVi+r2voLSO5yB0IPJ8Ee376i
eQER71Eq8CwvchBzeUC9oHaOHHdq9xR94WVZwz7qVEhYALEQBHfz/65wZYVo7zUlZWu2vYVAqKT7
0zqu11oyj5Bx7iussLzuoyDh0U4ymsHCGrvTGz7RGou4GBCIjzqfIL1WZUPW2rcL5Lk7fvJjc9t6
5hgnhpg37FtqqeaXBEngxZxYTFzDiprXJe4V1iLCKQevdFKA7XJqyGFiDZZjH3DWL9rmEa8XG5lW
d7T6qt99W/MTKO8+SHZB2vO5w+TfRSNtWNWuYRSgJauvTTDssmZjGGebJO2MzbDm+csLEk011Sx8
jf+sG2Gx6w/OlOnCP/ajQAQ3UmLdsJThB0jSvXMEYKnrVbJrP3sTHkOe5oyUjkOoZ5R6+id+frTL
Szwe9jSzy8J6G3KP7OV8gDby10b1pxogNAfF7yf3+mS2tzjrMPMzODhsI2HYevqfcDDKh1mRCPJC
xlmuGbRCReLbzlzjAz/DrzKUldooRntEDK68vQadIC2YDtK4hBwwexdpEfhH+WB2E6CmARjoZEQA
VGxlqb4xiPdkBgPKqltUrkVtKhyhJcZmlYTFeBbukgWVgpIcJM3v1Eu/SU4HGUiQ1mIVgi8OQgwT
7O5+0JZDyzE41NuyLkfEEmsOSbS/PkSz7/kckmVMCU08df2+Jqy7TOpnw9cjWwiDAu9UKgDNDIxl
CSEnDAMPUCY6SOW6O2C01wVd4ohBWmezEB+xq5CLrnMjs9VAPL90kkiZCLXoLRdCA0wAX1li+G+L
qhXLO2QL1Ewgl9x8S6ayBF46+CE6bzyhTw1Hp4+IkO/9ht+jvXdPhcqc8lbNv/1qs3ZrS5cf1CAl
V521Psf0oqqXI49/3/Ho9oqFKUTlRJCEZwPERLnZmVeNA3vtbFbYNoj5zrNpOMxVM8on5lIHxNgm
70gysYyeQQ04QJ+PfQ2zXVJ0VFJhJeBSZxJN9e3ExNtz9fi4lNiYKCXFfUd5jvwkrsrsxArPSKYW
lo6c52mg4hqqCkr9UHE70Syh+55dTzNVT2rY+Hp/SvPDl1A5Ze9obzemqOtLse3OK38/Aq3FcdG3
d543CiPlgJ7MuKpD5APfRP+hMzno+d7OGOr3NdpJIk02nN5aIVz6wkxwAI1UPdz2IHqpCTJxDIrB
TykzJxSBWdd3GMUezBEjqxxWZOQsoT32+Eyfr0F/k0+3T+DDS5xKo4w3swauzAJPj+0FcS16b73v
/zoBzkB0WRpT4oA0sCe68Wa90msR2Tzd7tOcH7ooItD/NvnY5RrsunR3xkx1HYh34/tygJO4ZB4Z
elrliVaJYgKXTQ5VJLV9Uz9j3ENEPVh/WW/OK5IO3rt4gWH3xSZ5aRJcggyIVajMf8wRFIkvziPk
CWFOf01+jrp+lHs1YDs35W7Hoj9f7TzNHNIsjyWUMs9Uax/yrzpW+gdbjP6hbQSSa+Dc1YBalPPC
SPKiidpKpNZ4QC5xtIaihhS1wwI1vEmY9W5N818+PNn2FMoSqxB1pTW49wiLdlOM8qhSQgpelS1E
jW8d+6h9lufZTSt9IwrqqNh2sj2+D2UPTESIsF2hlzK18r4nwgdd2nBctAStb9m079sfCPCeqh4C
fbrTsRzI7xwP7oIVKd+ZqGXqb0K1Jwb+RytiyT0rI7wnmam3DVQggX+HvsfI00qDQbAiyR8PiZdZ
IWnQFBkxJtR5BLOF/L70U2FtzCy4sl4bW93J45doeg8uK8LsO9oddK95cDSCt4+BpkBzb2xQloS5
2UKCv3pqwetas3qp/FCZd8tr82Nk/YDXqo5gCtiavCveFi0M6LY9QYPluxTki7RxYkUWKds68ors
gu3ffsVAxAG5NGd+Yhhqia78UKlYN76RqZzWHA91Mvic+JbhbHsZFe+r1ApE79Ebbhi8UtdUAg77
M4bc1WRI7xlUPhpdMEdzJrLe0lDERHkNBOgO/vG8c+B61MP6BUFHkKgSYLDRmZbICwpvmRPop3wy
Mnfj5sw63vCLSHQJWcNm19dGNZ8Cg+IjebAosfnl2lm8BAEXiDJnC+JAchV8eJ0EHhJDGaAtamJk
zRGZNUk/DInv0Nb/aUZEVSw0EThWBLZoKxHQJWw8n7XTK/Blg7/2j9JHsMFczFBkMQtEJlZ4pFLT
4mDrj/oGKCuZwv7/UgnMDbyCAdr26fayXWtJzChFqTc95GI4//7xHXlc5gKc0mBuvLGfW6htSpMT
D7EVL4YNrdcGWnKIgJQED35umMLWixxCagGgZ6xV58NPL9xLLviplxPMRoKiwY5F6y7yVXhcrq4V
41qlXfl0P2Ib8D5BC1FFSYh0+aEq95R9/4jBk2csUbR303ktwPZTa9gcztxppULGyqjKe8LTISFg
w7NZRfjs0bpkIQyVbCEtqw94CMi3XshmAv+lif2OLesY2U8iWFAJ4YnYAoZKmz9h9VRQ8AB5zUX2
TfmwxtZUX/it6aSB30o2CvHTANGFRM5xYUhdYIeopW6on8ROWwfG0xq2mV3ag0fUEXR9HXCmeP/D
jgxvE7I97nssu9o0x3BQD/eQimXhIS6TvgiWOIkuP29HisVUMEvlVHWqcfH0MCBsNXiQLby6ZBpc
BF/d8hc8YJ9YFaLcNYZuT4s9BTJOFeDLrLYK8tLXEZzRLexv0v7CazhFz620DBhgVlkp4UCVtJzB
qjBdHcBO7naMjUPxRfW8e3OeTh7ZF+ciL7ftkJwihDspSBywLaw/FewKO9o4IQ78aZXKC4MEqvo1
/l2awX2gJSLAlFZQIpWS3LbrBOD1/DWVU+FWhm8vZHgTMziCYZWK7Ed03+PNz1V1wESXhD7hdM4w
qw0n0eYLtIgaVw5EsW6zur9Z65ABKHXal/aonZ164gjtuNuXaEolNkCxwFoIPjIlehPpttSy9Wj2
5JTtA+3BcEShw/dQ9Ex4iJsEbFbJO0UHO6yoKqSYlcVrTzkoriOBB2fu2IDeu9cKolqC0IZoV7s6
X06ADbNEn8go6g/iUTSt0qelpcck5G9iWQRHlPRRDJ1UBO4cei7SpHDRzOdhv/dvOx52XULpnTZn
7Q9YAw8tLC7B4z6JZi0KIt+eTRiu2Xgq3J4sTPZsJaKEBhtwFXWN5AfJH9Cg01I6EpGbCOMVe2V2
0ZiZjr1U889IM1pU6chov5O9zUUUCrqDS3IDkMblm8qb/2WNKPKoaNlSmjMoo9fHS+BBVrV2sCO7
KBhxcWnqQwfdPwwE/qXF2CHTdUPM17WIb7fNlntHnsNbJhneEsCtLbKXGmlYjuGcjB8k0OpHTpJk
KgYVPMaFb+nTW9TJZW32UoQtQtqmk+u3yr9YgExpvC6N9jt89JIGnLqAZquz85p+IoMBm4ei6eJC
plqERixHCwHxBQ/UW/uCK6ORxW6i8wLbmTCBfjPXhAe4f2xdLZH33l8VT3BFmQ/px7Yq1aFrYpI4
0Z39+W75JauUVOHj8cHmHTl3QfrPhSQx+4JljVSrpSJUJnvX+iCUQw2PHBQOR/jIjhLX9tx/FFdM
E/XkHQLX2C6dMDVFDA7hHx0kLVrEdeIWHT1DWl+Wo0YTGQwY38kADrWspUBIyGw7KeslzlaPJ/28
GQodpkc3C2UBkiOBq0dbz+M91EXJ/Fh56qhBJwd+cvqRq5IGrMhdio7buui7ev/QoqBRrQR6/z5z
Q+qYF26CFf/l2Fjdy5vO3bgPnaGS6PfkiDnlKE8utSErk9HfhexcImlGrwUrj5kuD1v7SHCY13ez
rYk0W1cXpmhcZHPV3WqVGHU2dAGHpk/nCnqOGQRMG91Noh0apef5X3eje8L021bxaN2C1ZpDthWP
P/7yet4/6yIY9lbJgB8h7MVlfIgoAGtmH7m1kTXvVvWp1irAjhPtHGoYyKVVxzOtoNnV8Y3+5Imw
8hQ6TxZb2SdXRmGTvP7oWeOXdDMjUOn1tLpLMKg0+HwHQMe0CJhu8R23gHq02Kg80B01ZdPhEEza
a9FAkdJ2pSFvnhzB/OoIta9baQpaKsSnkFJxML5pPMtz9tgZfEoVWPeCZghr/tWsXpiMgFV/y7+y
SXHpNG91MTyzdBbiBPkSO++qMBt6IqIS13juj0/FvAPM4UX9W3ueJorpRcMdbwqzKqtJ3vsEqNlL
0b6C2PTGMyB9f98ExkRQ1pefza1k8VSMCHrSD1fq15JK9ynLDSiRCeTZRpgzUXeo5FMpiow/RpRu
UXbHGxIp/ZdXpC6Ct9hEXf04wVlcEJHHVTrw4RWaJHjIWLKuG4utAguyJRjtqgYpW5zO6zjSF+mN
IEW5JDz4fYQSRwe+w+Gk9z5AzUlg21B4qBs2hBf4CDTqrXaAl8kpq7MDn+hPoDJMwR3qhWIw5gYs
RnLG6215aqCeRy/nLmYjwrD4zMcX4Ni7uwcxttG9t9SUeGfl04lwtvjx25fFpg6XGT4wuv//24u4
g7+fO/cJQ9rDO7Xeu/18GAxuCNz3gz3qyOVZpad50G/ngVNjUkRfffMZS3iOsshKo7yts52GsbGE
Wz+Q3usfdXXHoV11t8dtYWk+9nlE2CIQUoon+iXT2+bZzGON36TFNLM/iIroekcD6628+KwZqXbe
gpPgys89mCOU3DpEJZsVFQ0OHBjvZzhya1DxZPoJ5z7QGlFMqcX21GNrJJTkjEe3D7/HiTK1wcwS
BpB7kAy3q+NQlam5oqv8x7yptlUtXGupbLYctgAlRkqoAX2yyBu1+ddopy5znvySm78o5h3E3nAJ
l/tA2NtQeq6gHlk0YcSmFP9fsQqZZIXuAx5GzAbpd5lKoOLKJ95YypPR08rQlnOltvHECYW72Zpf
BTjX+1pCSa3ocqLVkuWZTVqG8t8O1KGy38jMm4Tra1f4tz7mX9np0d/l+A9RuwtlQREM1gxFqtwD
Z5vjcU724HT4FE8Wjqss541CRuXIG0DVgFnUmqMk4jwuJLFEF7cxp89reslpg7gBCWJ73siNMHtb
aekMTGPIocT18+8mRf3FuyJX+OhoJe5rAZd6+rDLEEbCUupi4YRelTIuQCA66Nx1LIPKxipo4d9D
dS34Vfj/GOqG7R3nrQBmz2ufSh8CZsEkVUlLx7GH0BkAncvg5MugUzu+461Uru4kqlDd86WHoy7a
Yb33Tlv9xc+TncGRD2WFekx6nfZ+y+qZ4UacqwT/kpm3vfIGVC2JL+YjnhpyWeBrlDosTKwfu3kG
au17k/KIZWtl/rbPSF1w9I11xH5F5pclLJvF1a7/jHUVY/ATG++k0HHb1WcM1CQeZNhM6x5d4CKs
wmgCLDq8sEbqd6iQIl0OG3weNUlmMnqZmS8pdO6K1e2mN8sdXzuSGRx5tyZ19mjwHGzHPDPAiLl8
v6LMz0AC1n0encgNqFutTf3ejn1I+HIrxEY+nONwNkjGn6rqMTZeOdgIaou5uDPNRL9P82fXb/Gs
Z9Vt0roNvP9jXxYISZJ0fXoSVChv75wUjcwAoa9pwxtjOMOECmse1sSiNkibNvcIf0T5AZZ72ltp
CvCqMYeh05bp0P6En8Bot1o6oMwy5SixdiomdmgnAwoATievUElJoPeYdcdnw+uoCBr9ukdznQac
tbNjva86eP3ilfkkhcsCwC2UEngGdg95QRmPqXfe8EozPkz1nM2wtFe1emJTmzwzG1PnYVTO7H3i
9se2iEqf6TEH9Kf6wc9gw8GPiplyIRzPIylY6hoSBRa+KtjI86ezcR3t/VrYVdyzT4+/w3ID3oSQ
XWY9/qgS6gzTznDUSbgcWkqFOLqTfHCvrhSkJNrieDNe9zcoY7qd8517cdjmkqIzfekRYbBK86ro
jQ7CKLEU9FlEj1dNs77vPwWCfudML5U4LlLzALrRKU5Szr1ccQ7ZdcJE5wbDKX0xgm5Gsj4U+NMU
652faL6LqFKM6abgZ38o0uO+uf/7i3976uW2PdFbyczuunA9YG6a/tvkz5ocCCiZHpJnB580wXpL
V+tzJhhYd85RBYluDQ59mWkt9scI3n3lu7fJpkMEI5EB+jdhi4tUC+kuFHPJQDLzyYacZjLQ6cum
p/ttGOxkYhklBLHNJw/5e+FbElOnz4D0zpxo0Eo25u+2lx0/2xHVgdGqAtaHBMSdiK5GfHq5Rqrb
XisLSPJe20soBUd9C2K1sGZCSf2Q9RfX4/NX2EL2jwUQy+Q0uCaiMOETPCUKUR+Vj0CdxifjInKj
KJ858XFarXWUP3CkHEQA6j2y5G4Q5tFrZlkYTxPpt0+JbylKp2KNNPB8Yf71ivmvIj/tJ82UbmPJ
hhhp/ZQMHvDV5GXWNQglSlhccWdyZtpBS2jVyAMOyovIQSSyMo4zB5mQX//YcaG6Ud+GeaRZ5Ttt
nPx7oCzmyZ3RfJyJ446/AD9b5OWtuz3fspqrOZjzjZsuiEPDGyFYDUvu/eK/1eXL6tlo0pT3Gmov
kOUzLWvRkj23fvfGcpv12xa+I8Nn2qCadtHKqsTIgV6o5XFco6KZqoEQV7pU0O/w6SO5zAI0TnAO
H1ZlBm6njf1zqGa+Pt8Vuj6RKhkoAY/ZVk0oLF4h/Ka3YbliiSccejrdc7lYFfDnYIAGWGaezLzW
4OJ3f22z3xhZuXtlK/kMRN5ELJ/K3iLl5jq9gaDQQQh2Vp00+GSiH98OZhFSMAQobp42z9NO01kk
tVLspHNDNCHMJj6dvOaDDJG5LVLJQJnQe3X5hob2Ut4lw5eq9DPOvaNH2zzc6SYfFHTueGd04Ii6
+ZO/0kI2TC+WEEUtwV4qbbRPFd+BY0f69NCvRKW0VZjp+/TUjegcFHdZ2rH24HhAPNnES7TPCCyC
VIoM3Xjlzda4fqq0Pefn+VS2bX28TBfXp5iyPnL4MdK9P21T2AkJFixSDkqoHuq1M6Fk0NyAt2t/
d18ZaG/IObGkJLteHyWsjIGMWUF39uVHNKvVV2V/fMX8nfsAHKZewVDWJn5i0cWT75FLm19o546+
v5wdV1/NOUDidnm9GlwnxEv1gO8IA6pL8+FpSqiOP2n5nwMy7IxEYJjrVfUxuBvY1DTaWvfGTBRu
zUqLBhZcu8ZJkaElXOWOB+XwLV6nPG7NcJ0gjjTv2vZ/KYy2FhwykzltU9b74Z/i0kD1h/otkOQL
Ew+oJHfkNuiAtSzrYS38fIJa/2rE1zDKH1f2jrkZEgKCAE0rIfhQo3Bpr7RFll38yuynqeVc5Yws
EWX/D9G5uKLUQbwDc/8wWstUKuAWosF7BqX4EFzO1qKBUMKuWk4dbsffKEj2B/CtPEh9mv57ACK3
sh4KtQ/qs/1XBRuP2rrX/I1yleVGkKZcffj27nAuvxMPQqpIViicoReLzpN+RBIEUMSKcQ/Ce2no
XIrROFKqF77DV4OaVNsmYqqB0MAGgPmZ9mTi0D3x0GNRENUKKu+JyvR0pkgwtRSnMDEEpZOVi0BY
h2qUgZN19GVWzcOSwKqSD3jFLxO2gz/IYMDTKlxy+64CT6EPGsMKNVYISy8rr3mLZmo+o7Y05rjL
OXfQ6Hm4z61zZ5ahbvlo9h1aU7c7+c3ECo6rHTANoD988VGVyI9EgJmAGfihkngOwa9gSgUGLrDj
wvRZfWmLKMN95QnkaVTzLpb6B8nVU/LX75sua3U3dPl1qpGyUELvlxBXRoZc08TM/MxhrOaarK+W
mqlvx5kJdzgWJL2JybAYP/yNVbRkPWMBXVo2dJGh02f1McjZclcxURy86NqBcUrppGY7XGpQoLPr
U2RXsbRdBttX+V4Y0V/+kWIIBzWKSPj3a1aN6hibptoHFsDVLC/hW2spb32EuEMipOcj/JDUzyPh
wrRcTxHn/k8lx4+jLFDIZuuurRix6ZrUMxt8QaB52kBDxgBQGfMRU638rx987wt9mfqYt1tsjoM+
Q2BBKaGy5gLvhvwBb3TPvjaN3xa8BEjvYMSmc1o+cDF60pdsu8BCqRTOCtD2UO12Ll6lGCYsXof6
PSbbysVPQpgUvV9LopXwhSyTvwiDEG6GV4zrZqmR6xQ3Gat+iIWtDRRH8wi2jiJB+04AX1iKOoL4
oKFUd+1tGfVQK0ZbR6yOFU95GNw+hXUWQaG2zDux9/JrySLJrgiMzQbHUjjjkSR4tCpRQ8QfX0S4
XopWH0nqsBHovxBtWTVp+1gm2w9d6ozVXZZm4ytSiK4D8KWggm83AL90vAu9xJ4WfZBiwUYtx/GJ
ONXbzMYdgDlmYz532RMCVIMZbIvK6Z4h9Bct82JToM08zxnyJoxlXTRF4EprgWae4tbh+uzZsDYx
i7FdgIhuE0MCPk/APmG037bP8ndZ58JvHlzgUB+2m6nvHA1hHJGMorUUOvhLD6y0yt/9sZ0m3iYO
udYAUr4DtWxDhDITf196rqpA+6sw8a19CrqwFvh3BsYu6nyq2H4uPVAK0LDD68BMCaaVVFG4JLOu
qpZZrZ7YHrB1zJZ36/JtApXxcM/fwSX+t/hrymx8mPt32KlFK2UlDLBcraHZRKD5nxqszzBBf+sj
NYsCmyhAKTr62UYuRKKFgfKUzcAyx9U0pfDFp2puMOmYmZmh1c6e0XgWU1fPIxFOrTCtTEH7Wna8
6rSnMDFxIDkonIxsFqVmO6oxst6Y3h4COYO5Gf0+fsK/LvGz0TeYc7jY86JGZtjW7bn/+3ZGzfg7
jj2q4LD1koMNdYmeuhGqt0rr5u1FF5EtCJ2u+p6zMkJCK6F3xGYP0rBN8fxYWEzGkQR2k7uRZIGZ
r44BUgZlb6iLjDn+Ie4PpDU4yiJ8R7oCf0nsw9Em5So1QQZVpHfkHea1ECdiNWSTTiKJ9uhU0zaY
V6Bz4iBgVPNvbVzFi+sajJnGWM5/DvWcc8SVmZBObIXBtylKUaEKlvPC2eAsVHIz+KtFetzL5cCl
Pfzn/mn8NOY2Rz3gkO8eMw4HKu50eya1n0LPe+cuEI7+LNLKFHOqeuPVnXHj3Lr+s73u5g1YfjC0
I/nfbcwHbYQXS16QCzytPGYR8ddUUcLo/uveNTi5MznRlrcs1+SOuLIcX5lKReYwej9h1VKcVx4p
TzE1j7PT30LM9OeGPF1TSzS1slBFnrNeSPzkjwsHaQsB3HtliehAkulgqGQgOeb7HJldH5dNxIup
j+dB0C5Z8x1V2cImTlCQP0GdeTNNW5kOSHF/ID8FLI1EItyAVcP/SpnBGreSYzi+rA//2VJ6sGcw
ud0NZCKgjDZlc9b2UHoYx7lWbp7umCsHxZlw6WkZbr/d7nmRrWwSEVDo/XjHoWymwu2fqGel3Qbw
EfnDUbdafUiyty5Yz6hpI1wODEcEWHhxKa9MzZv9qRdryCi7RNJ0z03EI98quR/BNVxHTN+HhdD+
1f1aSgyT2AgCTGl1675LuVo0Z8SJ6gl7vQOmLT+Z9mbKjsvI4C8KhHaOQPrHKSd9+4jL839wEqkH
rvCZF5ONyzSInQO5BHECq+CevNQ8omem3hVbzjpMWOraeAiFR5J9R8Rd5v18hlKQRH3RwP8rlCi0
1t2+UN6cz7GDvi4D7HE+/laLSmfL7IpSzLsompkqnR9F5x/SimTvkIpovcCGIF+NK5Qfdx3Kv2Df
wyX5NhKV9nmxIGZOhEWDg05kY0Kks4VB910xfagW4wdRg6l40Ret1JnKAiRQFLlQuuxnidFOcLhu
3plMCrfIBKMZX3EwB720fKJ4nX8lhH64wklRKvLBMaW7ZHr5BUFrkJWMF7lsvSOLNOFs7QQwbZHB
jaBGtypYdDqGNU7Yyani/6E8TbLTCQLMTIdmQpZL0f+W1oIXIWUG5ef0/L8Nl0adXQTPXrvsVuRa
H+pV3Kd9UaaymnRjicRsQ0ociNiOxBM6A0DJihj61gsf1pj0ixcCmMkV7lNx5YQeFOvta2Im3BAS
1Cr5TCTR9ZzlT+nEmoKq2bouJN/IkRdhnIEVY3dnS3E7prdEuMKmCdMnTUPj1HP+yUAHR5YLINlr
CFhhmhrgXUOWjiAymF7ui19PKZKbkA7GMI8r5xlR/DKSehnIAdJEPacIqZdgYqbGMjL5EgFmdiVQ
FUQM7OoofGtgogsE4+6lNr2xYBggV/NmcRL1iiCGJWIpaXdX53xVnqujttSwVPQKlEan2oeez1BC
bGm1WKKy4bHNf+pfUUzX2VlratCYzzvp6tU48yf1pvAiv9+Dv6lNQ+1wY5pkTI6uy/WTmlPteJd7
KIJp81z34mXQZfzUDLOXmXxviOuMV+0bJ0VJhJ8t8N1KNQA61qS4EqgKHmI/AHdXQksUYEVfcmKm
YYcYRhSrsyyWeyqfraThgbzFuklyTgJ0JRsoualuFPWOEzSq1uMaDeTB35K2O6HfjRoiUgRs88kw
CE/aNHiFm6xZl1EpssOo4Sm/Rhv5O/OYTOMSlCThQwd3N9zbEmW9ecaoAx8LPJVYB0WPW1C3MOQv
ypdACW1B4UW35QMPhoDLK/3BEBkw68MiPXjGb9LkqEu9M7lbUSmMLJIEE4rdr/ixPLyzYNHPi5mX
gVhu/lidxVkCMWsI9jUtfdGinAI5uVC/THSth4CbtB5lSZoMKg004/ZNIhmK2WL5UPQQks7EaYj+
ch6fJFC4v39O2xpn4g5+zJsSYBdBGUh8oCULmMjwFp06dK5TQrCce69SSZ8w7zzV4NxGL1gMJwqC
4daaxvgX4A6zHVwuKAr0midA1QBMH/eYRV/7Y6ghj9AzCdu4CiINTEsS509KxCN60jrMFJotp2dh
uvWYcnfRqxsiXKtg7i/8nGZUt+05qHESdFtIGJGE6KhR57LDndn0QIIatgHNAqUEo7o6eTFI3BzW
uvQCnUAQFQsH6t3G7GplVqtvDa7X6/jmKgk9d3QkLX05hP+u+I67HJIiRXkvfYWipYbLK7pJs/VW
SX0mkNhHAiarDZT/PvdKbaOqDUBMj6909+kt2F6bJNOIV53t/ih+pglOR/Tl3shgCaKjBK7RURew
bIK3WFUXh8hwpoR/ZonNo7YKd7rDvM2Tw4anO+TVMZuyJgeS/WhjcfDGJ8GAPbWRsaMS9XDONnEx
qrHEtJC0UVBclRIsXrr6LCMpv5E6OM9Svfa1QEpsPiHpQYqW0O/6p26t/6e8oNK/eIMeC8WJ+giD
10RZoWH2jl+P5N2Twej4FHBsCnUTD/064aC0Aoi3sn8+z1XWPGWwJzmIvjuFmlBU5ORtZRx4Wb8C
dmL8AXfyNbZxXSRSCPgRU3jqkJfN3UC5jCh5XbGAzn42g9pqjCxRf5EnV3fYPjGtKd9i7MlNtIm8
GV7uGPOgc0WfeRcQvuzd/uveen6Dz0/IshWs2ifGvqcWHUhx8LjAdf1J5ys2hkC8SYY6sPZbkTpZ
hDxffLMOX84s4CkNsnWqEdodpofd1mW4vAIMyu533s85wMcjTtZ9FWfKHBeu6pKlzvAP1UP7riIV
3cH14Zb7hsP1CeGCuIoeGY7RzLlRE2D38fBNs6Cp7tjZhTC19PfQ8gONHkrkUOwrQuGPsa85q46j
7KEhFvn2qe+zyHMAZfuZefhZ+QhhBio8+ONWwoOx+umxHPHrl+dd+REMDTZdQxzKsHDBzU4rp7D1
+0JDN8iDOeBrUSkoCHqd7KdOsGnyrOHb3wPdB2AkV6/N4vEL3lIsDtE3CAjBsazkc8UbUAYwO3BS
DI/ful1Bq0LkVfc5McQpSKylmGJ5YP41WoOcDBayJpaA9JpDj7BebzaWzii4cVDjzkmaqYRMKleT
T5IgSwRe3IwRR9C02hhRrHqj4PoNK6DEMGUph8DE3axPxBLuwGxfii8bV111jFRvao8S+BW9OBJe
rwxl23ZHwtPioqcWL3ItcEK4E0sV7eJqU7NcGRnwflpS/XIQKo4HtjKmwyjRVuC3z+8zH/ZmeITA
qDGQJ+22o1OSRLMGWPh3i0wyEnldpdQgZJrGMJTlu/DRziUOOZgpAHCGWAELhmAtzNP6DQeDnJXS
3ir4gW5xHoCq7YWFRh5YGOWf9LFhr3wVtzuUR/OR7I6DfKGjqxKtn5pr966xuukgg0bk0wgyj/pq
PmF0saJNrzah5NZDgSN3LBkz77MssNi2vgC4B1g+LJyQ+MavWpEzcvSQ/+MwzPBVo0kxX+4UyIap
kIf/JmivjZ9wMi+HaHZWYH1mvYPqQ429DlMduA5wHD+pVU2GQfKz5zrALn0XqlZxbSgRN+LmnpJT
PZExBuDlvpPpxizjet6JGnjZ/MxyPScJuU8dZkQ2jEFBxns+kO0WwAkCPUI3zw2lw3zdxLtYEGL7
RIpEDNCx/6V1HKmdsifFPYj1jLYqr4Mr3VPtge/VP1u1OsM4VTBip9z/hJLlUGLd4zkDtBewDHJF
6q98rcdF15Vzeu0Z1aYlfZTXEW4L61rE8QrqXvFaR1WmLktLKsR6zRyVQh4sLdenOt24PG9WN+0Z
iNJNQW+wpl8zthnylLSoZnyLQdIfew7bhd4PgNS60saEqno8H7fC5CVTwOS7pFdZGXteu9PDwDeV
bX8lmWyfabUyZWzDhEHIadCRFUAtQoDi45QzBjm1NhIYQcuMw3HqGu7niQzbhK6XhGrNSPTSMvmj
kV9lUmDB5Uh3baEbG3Y0SbzmueXAnB36ScTJMhEE8cQaObZhB3y54GaToKeQuvmB4k/nqYF4XNKa
yq6OH/JynWjqJ8Zl6yAAXn4GJ6jadFFQ4xOveyN9hKISuQmJlQiUQJ1yib/cxqa0fsiFbL7q1imG
2lmbbJeOgJfcfuOvuK/hs63Z8oZxT88wupCZd8oK5aWgjUM/ETDls+C2a5RspIx20bLRA+nYc5F2
pgT0yWrCrlEUzWZDjrp+y2JrFbA7gitUQ1/cLNiPErnArzOkPgZHYmmgLN1w4fe0gEoTlYXriFMf
ugSecNZ9QPSr4/vjrJfe0ZTy7eQWqjBWdbM+OO3OM8QFkmeetY7dc+B9xtXLJ6tlck/HBcA1/YBM
zWFBc2ckBtSQQr5gcj7rkiTwrQtyupXDjyj2rprWWVzh+CPmuMVbWNQrqg80qMAhNEDtzwJjBRBy
/d4pEJRV2bjADc6JK+/3T+Nhyi2pxsxljkue0DbUo8+e9RkILIm1PR7n5OaYnnR1RBfPjjHk0dxN
XRTaksQioew0Rt1GQGBXG5b1h5/0GUPzFrri0HaJw37mW28xjgRtS48RMLKUgXNVIUlZJFstAbs8
arN7RBWyA5Vduhs428Wgbn7Lc43TOJbqYRTxDioTibRz1GpmaTVllrcixaQTDA3fbtIV8j4LdVrR
K5sr/MSdZ6O+zyo5gs5x0gs/RTUd3cUQGmCcqkl+CAa7QB+qkwKIZBBphJaOigypLHvvCNGIa4X+
4udu7Lfaxjw3KGbvZIy2GgOoI4Bb6uxW/zzvc0PKDni9i5Hky0Pj+bg+5LQW6CIjdW6WH96mpjFE
PxOCaD83k4G+KG8fVFVv69rZXAgPN9/Sp26YEmo9AnW7qWWdmqFVHG5pKp47bxY7u2XxozqHWFDi
hLjR5it/yKA2Unc9knKoBAjFdrZAG+jIKdsA3Z/4WmH4Qw2AMbL7Hjk0h8PeeH0teBfbhqQ4amea
OY7rxo1R5Y8e6X/w0GOkKe4FgHgo204i3sTe08OP+QN5g2EOJTeG+0oCmX9HPjDNMlGW2bNrAbGd
qwG6SxTbG5Za81NWmJH56J5wb1As7gqS4BCLgI8v9jrosSCKGXJ9PWdCk5LYIRMDBoA3sksIt72H
71Z25/XPqBhHH5Lh0d67/wyaWcSXxgmqFkuFh/ZHv5jjJrL2KFEozcsjej7ZqwLanmoy/vyTLicr
Z6+D0FXYEEdrRbqWqKOq1CxiHUxJpQVr+meAZ07LvGi1m+qtJOC1DOq0oaIf0FdopMwyC3StVUYF
JHwtBuhbP1kbUAVMwASC4o8Fq7DMB9FcgNWDnzY3wBANe+EPLgxvs+x3Hh9BsnfUylGaulMBfECK
wUO0bVHInKUuhbFByLtLP3SN5QHiMKXqdWT56Qg3HM8LfNGjDE+0/PvaUQvxjEfnKUU3QT6WMs4A
P+7UjcJ+x3FpDaIrfdDfMq+tYoTLPzD90ptLnfoPsVtL3BFsyT2rGFAKe2QsoV01/5GWvVaRVQVp
iskccEGPNkEhqQ8WJd+hC/I7Jz7vsxrXr1MsNRWeYA85/GAGKW6ChFPijWzMAU55S2QAo33n4197
7ua00A2cZ+9HWI0C44kySLegcGqgFCLkZwxtXJ3c06Gro5Co8P2SaObkT4H3Sj6paTwKc1p7KYTD
V3oxzhzuE8hlrd6lr+eF+uKOG4ZTly4uWc/IqK8s21V1GrBnOs3UxPBLtKDIzn7eEI5MW5exiPok
1Z5T5SPGW6gAWnDVbQPGkEPL5WWpW8jA2bqexuzUtC4APim1hTZvUMRBugVCuakedyftiQCVYN07
kScCDKRAQ4V25G9gwydq6wtrlx66uACVlWkuxy+TsidEPSgToyzFpYUaJOTOckgG6jZp0l6sVD4w
/UvioHDt2YSToh6zVLxB0lcIHpwAoLOHnMfmKWXfsEKJ8Hh+VSyHT45QBacgKmbZoHyH8wfVo3x6
cINtR/JCTsUjCMvocc+/pVK7EUhsrrQQvzpg5CeZSJY5BRhdNS+HfDILDxSNmv4rrVwrEY/74A/J
eBzZAnmVkcyPnfxvlX5WzkkbRRRyucqpJ85Mxyryc42ILI3Q8ov/fhC7tEAHtXP/mEnkjxkjA/QB
fVkTY8ripja3GUiDSbIkzbSQ1IXk+7Jz88gTCPf6sH66RxSKFoL0/juFVtVNyB4md6haz1BzgpeG
5nbiKdSArQHAZv0ZSKOUVMMLgppBzv5Pcgq5W7XjwBE2qnXVtygxXt7mUiYE29LX1POft5xI0Nd5
xL6LLksulbStmKQ8mII/QaY/tuh7AxlZwVnVvbi2vMtFAqIto0U31okAIaioIgcDrZvMxLgeHw3X
3yKv7ZsEyPp9j6LWH0/mEToAOnYaJ7nAAml9RmRgdbsE4/zZTLDKD9mFOF1ZUBFqGYc0v6MHOWif
VKs0zQBTl6dZw2VQu1cEiaNr0P7TOZWoUw7TA+5Z16pnh+m9WWDD1prDy2LkEC9e3L1N7Fj1vzHc
tQLgYAm0RR3cATMp2/XN1qr0EcoA2q4pWqmBDxvpJ7TRrXYxA9T7VgUjf2Yg66RAyDY16zgE0+CB
0UbIA+Ry4eNhDIgsIi8jiutVptCkJq9GcRO4zPHJ3y3HtVnmB0BZDTbk4ErTYawhmcSmrb3/qjTd
xn8Ia+gVgXlIfp6GiB68LUEiZ9uwCOmiFJBXuxbO+cIavtejLTCPDiGLROKHFDo4jfOTiSY1HJfq
hXfl6dnv5gKeDZE3+ocE6ZnrD2Ra7zoaquvugVupuHzW/tEvwWJRproMYJxvnyqG8qx09g4ruL7+
UTMB5YeC9np+cIUS6c6DmZhv5vnSjw/5sy37erh7OfM+jTtJs/wlzlDLAlVgLQ8UW/HxKGxzpqYv
QjnC1hIo/cPOGVjK5VsYhLt0kJTkUeMBdJK1Kn1b8+6n9ogambq3JTmtbNA3GDWQF2LiSZunAZV8
Zd1mDjudXgo2FfKdoqS6vUmcF6D/Zxt3P5dxDLSbwyOjfCrQ7j3N4qLwh8P0Ib+MjW9uBHsqAfrs
aPRSes7n549MH1HCCt//mlWxwheZH7P8vU+CjrRox87c0LKCJ7wqGCcRPutezZlSjwKSzJ8Bbsk5
OiKUHC8Dna0f32nuaYldHMgCfwaGAZpp6ysHW+6NMScSANYyV2hIgQjdakVyO/TSscrZzClSZe9I
P1aXhKNeVrDPCFMJWlpMSH3OCryGOcWKQHAp+ANWzRPEfJqheCoxtk4UrON3/RWQskEgZ5o7ywFW
5LKWepkR5hYf4CwgolFviUKej/FobZm9JKtYjPXGIiobCmt/gCLufRYHw6Rz7hZQ+CEoImuaHEnX
BC66lSZW5PpHtwf9ExDkufIV4W28F8H/gsBq4ep07WdQ2GtUPNgXhpIIiVtje346vTugnxghGiR+
qfJZrIXZIZkycV3VpVk4MXvFwKpHLFmLz92FioHSVuBr/zYF9Z9Z3p+GeJFKTC9wiK93ohq4/Lrh
unASBiGuLoWoWmieS+6aOCKURakAJWaEs3eAcORa5R/Pqc/NJvK52Dxoq0EsV7jkKbSDZwoHuywq
cBXYsJjP2ClCtKiYirOgs0slcbrBvMC0UYFYR6RVP2nZad9JvsDzF4AE5vnZ5nDOaVQDIlUcKhri
Y3nLUSpv+eIHO4ceJmKOV72GOjcQNVpzsG9ecU4xspkJvWmIgDKvV+VxKCIbUfA15FQNt+mqt1uD
+agMN57ZLmVaHFoAj7EfkKPbeToHWpNX0D/0v5mLGYYhjMty/5tFcuapgV3QtjRjjrd4VuTE3q5Y
hPIakUgD1r7y3Lwv/EEEYEhhXSauqvmAjD0WtXI4adnctojyWdx9GFoIqY2zOwZSye13w+nlz/Zb
nqcU/dSAQlKalcKKQNEM6RXa4qbrdTl3DnjagQ9qFgO9w4PrE2ACkpnQZmrbvxUEADQZqOt2jc8/
9wKp7bDGW4sxOLgSNW7vWJtuDtZ99YykxCvBXGYZ+0vXra+UwdTRQRd9y8BUTL83wT5hf+xk3C3u
ejBpF4QyeM13GJempG5WpyIRj5VlujswHm4tphP20yI1jSc9nqQmpEb5I0kdGI9gE6XmhSAHo5+N
egpnnH+qZiZHV4UoCKDS2vcrBN2M5bcN310EsuCFeix10eHwzVfugAg2muCPwWLp3YzmrUwqffVp
AtheTGKa1LBAIpPY6WvFzfykJE0JJD809Dh1fEdEthTwZ3wUlzfqLM7fRIbW2iFeak6uRz/oHMZU
qlFBfSOTdWZl/WTQC8QqHY2bg/3gLBGCjOkgS6cjAiOOyQzSBJKXBiBoM6Dlj0iD+QZUumteSdwu
+mNN46T9h+bFRqOco45AHcOwWIZv8TJmxPm98kdILw+VDWk9sOy9VUk9bWj9ZNvWqEfDAjr/OV9B
0M6FGqeW4qmO/TyWWqjZJct4MiTinAzKcfUgfzdytCQSC1ORTO5O02Ucocp8mKxrsAcUPKOQ+CDH
62DEG5sftBpNLai+NSaIazYhs75Sdp8yfCF5GJ57oymR1Fn4NG1lpc/5PIAa9BQ+pnWfmNc/0NHo
3/ZmbLkshdmx7AAJqXhBM3+S/pqUnk6folhBkh1a/PlYtY35CjK2UUKFMp4fom30IYE/FM189dHp
O6i7eF5qKYrVtpnjLSRkfoRhi6DRh3C28SlCmMxq/dxZvEi/3rs4WkZTeIvF0+xkLFW104Lqu+o+
0eyD/s+DqPLC8VrIbOm65wtWw+arRFWKfgK6FDnMY7KOMaLJ/WNJKIDk2XE3uBnzDSw5Nml1SQGB
kWQCnZIOPhW5b2jozE1cFFrgieRmGiwQ+A6i3rApSZCeRVF6NWLqGVHwCTOpuWM9dEDHNSzeakTr
RiK3s5duITN+XAkIZ4vHR+qyP+wbb8bG2OiAHYJ1bU2piyzjoBqT2WQV6VFc7RBRSrdBk4QH2sD+
+7G9EOeR6H9THg++UTfj/YppCrfLVYz0mYOdQA8GU/IiVbSKn6+QuOD28T7qKh/zQ+7RAGQMWWBc
/vAtaoWkw2gUZ9vN67Wfna0Ca+A2r7+SI3CkU81XPoQo9iudaHkD7Hm6yFCNzpaDVXrwZgHyyktm
4vsDR7raGt2MvrjG63zT2s/rY2BJNtY9oa4gINXApIx/TGHvu9j3J7LAj3e4Mtt1nOyNEyotXkJh
g1ZXgbvOB566BBB4nH1Jn9MrDSeKlPvRtW72PNOlaf2h5eLxceMefsfH1chZU4RfNB0Wq6bdQL0E
fOO9HZzmFa15AoZGDc2CGACDIXf3MARHZ4hB52BEbJ0ZFQUx0mMfAS4P7vvuSanF2P8m8I+3SKq/
3ho8IsuT5bRQ8IadxbskgFXulIN1nNUziK+gAKTCixZJLsB4cmZzOogeKMSXrknhuLkbtEqRX07K
IxyWGwedcI3lbysR7FAnKueh0yAn2lKv47v9kuBIQmrwIL2nbb5YubfV5LWAZkLFMAa6ERLSTtcQ
UeS4GaDmCzx/m7tbCpfGErXN5thKKOYyUKeYVxpaegZw+TX/njxrtYvWz53FLMPyFZPU70kBKQIP
aGZ/OiS7/68580fw453YJb7J9Fdm6F5dqGx0Kvrgm/NO8bZp8rnoVHgZw0g7Efmd1y8ZBa/Nahj2
dFbEn/dNYmzMHfkxpXEeuXlamx4r+NXP/g5gVnVvkZaMG2JX3xfBx64/A+uQMCQw7kyKM32ILZRG
0MqD2NxkGMSSN87gnX9WuQprJxAOrN2VW5zeghZNg6+qEAy7PEpMPhEGOd9fmssT/GOZHgKe0owS
xmBDCOUTP3JSVxaRtXMPzcx/P4dIRASFfbLuSnEMxeFbQVK8CkFfN1PlUUi0yvqHSPF7vNiWlEbD
7e+DR7q8LTTkQdxHd/574Zuhlp96mg7sqZF4fyVSRYSChfZhjxtyYTTvzx92CUHACKLdIiil9o4O
zoiADMtS79Mo6sX5IPxJHAS1HVzxvuuNPaG4SzG39dSPdXcgE1YruqefUmIYZhi6cgpExgYM9xxM
0V0acFSGqJpFD1tuaFdodoMtdmpE/dr0kdGNGsaurSV5QS5byIL3WJlabI0D/Hg9oNfmiPLWNx6Q
ucg6Dq6ukcWX4MwZOmmNVVUbNjVvHzhS2lvrMya+ouWMdY656Pm8r/bmOcUMI65zHZ90l1wueZfq
L3yGoKeiCLuNN2KBgq+RAfJZes4Ty71Crns87AnALnDPSMBZRJfWrIrC0fwXS0cZnDvHx7Om3ZO3
2JgcZyAmuOJnd9gmGgNN5h0coZ3cN4zBzCLKI8mhgab+5TvssJuSPNmwi0DI4i6AfhLYaPT+k9sk
FnuApClb3WydyjK7Sxtv0TnPMPhQCevE8aUvacl9q+WjLt3iPmBGZUXpBWFUIQ4oP69tIV6NE/gJ
BfWwbMYCLlxhtqkUYT8l5vMWH4B6EoX78W8icd6XLlNOXSjen1a/r46wS4CJTyZykvFXYC8rAmag
HU8zldzBL6WKpdMxsKCrLqG8AZKAjFQojFOiv4ASQTSZCn7xt8C5YeYhkCKlKxUlmqrspMJNokJR
CsrR3McKV9r4nLDicBxQDe1JE/zJCIPc00TQP/sTXF03FEbAdqWeXqgNPreIQKCYqz7XGhZKVquF
UUCB1DdabHom7tDFlifcaFeIYn6T77R4i+pL9Abu+SqkELeiYhEMJee8D30G63N2LMQ18FA14BCH
nDe3lr6bUKkH+E6SXxyRJGriIaQhFdQseUWRU6zECz3obHHG9cLbSr2s68n+YHztrqbDD6Qc6nFW
qZEI1U22Ws5N8u6TjQDnC3iC1zt1ZlwtqgxGdavvWFx1+7WycM1NOnHw5wlqt7tPsPkpnKStIk5q
Jz3FFcKFjhmBpAhthE599snlbAt6kq/XQYIuVNA55rtNf95VhXkvApwcmBznbqk/3LuKPbbymIZF
4X5j5ZxE8yT+ziUs2Ck9MCe92S5cBFD1PnRIahXc/lm6kC21erDt06lYukqvvtmKcoA3CoUonmCN
HyMz3+Ogbk5BzdUPnCpZbuTRoLF5CsOAhklwh8aQp1CBlHmNwoGPI0ckwUET3cZ2l4VEwuYs2lWt
YDHL1PBmRMgL9vpaQdofB8ZoyzEDzDevRl/lcP/+pkqwrm7EMjwwo7AwRd1m7s3MBMfUO8T0bIaA
0L3YFfzaArhNEbFjl68jX6NLNkVJ4O+CBN38uuJkwdKCDnV0R+y1Wv8W+L9OFhpiLHFBKwH14s7G
CniFQtbeuNp3ZChPP+8wtezk+QpR3IMx6VVPPDg8fR4Gk17kKSGW22icztYozOsSmmyDeL4XBE6s
e9Eye/fzTtQdBKOcsfTDXd47Eg4zwsU9uvmcJBTJWC6etCki1Q/UEesCepZowFj8d/+ZCxmDdXa/
y4XOCODdvuiUIwpokhS8VU7ZzpzzonakQx9U2hwPxxp6Yebqlb9qB7pVbF1tw3cvZVJ5lGe+2Ews
Pl5oS7a1LLCqYux1+VECc+q+ySm5OWeSX+HqFwrfZR41yBBU+MOv08im9VHFz3+dakXo8HgQ5zma
njwUAmhljHxLROiwFSF17rPwG8NzJYnyjKU5AF31gF8q3PMWX+Yi9opEBtOVqaFN5fpX655IB6HG
7ROCMlRVJP4nDYI/UR8C78DTH1lmURQzK9GBuUhusomCEfoX89vqDrIwHvoA5L0xSsWU3Rttw6AW
mnuo43cbLC8oB/jzM2z7CsuH0Y/miVYqFtDykYuCUW+P8b+l9Xjqie8KuR2lXgawUTCsiKshi84H
3QpNs/uHPs2ptJfPuSYaIpHrNcCR71YiIORw9TlgD9zMTkvxmzEf4OLIU2uCmQi62DkjPXJj4B3k
8z6trVvXgmFcmBAVXz+0AJ0nWXBvR6UnsavqE9KynxeBQG8cE90B1rVzqJyW5OeITJE5fqA+AOvC
AYfrCY12G6qo02xiHTfujqPtYbC6LjUubXB3KH06W1U2fYnyPiM36A5RlJy/fzRGVBYyTvENET51
4fp4OFKf8QccpCXwLvMvuxDHYw5bezgKVxcDQRlC5ycv6JDiKZetd5UpF6TtshWuyoGI+K4x0Ust
6k6SUaNaBJyn6K19J0goQVRpUAaa5swwvxGEmQ58oRSmECidvpAwPy/lCrxMnSNJUSz5UC/qEYFH
8nd49b5Jq5qDtP0VCqTbEdsuEMDnBtYAeyyZlreCkYXV4S+xwtRRnreQAyGYGKX2fTsnmYL5ror1
fJqGDRo3Ppnp36S/Gl+YBHHVmAenxZoiRte83zsHgbgGGhtVuvqxHUSaUArUyQiQXnuybw+nuPNP
wf7uebSvYlGXX/06J6DtBkPfQHrsMjevw0gFg6qzJv3KX10IOFTuhz/Hwk3dMSQ1sB5zT4nWj0JM
CKpz7yHveciYfFLDC3cSauow1B5cPxuSc/LCYsN9R6H+kJg3aEhq92wpWtd3ruhrC/Dwh6cmN2qe
b4jkGruEnUy5egZzTnoaSAa5RtysTr3qU089oKGAfuZ0/QPB5A5GoMfMNHoaKhvcuLITSD142lqZ
Gf5KWtW9AV/DQKj+OjRopS58ZWeSCQMRofrgbr+YPkPb6aQeY0J9P8XbSlGANXR5UmBDuIHTapKl
kfkGlyixmVCU1pPvb+5nYjTzsCMZopLitoZvAnl0JdsdM1RQvcBgCffzT5kLCxsZ6779IcoE8iX5
wLOcLjo+CZHPZI5SOvNha6+gw5+ik9v6DVQuWqRjnDD3Rr6TBlgnyF/Cz7nVtW/nsvlzKh5TCF44
a/MgMcf/WdZ23cnE9zCaPn5DSKMHZubTIjHx2drCKAXR9325iv2vsrLOSBXvDW5dscJ4T0MnOlww
WWYP2Wo0zHmBmtNd7Xoy9+6k+Y99XzkYrgGFyI8CUGuIrHRy4wvojYg0W8hD2hjy/4GdsMa8/JIT
yrWEFLQ/JxqeWYF3BH3RhcyFfyqWajmX8+COFL76y7S0EiM0pVXOK79ksIHsn01Ne7FJtlsf5EW/
VPRksXzynUkH39Hub3G6HUhDLfpCJLUveNqOA3tnVs2VtMzSL9B2WJqNBkwnLhPpQBGB+46c5kUA
+gg++CneWlRcwoUFOuroRRL0JjUmVi1Qu6F7/k5DD8i10jC5sdqpnhl5U0pRIg7m/IvrC7Dsgc4f
OEizoW4JisUwXjQISxopxh/QgShvVlAo6+bkz2nAE4iuyHm8sSaOO22Qfoc0tCoo7x2UPnAL3ipg
k9Ghk5BQDWrnMdiK5r4MfEPCv3zD+4uYsL+02dM8ACNkT5tO3QTBA/dQ5TduReXojRpqdknr0u7C
iwedug60vd85x03xLCRQdbb5XDfdw/kg+IABz62Bc2OOJTAMdwHlGpIeJ1Lhz5NWuHSMQZOgoTBo
EOUcJptyk8OiDtuEAQ5WzB0Di/i/qZ7MN+YM9P8l+YvRp/UX1LQFDX68CVIL8tOlJGmPqojG1904
AU6QS0Ff2KRv3CxJWaypawxMdrgtj9wQqsnW7soyWnTrlPetSIImREvPzbllewWZ7KtJrgLGyrye
RRDh9R5VS7lqSXbeP5TyMQYxnmaNDxQk+sV2XobwA6eNx1JdJBT6zqVCX5/fIdTEqLTTADcIUMwl
R06kPHN77TVupX5ZAmQbpw26kK20OKkS2S6NVcVz2foDL8v7STi+RlGmpnxsTw75DJ9xuLRVGkk5
ggX7f4QtJSsgMtwXoOLm84BR5of53LQZ+rny6MxgD7599UgxTEJVmGkLGk159fhDpTcxybdPIpV6
qNDK7rKmv0MPpckJpbBN6jp7G0mgp3ZHrTZrK+wJf7hGl9G2Au80UQpvAtCS61HeGUpRsCqrGsWf
n1sHWtK99xQqdYdJkrMEBdKDIwFprJhUnZ12yHgki/VRRF6OfnoWUpwb6Hz/QBcGy1aoPzLFFM7a
Qhd8BAcv0R0DpOs3mb+eAIHK07+FKbakNUZUDG/1QYA3mXlKPYphip7cWGlTzMpGmf+LBqP8Xn9R
rd73y4hrJOlUQUfL0HiT/oMryL3eRT0jJoRZRB3gw9tFqm2pyKUQ5P8yrpIE6142xrPeRfEcUhSG
wx6IVFKyB5nxaaYzvKNkwzFOxBEI+KaPD2/vP2Q9QBydiZQsJv6btrP2CdUOGTGwQuhlrXmDB2V3
ayECn+7l/yRDuP7/TipsEc1DJDysiRCcUcpq7hjzDRDyRKMFJQOufZgUAMEaOuLGXTG0HRxq621R
qDmCROb2M+uX9ul+cx+plbW3aEf08U3/WxsFNtIARhIM2hO/7szAk0K4+FuU/1DSRzPxe/J4jcHQ
1gk+V3Mtj91ERKGdyx6ggEfqXwdBD6Vgnrkyy8K/kHucHCG9qXSv1SwzW6QQ+IL0pQaXDoTuavfa
jpTpPxZ8KT/eNCqAeaGwWRBqF1dFIIxtD2JTsdaVILzbkaAwTFPhb1PSWl6WNs4jabnSzvwGr9G5
pp5tPk717k6A4vwZxGi5IoxGiEYYCiSGmo4kRALjQVX8aqIuTs+iajhzvvIaAnXt7V5R6jfD7iIP
Plh1ZcuP014uC/tllva8gj7xiqKbbHSppq2m3wuel7f+tQHxYbPKU+U4ID4RexnSfWiFS9nw8kiI
1rMj/TAuJvkzFiVqn50TZ7vQ1m1nfcZZQORQjLHw2EySb/R2K6/npeJYY7c62pdkLw3ogKpn1F4g
lVuhK+lYVHeA7K7e9B5WJhflTOW9nkETQ4vzkge/Jo1+JjCzaqJkwkwB4/MQa5mUr70wkTP4Eu/M
+skssr03rm49gxUaWLcpcZ5Xlr23GFSb58FQtf3zn5sAIi+KYupkV0GLlyQtc1p/PAitpEQsxOBp
EephlUKzRv6kt0SOkI61NIYgAI21D2YdSabJRnz9mznXvNvW7W5DhfqTPn/TgHXMNbV5eSPruP5J
qGyWY9kOAY3lEM2b5Kq0eVciWMf4OqfzO6FX/B5gT8SIo4y5uI1VU8sSzQ97Jf5lvZnGr6uq34/q
Ho0spAALFwJCYc9BNrZyujFySF+W6FH4iiMch+KFpLUwemdzfEqO2sPo23S8qaq0kj7r+qaKnE/K
JTAsPQct26gcaG6cvicufm3LwD5XDIC0F7rIunJfcLHo90O9P6Qtjw4OILiz0NgLhnPrW3+5ppwg
xwquh6x60IWSXqZkFnJArzqMlxQfKPa6qVvluw0fnta85FNAARKGHez8O6Tonk5qzB75mCRynmHQ
FVeY2AIKScHLBQA4sVuPfYymp1BZpA9mz2yis5k82Y4BJGAuPe1EpPvqtML3k1aQehsykfSzDHl2
SgL+ICDMHMcbxHNrP/av/G1ZvVKeanZvzziHy9LIs9RMyFwYxGe1w3wRbn41SUU4eebN9ow4npFr
+lXtZbTgAKM+Nbeg6IKK5IUHehL4PY5VU67vq37uAAUI/vKU0Cl/aHMHOLQEJdlQo4x1Le5mSuan
ip/THpIOboY9NmthGCQkI5bISMdsBf74KRkKHVQcVEPA8fCkJp7YWkvFPvDu8XYhp8y/m/H0XSfM
LvXB/oRPolHhbOy3LNw4MCVwdfQFxLesCX1zPn2+ascke6RQFvup/jTPiMxob24s4Gls8e/ZAUtZ
PXA8mnzs4j3XgNj8nj1PIHh9gVtgJbkJKr+vGCZydECX1/lBM7J06toq7Hqo0S++GTDHp+lLE7ua
09ktgURI349C66XvIZ09G1m7T4LS9ZcTb356hiKKSkpVlkU5gbcEJxiz2m0hmGaZKBIaUAc1Ykcd
Hous4zH+4y/kL7hxFuq+GmAY2OKIzIcPRyi2di8sNJubSFZkX3rM8COUjxD7ujOoGQ/q3xOHsbSq
4xmCdUMCI2BQxu7Lw4L88BNfntQB9NSxPdekUySY+8P5/R8KE8SSoP0JOa/rTu1guKFTfnQOFMYe
RAtx8xIyvTa9bfaFp0hAAl8yh0YySv/3HhEE/rikyRGA5YMn2XV14k/6cPj+mobXuZi5SpPFUUCJ
Wm3Q1i790kon/O19CkN30nsB4UVgOfxLa3VSxe/iyE0eQ8TVj+S4LVRcbe5ByjAMp+NHVU1PwtEy
7GW/6o3WRhEcy16PPGiENGyaGJ8LvGYOGy7ddqfeGKlbPlxE44QfVRmR2fi22JdCvG6OnSgfheIg
9nkS90CppMtjzXy4HODz5URyO117cdKcSYW8NC7iIW3J9q9G6+yDM6h+uVEqIlfIE8X4uTSA6b0a
UuVo0xlW0cgz/V7mFjheVj93P9v2f8XnceCq5GdjZNBGH6Es+yF065ca2EUzbKLHysfsLtC3OVZx
NtVbqid99APRQpsrttIw3LTmiFLYYKPiI/SBxzuLL427zPUfibwIzxu1o4iQVWScEfRX2jTsEl7E
MxTRfkpnSCAPNJ4haHyalrwiIBQZEfXp8/TqPQuxk1yC6HdbDYyuS/qExKwQE5NYmDdot8GgQvCj
TR8zGeapMW6VQs7hOkMxtEDFqb7PFOF4tRvVcFMk7SL4MN0AzrSGROqEioLlm/dgxz+92Yvl4eQl
f3m9vNOWgF6YOH5v769uIeaA1TpQXcUmIMD4VZobahS9IQSzq7u9ZA0UKDwADzIWkqHD2rEWFH59
mI8RZt0H4S7Cdt1O8pvhq99kBM6YllntyFM3aP6l/zceydqoMVdYZb5oyz7qrRXRGGT92TW0NpqP
rNXqF4NhLQP5LvUXXSwKy5Py5QnG5Hpvpp8ld4goQoGkZ2jGxNr18C2S6u1HPa3vjegKZsMTcFWh
khObx3h4WyCDRZmx6wadKxRHQcA16vqnI0tfv//nYyBwhzNDFONmZialEJFZHXVsrm7UyrEXigvO
mzbeGVGAwVEiwiR2JQKYOXBdF/RNRfUYDRGw81xL9tz1/CN+SAN2RkDVTiEMyuCSG1QDaUfzftO0
DEeLhbLuT2z38AbmpKKCFbghLhz6CBtqvZGSgqMN8OdWmt2xkx7fCkMpq0dkSH37UbTeKmYchcBe
ANZWbamRotbtEorWPkuOlNNTXvwqnBpULswi9NK1qY4Fg01Y3m+wikI5RwIi1q4g7sh/L/q60Ehr
xC6P3NS6AM5T59hgDbkQ+OwvfFnZ2kjScS1uBHSClGCSNZlh9IYCucCgOFV/y9ttCgVaO2F3z8xD
kn9UmOG1KMTeld6MDCjZT6pcL/CHM/cMxNkyrY9UJ92r047lI+TUtx+ACAE5yRsOV6UkpHBwz80h
dSUz5ubZ5TSgjAZFh976biVx8Vjh06e0QLCYk5LYL3PM7rfRhVenfxkfSQJ/kNdnO1JvI9eTe2Rd
wiejxTbV6AZnuDwYIjALh21yFAOF3mUVfII2gw7laCtTauGF8PbN1YpVH9j4o0YZHeU7MHlq/gxm
9kzxeQ13A4jlQMDRQHy/igczryO7Nw9HP+lt0gTlQhVQkDtHC5IP0JbT3RKhsMylimDoAvpKX1Vk
Src/d/BmK6TIMuw5+LAp0WpixbAUULgJxEhrbgNf0Q8OiXfmareRrlCdYSfcqHauQcsRo4otwYdo
+AipPt6X3hK0/LqmqyGrzV0lm5naTa5tQcoT4qSBVi42E2Hoab4FVPiIFmax8YH8zBjSCdBvJykH
TXA0Lvah33WgPqWsa9FlnzSs6PA130nGKSZT7l5ZmnsjueANWW7Zlc3x1fhv4T7YJmTwoFhPiwO5
+5oRBZmpngvBrcuAMPQ0rFZeZvCGR8W9alAdHjGsJDDtVz00BtzVBDhWMh9MsGFxkDfFBpWxREpn
lYq85YBOJyB4d9JbX2aAJGGqFP9xKT12oEAlTsJVxzt8SNzYwIMyYop0BFTCFblTEFSYoYEl4GG1
MlioUERcGROVRr07H1UMHOoigl/pGC10SbRK6NnmxiHsM9E1m9rqdtXTl04HcKLf7AfLNm1QPI0s
wwe3t9l1FIwP8Y4Smiv4lSmDmWEYNokTGMHrjjM5d/luxKFkqVyKqpMOf3wevKPaZyhLRK9A82Qi
tcFEbCyJSKNgLF8h7ctL6y2nCwjEov/qbGd+8iCopkRN9Ij1mQvwhrycMPmkOE+pjm//1ak+Qzmz
ulvsTcGXy7AuWGL+2EvrPYJfX8uv59LpcXYbcZv2ReeFFYp5PCFQ9ViBelTnfPuo7Ue19Lf15htt
YPISVoQZyjeFa3CHA2Ukl1nC1bB9aZqc8RkTN8UJ4bjDriKIeG5jTNpdGWkXwgoRZkqiMnl+W7Jg
5apF3SiLpZJgeaMnrd9b9QYXulvS+i+jyAEqOXRzG0xQEJP7wbqhbYtio5CdDVY1lTk53L6gLrdy
MrPVF0Do9r8m/hsqc2moS0AV8gNFuVPwY917e9ZbP289d1I9YDnRFm6yUF3LAxtV3pnqPQ0HRG/M
5lNXSo+hiG6Gv6aFNgrzqHgQLn/vhJvO5rU6KDfdNECoYcJPEVnnFEEx1vnIQVUsWLVQOfisZUYO
0NblwYVCZu6jqtKRSYtgfNnflCnSPlMSvsrTZ6Wtfdnpz7XK2zRGbBoV2EwevexYYNfGaQyFv/nD
DczDc7rrzmandGOdqOPQEKltM0A87tbQK9W+Bw6dcZMUw0EwTKABGXrJKo/AKmWCSV7GfZPmm2WY
QNjyB8DibzYMAcPuQiT43Vn6kyLEcniJTCD/fpvz8QboZai4ZTqgDJm4+SIta/6VstHmw1FQqvSy
2/S5n4z5GKx/S0BrQ0+eK23d7ZgHiDYMPUShv8kQa1q6ir6GGt7zvDnVyGjI0K3MjJH5HEC4SFZV
MWyaLUXdmoyR0nkdZTQl6CpCkPfFqsWeFO95bslnck/XAPmjhIMbdkZjUD26rx8nAkvGViTBClY9
6rfB35VrVxc2878xkqDVx5guWdU+h5/9ws0WIwODSDP1kyMCOFV1r7YqlVvGVOdrmAv4pUFJAJMi
Dut1uD4eaZqfLuZoGn1wcbPdGHrLznw4HPZk7oWTcJpffScmhAVJs/15Q0fb+4fGFJn6uHf7pxcK
+eGn3baGVPyFjyueT7HDF4E=
`pragma protect end_protected
