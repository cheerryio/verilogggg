`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22208)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpIZ7Jv1l9IiZKpSiZkp3Lb77OsvZ/DQYlFXChAWnIqEBqnblrZi8wQ3RE
vjfgmdYRKUXJDB9HwPTxCtnO0AclCH2/5BONP/IxO0W2Qz8QYoyyb3S4teAexWbMiuJemnp4LoGp
PYtgYJcx+ttu4rMiRdtJ9ZjY0mNiH/CHUeaNqEFBZmaR7atNL8RYbrOGNHH2JiFLn05NolGgjx9Z
Jry5a5wEzojTtqoFgoVFTujg1xUxhBgsUWEiNPfvikYsGV8XB79gKTEXvULF+WQS2y/m/3AveuIl
WWnBOCKP56YxjQaKHhytthNlpS6ZLLOgMVsZ9pfcQrcIq6IWrHH5moLdcApIukYmFz4/8BZ44oE7
ukLUUnTSV0pTlgMaN171q8XlBWwYMbSG3KLNgGARZhK+XIn1bBdhpGkIKqSYz9zrrYrJF5SwJbjd
rEkOgAR2xfGTdiV8MMnDXUu7JpUSmJPgVQQJRCYfGKkSlbc3+cQJX9BQa0AdkVXb2/uAovCKnKpZ
D/JoVE0FvXLJTc1egRmyw05Zm/JzlSme0Cy4/F+W1f765xD67WPjGaNacqoios3ckoe2gnkNmNmS
fHEFcV2mfSKSEEMmLrZ9MCUWiBEFrglMbB0kGZvs8tQBFH5b/r6j1X8ImIJAJpR7ATfZ8MToZlx9
w0pTqK9bmoBpaDZHWVmaQ4ZRUBZ+GlE7mxMWaX6/jLUgh0zReghvmLJl4JrbbBSXFMEMTHM3I3Hk
RtudpbaZgJy/q8FbBd7Mwke9Voj037C0CH6tTjtHuX3ylAQt6jDOSC5zLZIoqeJZ7X+6GBt7AttY
VdOIHpUwZeQpUPSR7EQN+zeSofQIQDtZmef3OPYuhC4IFPsxPTmtSMBohQ8ao+2Nk6WYjcMVL4zU
vfGP/HQRCBzUIloz224mc6Yo0+jjv8+0Df0Et/5Y6cTLkOEzHRZI+4srAZwyiOAlNYOXYYS2U3WU
gRMmpkeRYPdEuQV+ywghhpmjEE1CtYhj8R7Wxb0ymFFON8XXHLIuDxUxfeZl8qfSNRM4F5QUdwB7
bTZNHAKJrYcj1iM5ew76JZkd6tc3UVnh0ZmP9UfAnUnj7umEjeu0Evkq778JvoLcAubgyVk1DtyM
AvDb6pZB/mfUEyqHhP4gH+5Y7ne3FyDQYPaF/A9b6SWVJY+peLoAZg7XhbTuqXNwGfYeHml5Zrv7
J5Qks3VcEAnKTz32CYljyGMkZH6MXkwnPkB6zLAk7vBOfoim/AvacCzxwWIrswuWMfW6jR6gpnHl
AaZbOOzqzGU0MLuF7DW+uzIKNV+kGPIFnjfwXCz4/7efrSYOJfc1vsj/jaD3atsscOoCntD/GehY
JWimpTUGNB0LfoFLEbbHIWe/2PRlAeXxPXfaS57Fcn6e6SwWEuPC8VZ37YIkzysnYW0YWS/B97tW
Ud7jITkeIMyAv4eQekAnvAEQbjCeR7EvbB1DHLpIZrm5nJy/NhUMGp/bH4+9ecwe3ASu+qN9fIbJ
OtRvs2KhhXgkghTrZAjAH56eqo6JT/giYZuejZre8r57dsB2eYEvddKM3qSafYxK0gjp3TqMSIu9
kBsZgwWCk8McspLxkUoBbEBszVLpicZtH2rqezaORi171vJCHFlW704EiYwdCBGd74+/WY+jVE0N
IR2Zgajg0x3TdJEj++x+glwEGZy89rfKnUhatyCAQYZdn3YR/xbssrTj9h3IVm4ZQCVo2zlkNV2L
kneULzf2JN7zAGAhxRyF/70kPianlo0z4DjHBf2qZ9/tJqtSoKgtflfANkXONp+fHdi9nrl2BBzI
5f4baUuTq3NxvMRxHzzXeSHnNr4HJQEhAnhLCLkB0zMuvUdaIZLg7N9Eoeibnjxh5drkrSWtujr/
QObClFigGoLifvu/AmLDIoigNbF7cN2fNGjwrgfSqBLAQFoJTAJnjHKw0PpNUcGarbwpMXPHjnbe
x7F5t6uXR9pUqtme6XOHtouOlb90tNXp93H775kFA6BVIlYAO7XBjgh4GwLBkBT/W/HpUJDkcZeG
SdKVl4URCC1EB/t4grLSpYnK1S43WDDD3QNVl023JjiekL/rkjam5AtTI8HpkcxPvzGz/xdG2gi5
i+wceyHodMlbH1/9zOR2PwMUzFVaEW/4kl94oS5WA8rBCyXijTvJxAXml7IbynlSBtb9o6JthKAV
DTDEJPw1QSXXtik/glkrzo45pS7MX8aBj6pNrpjYSP4xKql/mVqzQeTCW2gV2kXc/Q51Ji8mpNN4
Jnb3daaInMRy1gZnexNrwfnSX36UYPiIYYz+VePlhHKidgarhc3uqWhYPQfcEmPks9qMLAImz9P4
K94iSwkKWxgMUuacdWVoXR0SbBGvTCnkN3zH0oB6kRtfuOeY/fEnhbWsZSTueAEoQGyj7ASycXby
XLqZApdZdJleuBsG5WJFAuOq/nvonTTp5BX5Lufnxz5hj50VpHjohGsSki9tZc0nbiOWlhJAS2Ld
k0NzBPiFg1j88YbGJIsHVf8NG/TIQr8B88qJzXBNhv30nEvcEYIHEXKhnu+3PjbA3QQzpn/kUwsH
3CemNmXL3cdDb4SjJO9ImGpmvXF1MnQWS0xZrE1B67unvX+QI9K6Vwo3zjRwHx4RGPUVC/50mkqJ
aT37xOzwr76RPwhptguIQW7Hei5l5LUd+Zgu2LLn19rayhI7YoRH0pqxL22Q9DDeiaAQyvslyUTX
/o75d1bIIvokQIYtUDaEFru1xv4kfE7gTOdKNWoiEOHvugQrAbBckeox3UPDxMmC8E9Rl95AHvH3
sM5XxWcJqyukoktdj2GF6OuRggl8feZPybYgtcgEGyWrtDo7xnjPIG+oozL3px4Qx4spNvpSwkFn
KaJz72BUM7rWx5yy3Ppuo6oHQICjT8jVilDxBMJ96jkJdNV5S/bwuz4PqczL3dTww7oRHv5ia61P
9m3bpQcaCtuyLxparh+wx4syYMISg+r1WZfFDdjXGVF1PoL9SX5s35nUyIha8zTtPmxIZTq9DsBP
khRAvGD84XEj0rihJ4rG59sjSlP/4+MXjvKGKZnKgopLjjpIycXJd/v55kUbjA10QeMmiURCOzjn
lwHGgLeCtzYzuRw9Bs0x0lIWWgDpT0y4/yCMgwwj9l7UmkKs4vmYyHoO1D2WvQEoHtxSo+fSX7lE
wxfBP5Rp8uGRR8TnHNvqu0OFC/veI+4rgenoTyfmq697qvimedOL/o+azbco/of8mLzkFpKxglam
QTls2mT7XehyM1mZz7Uxgr2JfWYyKblxK6CuBpOENrK/x/ldoog3aR6ECIo7IP16pcChFgQZkCaO
BeCqhapem7pQANu8+l6QBFJYcFmv6gjC7O/a3GLJ+Rssezq3DCAA7DfUjrrn+c8thBiKdm4MUfil
h44MiQHW7a/DVdypH/G2lB0OiTCy6j5mmWtK7idG+NLA9A1gkz8+PMLCrd1GnBrwXVhqX6KF3VoS
AakuEfwOMwKH2nBY6HmTp1vB1dF9OMYb+V7Czm7WVS6/p3u4wG25gNp6YhrZU/5D3hzZs2Ij1loh
ae0oEWYRrsvARdaQMWkQgK2LHMb9xwxLVbwA8lR/ufUyA3A62bYdfjlJhZB/5Cr5EhGnsyg6gAEl
jO+6I2xFRttuJhRodNY5QF2zHZIvd6XJ48csFKLrxDLgQ4Nxii1YQq0zG9W4DY/sfy/rDyQ0Hffv
dCbSXwl/4G7IeaDklDpJI9PscvjlN0VlFj5DfaC0Tcep1CNjnm0dSiVcpaTO/gyTJau3n/81eH6h
ydE4ir5THOUCBITa5wDOOuuySvcpvZjgUDTtMNt92OLP2JKzrXLFN2vRoGrBjL3fhjNy52ui6ioV
bWLmLZAFnX0oxWfHgnPKdY3vFOjx0R9DR/XuyBbGIdRW1NaEx584tkjQ8mR8SSsSKihPjK5FbZtK
B/M+XnEDz8fP7CvDF7AHN+CPTFo2lqUFzSL2Sd0M+hugRNXD+j7j1TK1/A2WZoUPcS5iTmuIgMfo
JB85pUAIwXeEgV4j8lp6wD6S6b+Al6P1Sb4tN+xmKWScOpQJBP1/ifme64m7x2QkYrTfRLaLJSYY
Ff7JqZyCAT6LZEECtUeW8my9lY1JcqZej4dIFAxv6SIU4ELLS4rVYHzM0iSPqOMEqLq/BL79mwLK
lMSj1oa6VlGrq+NXmGY1tPg7QQVS36NZAyZx5ddRUGbOhEJuHFmXfYorFwqmr9q4/d1RqwbTwQuN
AatHAG7g3n7tDsaIRm7cdo6x+l6CCDmsSakvO0oM5zksX+ny+ZmBJqgAAwzcwvhAXlvCKQVTSUa0
ecpCN4wwpxFftYncWS8MZ8fBheaoVgpTKkjQ/DtbZrlUmJcVvAHvbCjBfre573x1x/rX4D1c+Jfk
FruXS2Br5mYMJLKyC0R49kEQv5Y7YL82bkIxYdAmVyV9AKqFvz8yX52Z6Yz8AWMB+C4ycq5N+CBN
LDgEYyDqZH0SaxJ+3wyOkpRQd7sHT8frPOrPfMZmRfkTqNprly0DNxR0n8wDVwPM28FVStskR6Tw
wEfD1yHLQ2GZTEoSa90gOxBRXBl/5VamMDBSBqzG4LY2sTz8Y/doKP/Cocogp7Xl/xkrrGASIZms
uOZHjOfFqUIdy+tnL0Pb7dNPTw9usHKdENDaUdn4LQNKtxHKfoGaI3QrnvaxvychosceN/LF1qaq
/ST6fE7V0J3ftDr6p8mAqWiYouyzG8RrQGJKvIcoBV3bxJZFlT6mXPTM7DJEvULStiTGfdpmlvDJ
Y/58hRGryOl9xg4U0ufTt+EV/J44ULeXqEvaARM24uMcVD3p9xlH0eGM0qEfvasA4uitYx0gjF53
xXD5XswlRu5OylcnoenePVMvDKXT+h3435ZIErjoLb74HnNcoXP1xJExQMVwwvtcOSpshOYjgbqs
n7WNvQvqiMU+iyzV35Ka/ljsBKjb0XjyDCS1eUfGYtEnZYduqHtiEj5DIQ2TBgdl+epCw0AXmaK/
ghMvffyXCvF/wBjmUrUXFeEu4CXEWN2ig644YgPmPimCQvY15ROZwZi881aUSO5LLKgeO67XkjoF
ZfT6i66pSYHSZRaEWleFPQ+CuPQMcLD+HP28YISiQLj1FNk7yPfDkpQReyhssIVuLQpvDV793Ykf
Okmj41Qck0Pvem3+6W7ep4xlwZcfGCVuvIXnPRfA31MI9D0qP0PDhLUDQlhrCj15zEHsxKiGpGKY
UwOs3NSrT6EexAXxNFfrF91+liRyMugyHC64TqddIkHdVBuACR/V8DNUwP0v2lvWWCAvOL+zLuVN
lZENYNi6zOgndmIi6KRm6xEzAquvbitKjcbIgVQ1HVDitf94uR2PkgLTMoHSS4gA+o+ttKkFyE6v
LoGt0hiZR6B/7xifmNLw05xsx5c5esuRPe6XqjBzpZXCqGjGlkUUeqEThRUr7Fk9BisT/aJr5/xJ
dEZDqy+eKq8JKVjeCBAJQkmV3FxiifSnuyosL4EwVmyG96yg8UsEvhFH2JTtDEf39bX2gljhh9Zw
m74yR5Uh4M7G/oZ8dmYL0Y97xIrTrYQRUDMT+DR2yfiisfRPncIoraatJ/bPGUCWECtEG0+8TnDD
oOQs8UttR1MdcPb3O3ZOp99NsZ5+AVXhm+i4h2mnqVWVbzlQlhW3N6nMX0xfdATJcs0d2U11i0Kb
gH2AY4eBwIe/ox3C4rHFff5NKtvNcLJwDW+9sk++8ouMOt59uzpUX7xdC7yWCP2ybXj8f0YI2AhM
3/io/Uxu0DnDn81i0igHP6JiG+vUeGReIjo041boVohd9Hvn0CdDQy8EqSOX+AtoaHWn8yUJZ95T
K25/ITX1A1hBg4WQ3n5C4QROGUjK3Bg2PGck6SdFLMUxIA0i93KEfg/dc/7bKdgEkU3M/Y//Gi6M
lSlOJ2nQ0b6jkJPT+0USFVglBRK56+Y1Tl0PHYLTgYbkvw21OiNWOOEt/8JdcH4Ozr8lXleMLyRr
DG2jwLU/kWfQEcfOJ2YTayx0rokIXaVw0QeLZzNgFkd1b7XsSX5naqxPJHKb8El1Z8z5p5PyBARM
4yv5E6CoshjpC7haqIrvPhyKs3UzKRmYK4dabZEN6bvauy4iYPC/xmK8DaZ44dHiMteBheUmCZFE
J7GY5w8Q5mI0bJQ1QtoP3qNpk6jZYln38rXYEIpoZZbdxVvAu5GRfwTLWm0uYhwJZ7XOfQDvvti2
kYx1XlspS9bFFGv7xAwWUpIFPcw7vX+U03YsQ7CKuariQ3bEM38aWlCaiibl3kxbYkheArRXoge+
JpvJvs+Gwonc6IO4SUoEaeLyRJPPLKoAVy2XyTEdsj4/xF2wIJ2fQ57p4H+tzGfsbKfjAetet2Cl
EjASqoPXF5JzP3AV3hCPDAVSOTNV5atkerdsXvcpQ1921wLZEUQ0xgJ4yR2fi58/DMAi6nKcCHel
zteRyi5dy7rvKYSNlqMgSo+jdoc90qFZXOX5VBeaEuHloemY9k2Z2v4P/38BBjQTVC0mtgJffpHi
phuShB8LIO+RteW/Y1vrlTBphDi2i0H6HVS3sxHHo83j6ypPgJTfJFzr+ulqu/S5PJMpMK08wSvm
2nimRvNIol/KqNVO5rSIP2FEqZiHTf3k/bX0tmOs/KT1ZAigGB2DiXpFLzmYSyUmjL1usujmNFOi
26ZnIyIYKgYdX5/z7AjkH2yPw/Chhc8FxJHCA1XTaOH8pqMTvJZTdn+7gbsq5A7Q9WJzfvqFq4UX
VTgN6wqg527xZzAA3YWfUb7JMMY5uhzigh/T9OSUCrepWESArrTrLyhxWTpltRd2Yue+mVOZp9+F
KlywP1iNCNAqROCQ1uBPaWCr71qRYz2/i9/bn0wHd+AcbgU5YdEkUQXr6QM5y2/Ptnf9gBzxKAA7
Dhhv/VycTxIHWJ4HMZBaBJSGJMsAxL9IWfOI3YzfqWtd+EzOdohyNKURxE7CvfBxYBlIHof4Mm/V
6N6jCkkP6Bj2cdFvX80vbNTxKZJmsBwv7iWz9RWx3WLdg7KlJc0y3SpSiCJClpQ28Tet3Nc3Bfy5
NHylB0jo365/JOTBUkt7+BTc1mAW0Vuhi84doaznaikBLgbX15dsKFl5pRAZZ9koLzYAPFNeUs1Y
xf7LC8JV02qTOR9ndr4qycx81pqLwltbnOSDjG9C1HORbVhGwc+lyb2viKGLgKRwrSZiwr2q3ork
ato+kGnGvYg5veCnMdhE/mFkTBrVzsI9XCkJiz32tQKvDnRXSykGAp9HnHCQ1qRNQKKMbZCUJWD2
7yzYgRS8KDwZ2faLQN6N8lLfFIo/gvH6qOji77B8aU4McZvJC76gxKEjP1PJWW5OiIvQmqW1mgre
QLkqMf79tspoGhXMd3GXtyQg0JKQ64qgS2Mkd5kWRrvAz0XnoaL8AGUD4msakUUEq+zioNmcPw2K
+9ohdFkOq0QfPu5PDtPnwFWNlCI4Ga2W4vjhZQ8bwwu83RtRmo1QVt6rr4BppPl4ZiuiHD9jrmKh
g8GxcyBftYx3PFt3duSCO9GNd4A0/ZP7xfa2R6O7LNFQVhge9XyztvptXOSt8vzgNELrFSlpEwp+
a6OzTquZFBEE370/mwrFfhoM+H751l+aJ64VxNmT5Vsx4m7sCGukJFvVrl8upN5yxjKxrgl8IErU
+CWm92Wy0xL6QLmo9lc89U/k8HsB0uviViUOFrMSSye1bLzZ7+eH9q8PHCHdJC8IJ87cT06HQE/4
hmgTKKnVeJ3zFNjJjGsyiEsF/SA88DRqB3iv6j7YCHchgL+M8WA7yufa4Uj965zR+oyxU76SLiCL
9r3kRGzo16HiC6B4Zs5ZeFgndYCERDs5ogLB5IB6ZaXZYGbo58gPezRP+O1subvyRNtfyyMybITO
0ffroD8VlBQcojRvxAvIxywuRIb763ijzUb4GudaRP/nDAjTzo2ABPDLnYM4fD6P901xR1kkH6cO
4PwAOnbP12IxVHOF/Owggop4sE0rAI8czEwQFTxeXIRAZz9cC5UtyJY6vAlzpRf2XNDCT9l6FPJa
ElRcxlWy4rO3GN7VtwqpyAin5I+zn3aGSg2/ZSOGvsRycMU6pyJ3WZbtCYQqAwzpC2PcUUmfUSIa
4oDcJyFzc70CoouEM3mnCSQXGisTqpq4/pIQPr1145EDP395DStFsm4meKWoEpBkfAzX2pOX2hpX
9vRtixaOaf0cDBdRl95aXg6KROk6D7PdxAYhPdI079YVO6nNTkrZw6N+0GgH87uXJG+cwbyPTHh9
M9einlkVOggDEspcOfmZHzGDIBqkTgnqVijsZ/h+PcYvoByl9fDq6CGAB9nmWvSOeLJcG8hXSSGu
iuUyGfWW6LQ2eltFOhdsNvGNzm+mAWcJbDFe69gXuO7wIEGjLisCr2Nb1ztpQgVPmZjM1OY4Ykke
mSv6WIczmzK9VplvfkZfHD1zHku2F7DsKJAeHDkWDWAsgHeLKDDpPBaltUoBtpGllqjxgWpNmzx1
SUJnvn6VKADL65Jn5TP9MesfA+UwQZwd55loQh9kNl8LOrSp//5QBuTQ+B+QixFptQer4BK2keWT
ROG1qHOuopdEZAjZeieJa4dBHQdIMOjSXp7wrW5+WyygPxeepownmQsR0Cc5U+5UV9PrpYArAPui
dSX+/SYubO4aNVsDQv87TmUpqlcAUmkEglYtGS6c+PUuYqlC+bIYNyRTbZ9LG3KAIn7RBTkHqmwJ
kE6vp5QOkExDG8p6O8h4LwtlUOo03iR1/ccVW1IlBzv3KKDF1zFbsrLXnF+vmY1NuAoXJECitVE1
mgYJ4w0yxQVJvnwGOZUMikJoyFCWDgxOJqxisaT2banf1uHTMD5+t9aL7Lgm1ftzrqVFBGNcJ3AA
KtC0mTG15ZLqEZfJdbxfwySXdKzrgcO9TnfugOs9efaXNRTPoF/FNVIKS4DvhYiU1bJeMONhLYMr
VTBce5hNq5BQAHGczppiFfxlFpUeBk5HDPHiRgLTlanCxIp5NH8yH9U1DreOQ7xtglUTwF2l4dq+
J90KXPAimnqphgXoBA6saP8ZG/k4YiwH/d+IFlruxX8a2qiZXd0rRcf1+MgfuNuLU28RsrbkqbxM
gJ9dNoYGeXvraWFAz12o2uP3oPyZvFSBXo7ICnWQMh2SppJhrJF7EyFsgk+QyVl+DVif3ALgEO4p
XryTcIFPTbmK0n40NkKu3iACoQ15lWeTP1NSvZOkzdggoc++anHK+SGBA5kf4Kv+EH5rVbSL1l8E
ysxGp87Wbw+1xqWPHME/FF4mL7fU7jnWEA5twL5/nJM+m+8VVmdPTbLuZC8veNOFCo/+XZu2sPgp
WJge9yuauNRcJq/YQTGTh6hxQc1AzptUTjrYb++RTJj475gZcgLXMUk6avynF1Vee1y9/Q6SthfQ
1+GuVqqbRyQR3zwLSdx9R0RrrScEoLeCnKx7MhuiwlYNvoN3UIZkAZ/3M3yfmKD5NUiktTtO8JD4
kkyCMCRP2+WxfXWXGiBsnammVICByGTbTUTOwftvG/NKFFE5Jgz6GWBUXDEvdvkiv0R494RksdZT
DnMe4ZbtFVcBCSn1FVzG+KrHv94//Rm76bSd7I/2n/dZdegAQzhyD/aO6ehYHcuT2KKVm0C4J/GI
wXTisjiyQGw3IUvnkOQG/QNbrK9AAxvCnpzC6xKGGApxGsbCcxwWJkp9mhA/1yDd1DqK7XGBQi9R
lvS42pRAfXb9OS+5XTXTSmqiTl8KgeEcQv42kdBt6bwvB20JNPfIktoPiELopJ9iK7TXe8TmLN6B
kEZkPHkjgl5iCUnWV1HwGx859k91clRYn9ErdJ8u/Zm/4BM561wvBMqWxoDPTj0HZvFOyRAHkgrR
SYrqDxyZZb4c7k4k68YsPN81kslP92MJAaIyusXwoBwGuiD7tVeZVdCJzc7IU6C4W1sLn9yzPCXM
9Islue1ozGLaDVU0M0XEiJ8jVai/QzGi8Yl762kXU+zntOsk7Y5DCYZeQp0iEhrVh++G2ryvSsFk
EMhwfVXO0yYRPuh/qNaOATd1AKSAo4iFKbnhyM7WedKK3ZIDvYbXlO2t+tJRTJCZym8HECp42DJz
OpDR7c//IH9p0oLYlYJFk/s1WEn01QKywm4dulCKxzwCwBx0OCTx1TPjk+mLx9tCwTZkXP4O2COY
JZyGaaJ1K8Et5Rm6ZByMTJz574+USHKEaghUgTIIxAXikZClPfD7UmnC3kJTOFPFpDAvq3IHDslw
FxOPC1A2Djak4tPP9m0/56xAeGiz232mDRAtwD7IY4PeVXsPTbnKM7nPFj4WuEiCted5VnXurOQL
6DuTL3YUUkGCeU8B7o/221Cbsj6kqm/HIKzOFBXNFggN6ehNPQ4SWd8W/w2sj9aK5Jr9LxgN4e7j
2GbKOy0ETAvCE2KhF/RIhZZFAjVm5kL1h3BNPNgC/i0eIywkuCIYHG1sTW4RSSGTh79b7f07Vg7J
3F7ZIlgCm1JwGOFZdv//0ToZUNWMGt23+IyhlfuUSVs7//idd+grg9P/TIfT3nbcXuh46Aa2grAU
67gv+hD0LD0Y+iw318uhlHlOY/5teVeIFzcp7HTASAKnr4OS8WLiOVjlSf7r1SHevhy/4PgUmXn8
i8/Dpyk7ovIk/yZixYaFCJGILxMhSsHbZq75M7frMJ3to84J6vQ6VWKdnJ7Xfx00l6REdHDYcWUl
iuR6xC+1vif3Pw/NN4ECR1ABcsLXnXS6Scw1PlGTa+RIo/1IcWcrfu78z/Sgdjfk0yaDn6TGVDzt
Wk+q0MPWUYASxdHCWGLOSMfSbCIzGSUoDMI4TE7E61cYqndtn/zn3mWptb8uuGWZHMJ7DV1qyfdr
sUc7PD7lAv089rh9HDkOVZnTwEY04ZhPuVt2dVpyJaY+6cKQp7gI29HIcUPN+qEWXF17gYW3BRTy
YpkLwZ8vAJDswHbFuUh0cf9BjlgqPE0zKOpPFfcvGG9fJrkPT3OGdI+C2Md7ae3Xvx+FHFbQK5IR
6iz+mvL4ARIwDtu7u9gm7dbQ7Ek/ZZiz+9ClKQPP6mzcK8T4D5tAi/7N2hmyp11ariI3yY7s2HO8
qCm4P/A63yKaESE71l8Owm0D5XjOzEq9MMx9GjKZUyBb2sqd9n3xWSCRt0MUZeRHpxszeXMlUgjv
n0vllW0rywmaCGQ5w/Vp99VrT9aTNi5lflxSmtp75kFXx5bum1XOwntmBuuC3B4f/OKxZV8Z4j4w
xp6DLROcR/P4+XpJHDA5o4woxEH7yfCEgqiBVvbyNvZ5euWHJAKKKM2WLo37RF4oGKNiW/5CXIpX
ZeiVLebYq3vZgesfp4O2b3SY9T1RhIjanjXqPCmp3p3UPnnzpRa5aOKEu5L3HsR+IIlTBwY23ihU
SUNTNpup4Vte+OV7lZXe2KA+J8Y9SRNzI5RgUDAoO7gdkA0n9GMbcjwiRLwtM8XE7qkFiltrqzGe
NwtsszvKH65OW4yTnXoy1lDnjdjUNNtVavLqPvir4hL2CaCoPIz1creO2JEBcWAE0lk765jC7Ok8
USl6T9kWYWzcpgeNLIIQpNFpZPnFEadVxlnoYT+GRy+yHUxj1cpoDvbtbhvvghv3X0fRhCsiMe+0
UIRvja2qQuD8GcdzLONoowt+8AjJB2X5gfstZerZ3QRyNpuuxg+Xuw+KTlhd+J1AVKv1VPf4q0Ji
BRnk1Nw2ooQJTJ0/B2S07MTtc+++0oV+gsUyv/6EpMH0ckZiFVZnrFlMtWkXrhsc691IZiSymbmY
5hynWqMinKeAYLhZKDI3iaamJYZ3AKMD+J6jGcX/9NXzILf3LI+yJcGTmaB+eLDg/l8Wgc9vOr1k
IACMAGyqeXgINXWhWqSMFLJF5/rb7OmqWpyRxBFqmQFQetgTKRHOtIrKEg7gvyJtdencqcTexYC0
eCmCWCq5VwR2fZpeA3IG5geaksP0VOy7uzfehUgpES/+kvD2yaPohdSP1/z2CYUOShBIGnnYlrfv
ZUNJbna2YPCyZ0LZo9AFGJIrmy7yEZK+bbA1iWzCUH/TwJne94hmbhZhLp+ndyzLYidjTIFBpjQS
vJbyBtljrO0RJF4lUcvNCp2Q/P0+iJn84jG2YxpjdXim+SmnQtPxturCGdIikK5Xh0OqyZMEjrqI
Yc3SiMsvtttRY+JBrn/nQTPRFlFZhxMy+WMn4p9x5WkhlP3iWpyvPQn63tesPU2/yWgUpyv7vF4n
u3yqOaxSJqgJBNPR2m2nET01xNsdvKSbau3LMsZd11GBlCabXzkvCW5jWqtewdob6F4oAoQa+psk
lui9tEeCGT8D+WN9/6k1n+oeQAk2COZqkib1q+XgRjVIlCsVcFalPxtUx8TEcrbxJ4JdVWWVxZi7
0VF2hAt1pN7uot/HVVHzPT9QUwLMWmdvEFPY7Yg8jRx+t4Q2r9NsvXN8565Tk1xoiTsUUy2XcZtP
ZuK9ayor9tjG0A6+2CJlulB+EVSiUB0FvkWGRGQ/oHaEzHG/GOsqdrcD0BdSbjRtaAPYhhpHLS68
C2xutJ2ffE+yKoiIdQIPBMlN5pJAbjA+2zRhA5yMXHgaxub/MuO2iJunRar096N2+oV+w3p1JAoC
m1Q5bV7tADdd7qfxGc96u6+a30/RZpL+KIOg76bnrHAcnAgeALGxSexitCYZY+WQ4aZMHO1//hzU
+7Qk4UWLsXuuW3Ssi+w1KCq0j4CSDzuIvyyN/yRpUgHO6srU9NxtfpR/CwKs8qLZ+or5l3UUR6ol
WNCtNzIRYIZV8EVbwzMCDWJAjQEa24Uocg/BZ/v/l4Z5mX3T4t2FB3jeMRYBAKtqRKh4PSRptAro
7kjjEEJnWdpufmPqTuNBPt6SSmhJjDudEHHgXh5EyXvbnsQFa0xo/MUnzE0TrSYgmCaFH7OlPIFy
G4WUGQhfqfRiPf8kpN34FQJXINj6Hh3T58ITaCqIdwnCPKt+fdMkMtfRILy0/cgc/Wlpi/lIyGIB
IhXBtIrHvfWodqsIMQ2wI5lQ4wwjDb9DKijuwHjiKviELPVMeN0AGC4V2WJAH6tYo2Fl2P5iD7dn
BjQbaERiBfHitFqGlu6XD4+/1Movi4b3ppqUf91NGFELRpR43Osk3L0Us/rhbwpRPR3H66KsOuwv
7IXuLsTWbLUTecvz36ismNzaDAf32aKW/ql2Qt9ekjnmJk8SKAihOg4UTbjNhLpIa+UlGX804hFV
169Kddm4ckG5zEDKgQwdoiLfoZpyMiu/vdBl3ynKY+qwzQYfMCYSZakR/AoSoTXngn7tzOgpcf8w
Eboz50v36th9e5ej5QTfviArtI6V11Wf7QeeAVgUo2obvpguItTLp1MmCk4qWyXN+SWiw1LRI3pY
jw3wVm0dYEj3L2vENUW8lEcy3iaJxsS+Dgxm4a//XBVS3qI/JjfLuRecZkWKUT0o8Q+p0f+Jt6dS
OKwgrj/0HEiEJphxQCvJzkimAWSvD9VojOpecdVl9GZtrhHcow1CFqucPOuv0ZykGAjp1S14ZY92
bNt68+gYOu00KuquEZ7PwH2Od2bfQWYFgDNF0kJZwv2+/RBem0Pfzx7VMFp1Y0UGTf4Rdp6As+EM
j9A5691YnqzirLiL2CFWayExW87ndXWP0wLfdPUBI7Asr78EpyWwz5+rzwMjNJOQ4Vn07gBEYQGJ
5uy14c7Vbe72UsdOzVidjHtoj0lS1zG/0ygxUVzhlbBu+06HOgIUq7MIEquKX0n8NKCogen/ez13
yTT6MJDhbmt9yDtS1MTmRccqLroCyCizha3mDQkMVFy/X8rLoqknK0Hind3pZ1vSsbO9xJ1pUjnH
bCISYMFhpJUblKK1g6434/+bFq+a2411Qrp5PmWAL7D+DWNqFWr9d6xc7e3c3GDJAtAvy1uRifvZ
ZJGu++1pRB5obJDLTTcisZLZF6n3YrjxrrxDCI/w47ufFb9KnpJw2cPx7sqIWjQrtYqPTJgDst5v
8QYrFiavGxUFe+zlL7x6NpXr5ld+OqtvjWzsy9wPVT+gn0Hs2v6V2jwoQNa4OSYV9BjUyxdKQsJZ
QQVb4wmlV7u542c/kRDV/F+RX5rCfQIFFcQ3+YcvzeD/1qWk0C3GkV4mexhg/LtdsA+vQk0FCdji
+i0pGfJ88RMnsHaSS/bG84OdVcvj4l7oec8rO/yCRsu86HrxiLVbbkA+PMUhCK9pitvYA6Ub3Ijc
qg7SJWxaSIo/G8qV7HJwKSH9VVL/N/WHdMmUMhgiLSEJczHxQkSxEzvYKxCSengu0JNFdY6DLvha
JFtCpF50KgW/lfN1kSd2OzA1vIpkqWmjBpvxO9MnvycjC5CY/k0N5Y7Y3Sw2evdqU4wNGVNSKYOx
usu/Qx6OuASbMQ2P/8EtzML4tRpZwTmDJaZLYAz5yhg+WxP/ct0sCi3KM6bDy22xuljCUjt74wZz
aZJRbL1sKjK78t0Xxdz9V3/aUxooNP9pu7uus7TtECTEvKVydCDZfyfWpu9jWxmm6b3to3dZUHA9
4GtUHehSOYbmQQEHyJKkwiFZppFLPx2SO/IUjcpXQVS5wRbWoxGhxqI6wFTufMKXRlDHuEfQ53NP
2pxP64MW1Cj20AzvMRK+b83O5AdUY1lrnZaUhWp/Crc5re82FHC6quufaJOCIU8PGknO5RKSkHUL
7KuX8vgbujTuIJTY7jlvyBTAjchgwM5Y2U+NjdwG02+AJz1GaFxbVnZrFNSjbTpNWuFIlKdajhZM
kgOwucMKlD+aSMlCzAaBRDl/dSOu+qt4knUVLIPdf8/5NMv3Da9MjsR2dFRHospF97ZcteVgdml3
Q+028tsqFlNPxxS+Wed8VEahnPU0wHarEoAiiuBsWKuzZppJiy18xwYhrnYEtFWzSsMsLjUtm0Bu
ih6OlbGGjltL/CYXc9Dsvt+ofTdUs1pgduo+M+Jv0jERf8SIfzqy7KfnF0zxi+I5hcm3EwDOOe/D
nqgkwQW6o/4Kpx1F8eZCOl2UO0RJbs1KSpFp/m7KjS8NM200PltpRqQOU7pC5HAnBE3EP0BI3CcI
EXIlsL6sQsvCtHqcLJ51Q8XXMiYy4Gx2J66UeXHeJXYQr7CA/A0I2/WQcoFGiDvxxKL5enq7s0sO
gQW+eeiF+IH9rRrpGLmUtHucdgJQFK+NrjzR9dsuFyeytfNDlG1pDIVJosq9KreVkAJjWd3rK93V
X4ZDlQ1FK3sro2tmKGeBNDNndJWrjJHo1JVUj+2jdyXsIKe03wdOr7fnq4LQ8JwlCglJYCdp5chk
3Pf+EQcBI2u7pQlUjav8Sq/gnbMTrgVeKIN540/MybTpjoOBP2iogp+NwHKHWJbqB0JjEhkl3CSY
LzuVWW6FcrWIC+r3YUhHWcKujfOf8EvpAzsl/nhl4L+MTRPYA3tjeAwCytg8nxjSeXGWrsTmE+uv
xeWb6xVtyeRdaX/mWIuz0w3p+O+XV//m9Kow8uxgMpsdI+BHxKyzei3GUyWLz0DVyUpkxqPr75jY
R5bmbcauObHElfIOrpsKWsoDBd/QLTVntsfnpJ4/92mMN7Ym8wdAuXw4Ai48D0lTETNlF6ON1TsE
LG8QqeXuWCHk7PtSkihuokQ80Dt4H5jZxmMv3dtZbajE0kG0gHsH2wuc79C+kBDN6vwLjbKtqRR6
jRXFwj5jjEoqBEMUUMRcqpnADQ4yVUee4nu9JtNzREO+vD/CEDUDhSCE4Feea5pAIE8+pk0aFy54
+z2GxDD7GNuwYzDDEo1pole3FnGfz09nezE06fakHO+95fqC3bx7OLrT9nt8qcZTO1JXI+FSVOJT
Ick54FzP3k08whlRk9EiPtDpKgo3dT2xiWdTvBUMhUVQEzayoBYfUfXdkY8j1mar8yOCsnrPicQU
hDpwcb694es2sI/sWka0vnpyc0xGBvnj3l1HpfTAOaOAND95ntls4HNwURurp5x8CYMqKL7LUzSH
QGe4+hToGPDx7cyDkORKYtFskK1T/kpE++OsL4Qv8r6U69oNcr375AUhZ6dKV83BdLtiDR/A+8fX
4EVhbzVpxcDugcDtzS7bAzyYN2b9JUkS9cCYi3ZdznV20Fy2Wenvajo6OKk3aMgKj3jnfpbttJ/Y
rxDS2iJrYXlYFzR/BqDD46mCrpULlqJ+5luqIrk6ANbDpEDIyq5lE1T5n0ABo2Tfh9oNdhpygY8C
JkbuxCJYF3SQshrZtRZd3+BxHuGVcveoECm+kyDKTGfpKyG8FRBx2+N/m/H/mVhaUKfJ3eXcehUC
fgjAPEK3prFFCrXy0DBBbVs82Ayf5Y/hzzCaN4YsDkmM0BO+m6yExqNIm7/AneREGC173GwlM5HN
SR26PFDfuVFwnaXa1SXxEra7x4nBwez2+TFGGn5pMOwoUDU0oTq7ND1yosqz8fjliLJw0yd34UgO
9laWzh7CTvEZDYaTXdoEooHkcnBmAsgzgxj6vuH0BY1lPzp7mzZxe6RsiUHg/byJ/MIV7zOjq39B
hBZ7XBRQn6Is9x6LWzTPL2Du1GbXf1VbdZ+1YICcoA+Cih7MRiaJJLH688Ie0F5kB+CWeSY6p18s
fems1W+9sM7+fg1ytLpyaMhNpL2riMaemuEVxXSzBw6nr0OSmW84xyItQ98ITiVfW603dELqy6Kj
dVfCY76WdjVpGkT05UxbcDWwORkjVAIk+g/2K71m6uVCK+hy4dqyikeCicz4oeDZHNG5CNvvA3kM
0aD7+m475QGcneibwW/gZyJiiIm4SVdBSQWXO0oMEGkQrFL3btUtQmvzb/cTlOR4fNiJ7ckwuVzI
ugQA5NeqVmG7Ik/uvhWM43dqK3zoqoKmk+hwFMU2kNK8Rg8h3TZk9OVbggku/RVaf/Aw2O9tIcOZ
Na2HonBC1obXgb7E/fehVpWbf/V6Dn36KJS4nVUn2OvFpmS4B814l0TYtx1Rg+D7qGyvGMUn6yKU
rEUMvDUNsQOSP1UAYXyWgVvwLn4+vLyFemO7Yj+F/x70Cq/ItAeGZ3Tp/xtpTw1ZbXcqWHPdfYVv
EVCIHP/rkRW+B3OUymPqJ/J2vRQDlGrqMMdKDS0FuFHtobaWVyRvi9+hN3mllVUB4RCcbwuy5598
G8u/kOMwAGidn5rTFp3vdO5SRJ8P4JLx/WMH9iYT+7zEqAI5Tat5jGJTzEvKuQYWmV46/FZwzmZW
Py3mwKFtiLepnwEIxABdCM2+j18f0fd5+uS9iShBFZV3ooMuGUZYn7tT0fTUqvJ7xInZ7w5u5rJz
0s5JWQBQuFFQCfWpWMUxDq6EmJG6kvhUvTV/aXRvoSjR9Z5yxd4m4z4qeYi0C5xwLiJPiYKnOWvs
j1HNyMJQKz46IaQH+QPFt86bSZRw/CzQg1wX/1DDw3eUZHIXM+nutu7PGXGViZbNGtHujJcE0t5N
bYXVudUY/wFHimtjISSLS/5WHCnkSuPWhPiIME1ROqfaOS+YG9iSIycb5kMcR+qqeafET0WIqMqF
C9GqdwR5dsJnOxrXbiLWl4qIifRkJXfx9YCagYDidXiOc3lEs1S847ssuk1rLQ0+GrFcfzx3B/Vc
a9J+hjVunpZC5l6nJGmpHnBL+FSJ/G2UYpCBtx2vKlPrlBQ/vqISs5kFeen7Pi3CT8GZ0v5bfEz2
IRJdMVH5XWo2cepFdjYP/2HhZFHCLig2V9AXTit/+hw+qFhvfFlVmOrb5cxgcWpyLWJqv/UHPtcV
EhdcCTXuOJcBX5uy5b24yLIVrvbvS/XMpm0O3JT+c+S1gXqcYjlAYn70GnRRLVcWvzmybFrK9w9w
YF4yVfbGonk5QVeZ5KSzHJuYEFzFuydJHOCR36hZydr54F8E7ztgk//+PhS3HwjfLtPQUk/S6GQI
cmoJgKiA7LWmEMp7PDLV6jlombpUxn6i4DhGvakSSAEXyegPpKqcN6+37YCGgukIegKiOo2m7MEN
lZ6brWBTe1FJq9nIaGNGdiWeQAJ+vzFRCcDmILG92wMazD2YThqC9ruUMaKV4e63qgkegeBAt1QU
tLjy+AjNf/mg6tzgmP9t0KABug7maDjQOy3sCQL47b9YZFUlPD1a0sPgfzoXNX2++AkBdvOZoTEy
0o5umwPy7gPp1AYLOKX+sGT9U6KxyxyMDjJFsw1+KteIzU8k6TlXwxlnWmRBgCgjvzNzgl+pv+eq
+kpl2OTrGaU7zv1mX2xsupwVmiwInkxsmNtPLTZreKWa+xnwHnyl9n5PK257OFhSH4N1phKeZMIw
oQL83Pc1fO+rIaIO7YiRADkCvDWevZ2ZWeLlZy6JQRUl/AaIZVu6/B1j+S4hB+VOZwZTaFCbpugK
q+yTsg9zQH5R6KufVxhhK9Qb3G89eNwtPWxCgGsrlfGPDgj+HRQqOvRNteV3EwbSzE/6YXxuju5w
tPwbuX9JHO5fFN1YopLrd6+yyYrqKJfxV32RuAL6AjLXLPhDgyDSs0T5+Rfe/ecLDSZjfEugnZd4
akDC8XlHURsUOoqFiw8CinxWbItIugEJ6Yqt0hzZj/UMYxBWC9HhhMOOIu1peHkRqJGDVCQBLdKe
q+zTTflNhdNFOMjbM2r6zFDMHj5ZrhdlhH3UsiDoPB5+VF2F2K/wgbNHUrURnELRoxyKwFOT52n3
9y1kO1DA3yjE+2//NV7T42L1cTgnUXlSJ/XdqUo1rTgpVgEPl3WUim8+UHB7IDtTnM+uxryy7v3/
FWl1hvXmdZgRTbbSJ8knhnZzQJHK35Cn212CZNJw1VIR5cTaNmlizSCyiyJdZxBcHNCOeaiU4A78
iPl8zVynbBZbTcoACV7u4k0zAECg9r7z8R+Z4JHrYKTWyGrCBlIPvxsVprLWOQL44QId22XeHafz
KxzGXAorcvexuk5fAUe4+yCsT3BL2K4CvKLWn9VAh/creqWl+XLwTdfqMBPwn2zKnGGcNub1bN7A
oGwt8/E+NkydgAsJRHJeGIOVxQylz/aQP6Wwn7HUGtygyQv9mUd8oJJtYkaH9Gh7HTGAEXvWPoMA
kMaxfVzcmVhu08aOu5vaCu+DTLizxItSS8e0QLFYTYbWKXZxqrQ42ZDV/2vf8g+XwT7FnTlYKghK
Jrl3zSXxA8zkzcEX+PwoSb2ety0kH2w++/sO/VN+TQ0bJCFvwi2nM2+BnmRHl9tviYhwZQoAmcJm
rCHtP/aQ3hhI0Q5x2Nsmh7e+00u17Qqi1c7+UExacbjbbf1BDlTRNzXU/DYDT0h04jJKduEFzWDr
pfhbyZq02aPz1PqZTNg2TZm/0ac8t9YOaseXOtnrVJp+DjuU/ZWm1Q2mh6wgZTfXpgJLAwN+ppoW
QTlgYeSjxf064CnOPnlWRinCVjS1CNpqJiwdM8epo0GusiyLml1iyRo3crAa9k2BxC3RuOFmOkXz
gSvkNd2WJwufLy1sMgkVITdz9qaegaQS15iWkVG+TJGr423+l83R7FyYuJVck1zzTqfKaY6e/ZEj
g3wco32SL0W5HtGsYo+T/jhHDkNhpxwtzDLUVW8ShJhUA46ukHiwcGwgS65vH2yxfzB7PlSYvoMm
ztDhQwOd/yzmglqr5/ef9H9x8LuOm1ui0XXLcUAeGo9Wgrso6hwBY6FMKqNfjTHbtkif1afk7PtC
VSR7V4PvgvyDm7Xx8zjO+ZlB4IsXmynWT0cAsZ7SDYDbtwGRugdGw1MiS26MTqU8ipsGx8J3H67Z
VzAcB6S72s/5NUQ99KGcxluXP4k89qSadYkIXh2acbYrjbBJBLXBZ92OXEpdFxBWBUDIQcLSqj8o
BwHKGpJQxxyX2Z5KeaarQJjtrw5ff/KrFFPtOvf/vEwZaw7ffwyWccqT0/9o8MswV4x/64bRGRw8
zqJj2nBPQlTl8Y2G1nXd16lS6H1QcLmXw4RZ9ZLrfCtA2OI0//hUMJ55NuBIIjBBWgIchPoPWvk6
yZhZPgzSELTuV6xOas46NZ4OqVOq6AF0yCd0nA5s+PHzmmtycTKJLojVk/SpQodipaAtHUvdcw5P
rdXTx8iZU3h1TxUPBQ0596jooRnd9g1aPUEH3xvwvdqUvN+YC4ULMqDYZWOM6/fgo1wtExii9VzO
Xpn6dRem4/CACNf0ughzkjQoUsUr1HtFt3f6iFXs6Iq+05mTWHibQBZZ2EAxuA3by7cfYJ7hylvX
uwFwLK9M6gSWorbZOz7o8YWRDhgFbWxyxm45Z/kzM/bJJtA/sUhibxtLsrOAwkQpgeclPMXJw/74
+QzZGtED4UPFD76Yw1K/Ln4zANSfPFJnssVg/hbsl2cwQur4gzDePFBq07ZAdG0jDxsaFKyVhu12
PZxL/XXw6Ct4Arzqp3vDe1vDPpD1yPNotFbNusM0qCjBXdcOHQrH8oR6mJKivuVle18lymF3NPNk
jQQ5tu0X9USFlf4+VdnsOo8tTMJwVkfCKjdEMTPia66yuSRD6N9RIv+i8PDVyq+vKZspXdQt/u8w
Ue89o4F5sCnuOugiV/0gPWVHT5LkSk4DGt1vftE0FK3i0gXotIIbbQvfeYYeIhbqps+Y2rAWq3MF
sEt1yQ39lvS94rgNO+oP2+VjiazTj3OaJnN73IKEVdrG1bqJA0KAFfIa0N/idubZEX9xorl/hGZ0
RL1oiW5Pjkp31OfLZQfTUpxiAIWIspncxqDgTtdC8blenM9WLrA3bINhhCbX2/y/F0sSn33AR5DX
2DUYDKlqap9RQBAVBAUsGZcprz+j0atSdkG8GNW4EAqthdgHOwdN1+ScaikMVKWY7xilIeaw1tOS
Qmt2WP8dsue8Qu6D32m11hNbkVnYrLFQIuuUp/9aDCc33s+4qiq2MuaXatZh4ZtSNq/gG++Hl4Mz
VUxEAt6AImMOteEqf6NWp3tE2k9RO3E+ocqex52quHzPoxqSXxZ9PMdMXGc/4+HFiHIcCiUj5xOX
0tiF/NEUx5qzGWni+zAZ2/yrkRO8HZCw+lkJpEGFh44npA2gkFcZaPExxT8Cz8WRf74kEmg2wgcn
rPOdMl362/43O47nP+oW+J4lOdbNpNBE2ycSV+lenannKaObzp6HPH4TqR74L9RnUCb0U67UL4bo
00JZhSpdDK6Xibj0i0VY6g/Zavop+ABisrSANUI6fL147DW0/htYgcbiYINGzOs09liDutPug0PA
R5FEcp3nuH0wmEuskpb5nxrssVXTKgOZlK/WMfd/aH/+v1teAZhcBBDMbWTDtsg3WVPKlfFUqz6D
rOyZC+VSmpN5CNd8NwE4ErcdPqY1BAGePV3WidJRygcuLaHfq8z3LNWJREGG5ROevjUM614V/mV7
yMY0QFy0fa6pAh48nOTLBzZ3N/bNiEQl/6/QyNhY9MQLs+5nK0PfYRYlru6v6EL6+af7hxsZ9IWp
cwtUJ2BKhUWbnQictHX9aXG61OHZanGAvIodzay+CvBrzvI2R5B/JzQ6YtkwR/hXp5/Cpru91Ntw
uUi/U+c3NMPWhce6S+UjEEedUm7B5Hnb/sQ7M1yGMZmQDwkZnYLB0/VKK3uGWoGatbUVrSj8wWmw
xOzbhdg8l04uOJH6Z5iNGBj8TBWtiS0TMZyZ/vvvDKJqV0sNi0T1yE22A0yIvL0w6Mz5Ff0R85sQ
D9h/x4uv8Lwu2Vr+Vtp6gS53YZ8VpyMilUtbWYuBZ9rZPGmWQ/rr9cgbQ1VIkhUnOAFG3Ds5TFgB
eVYkQfpXA4eErFlUWREcluFan2mY292SY3yYBljl8rKYOnv7LHyr90HBf+bsGZxNgtsVAHBzy8K4
jaOZ7395ZI8cVb87+l4u+dtbFaFa02vXZgWcqnzFEJBimOEi8WbVlfXtpIxJZaTBGGnozt5vEzLL
s0/PxZfewQvFn0U58XZ0gNW3Ig/o7TI9BZXLqsSyzBgSo0kENDhsk7hJK11dSZ3oYaZT3HGfu0E+
z7obT9/X9YhDJJH0++NcyTLA9q6FMwJU9qLq/sC8pSbqxVUXEOK4n8IvCb32XRxz0U1yAaNKLPuP
K/n3A0nYt8QpVnRj1qZkIpP26Vyt5NNQbvb/42hurc5mNULbrB1iLuhbAmJtcIVrlflwJYz34dw9
zFDu+Yx7tpejHGmVDX8jHyJcEK8zadWJxgoibaWFA1jvxJ2+YUMwHpXOSMRZz6uSjEwk3MLWd2/T
G1RKp63em7tedZlsvfDlB0GmdulFtTHwC1oMl0uzRN6cvRUY/DiPHv786nU+QoKAlD9/DeJ/JEwo
xD5qOA+FKk4AlgaFu3VwuDNNohkPltzEnN5LsyYN2MhR5igFuS1noqHBMRVmDUkUmDwyBENJYw1y
7QIG5ijkWtsJzleQ5D3Axk+uXlUXdPwuEMwsMMWJ2AnmOmweYNS8eA3/trLkNjHHrLn6lQBfzl3S
2qsn8jA9D5wOU5yIc1AN/mH64UeVxLUPy2LdA5ModFP5tyvnQVX8xtxFdXdN4U1OqhDUtMaQA5D/
vUXRPoXgUEV1YEjyG7tffAs4NhZEY58jKNpasxHj3t9IrWQ/tejr4iv1SzN/VWjLxNklX8QAijzE
qZWuO2xfInq31alLJq6nt0t3bJ2lWSCCTSrMT6HLp70zJ73RGPCrbgVWBQQYIN99blx5RmrEQbvS
OBbXxVyLcA8vbyL6MgNJ1sCvpyNWoIA1UQ3B7vh6a2sOmHxlB18kHcY9grKZ4xRqoSUmXLo/QAni
SSxrfnvhBCg5CexaDZ87wuNq7CisVFGy7He5qxevUM5Cb8nNPJQwtSfXr8tYrrDRLY8mq4Tcf7R6
SJy0TDxisJbJzrFAslKx/e/JuMheeqmAP9WFzRrWGS7mTqh5pnL4DYly/6u3/8QtUssfHF+LSfpg
ANLVTqfGqXGPIpyEKFJ3sQkX7w5ouStwnFS4ekzzdl0zhiUuN+YIJdQG1t+1qQApVUmayTcyNM0b
W4M9OZ+q3h+b0OEKAhJ8biSNP1PapGJ+NPrGS7S1TKYPlLk+w+VHX6IMT8M4wjXJ6mwhXH2dX35E
o0Dihxc7ixfX2DCHNQB8PXKcVrwkMm9qlQuryz3AjvB6BvvWeDyL0Itwv5BNSPqUnbip0opv79bf
qrGxZVSB9a2S4QS5jWPZP/peYuR4v6P/Ek3s+uKwWBrJ17HwF9pcQekoNcR3+7/LEPpLEgbiH3+y
Q3XlNFiqzVKZsNi37pbZg21V1z0Z5TsP3sTSO2dkrmNngiXlTgcyjPSLtwuK3hIaFpyOQG/YRXb9
hYRnk9bEjtQUHY4RsGNo88tNeQepYF13mN9msEIxgpeTc16NngT7MrYNbjQK/fpD5VGEYNMI9mqE
6XR+6wYE/dXwAovUzDz34PjiySN/c62A6JDtDuh7KTnWovsJ/kH9UcMsV5/dOLzxJBt2qIDsqgfF
ejOR4GwL7Ug3kQRvfLDVf4UtvMZDIdZWHg1eSQ1BcjCb2aOSj89ZWuNMi9RR8yRszQ8BhQ5CBgFR
Q7B7qIlYk9DsphSdofjuW/8bJENcSjND/pZNej+cwZGKe/BCh+5B+DmS8CQRHhVgwEg43mLwm2EC
OHdpam7hqjJNS8KD25SrTvRHLZ63Rql3yEX0YPTiyuduCRUOKZOzrmXQ0sSnZ+7Z5nmtoqlCGFVD
7WQCXFPlSV9H6znesUMG1lNfKShmdBL4V40snqv1Q3P/X0BEOGWpkvm+7CPTAWnzzpAvBfrdUGf3
DqporNI6halzC/RddftxX6VJBRI4kPiZEw9OoL2I5o3r8aPotY1famyqOLHlrGJaWWfN0GMDxUbG
UHds4s0DCrKCWRVIRHEuCffshlIAzBDLjcv32dil0HefOL1ExnfNIFBmH6Msac5wGl2pl+yJQGVz
K97IDuQEvlLlKGRUW3UF74D00wGcc8ms7KJxMHJ/zI0xbfCFd9zaSV6WSUCANNzrgTxJiBKXkUz5
iEam2YTjy5Bcq14jLDoFOgoBnKWFOgE55dD1Q1KIu8Y6Z8bmIKQbZx15YyCjdcW17/fSXifx/eYA
WdnALvaJ32oGSVrk5g2b+1Op+uf1VWuSLLJKsXexxt1/ail91B1gzcC219q5FHXgDAueQvUSvvGK
IfIvzteb7AVxUB49WvnlAwERtrLMhtqcPqIOFWjucqXwPA4mWKnC+TbtSR3d3pST0kuFoAAlPI1N
1kjjVlF4CHWILKuUhGXpRrS63MW1Y9K2Ceg7nNZKENjcHwp0lO3GtwKBNneorZRxcVjDvY9UllFP
zaISU+jLKEUAmb7c/rbL1nrksAHnAWmeQFv6emp7lj2TascoaEv/0Nt7s7aNWwAwp9o1IzGMpwru
IyIMshMGU9dF4da8roOOI6hE7EACBBzvwSK/2BHKTL1dmugWyhbMirdoKJcMz43TcUdf+5mEBgiO
MYhINheeEAnYAoIGTQ9q0lOypWgjSK54HIuPy+LsjWVAJGfnVdf3gFHXgIlbLVswfrBGA/oHW/hH
CQ5mxrbe2R5Udrcf8Ovr0YewZQ64om7Pw+a4vq0k/4aMTvQL/ZbGOON6WyTHhPgmyM4rnxfl38Ae
muxWbxkuGEnd2hMnO1pt4sNAkAnIQpe6PFoRc+r9CEWVx3G3qzvDMwHSZdmVxbmwhtYnwLLHrK1/
xP6MFx/x2xdS8pNUub0P3cKHTP0MTnEvMTNvB8hykTYo5+n08KEpDNoY0+AyV8e0vO3I/cGcJi46
Il4ge709xKeHdJbI7s9BZTH4lE5HWZopjJFTtGdWQ9P4Q4pLNVFmT4WkQIGL/5QaHbthwzV15DGW
vbc+E4CihqIWuhYNnwA04Vsx8V6nwGi8i+NMhGKXs66IgQhwGrxnthMBtNN9ttSTbvrjkzDnrpUX
Cm8cQfcvOtUXNJ0j0u5wp8NeW/7qVShsfa8fYALgbnwcujTrSu0ZtAJX0BjPmqw5m3Z2li5k+uce
GGUO1pvo74u4caLuaLuzH9x8F3O89R0FRB4vFuH8Wi72hiwyTR6Nmh+A6slQELpJyg2bH2sdfN8g
SkuSMwRqCHJC7Ik0mV+CmVv/EuCuzJt1axaWmnxuYYTyCvuUg8v4e0xcn3JscP0Q2vjBuQ6dz7uj
7a3ObbMYBaKS3/xbXADdKYDG0g/B9w82xoFyUz27YXYsH5be4gbLZvXkDv1ouOGp0mFNxCLjJoYe
fWgTijSq8Dmeze4e1uctR/kMLWPn+Q/wkE42y5MdHjwzpCzHnmEdq+jmTX5tNk6FN2ekjsdKPNmv
BpgVpfkv4IgREYQa5nWiwIY7TjWIgfD7MvAElTu2zERu27iTeQPX5Cd6riRNEpJVIHhu1lAj3WQH
kOQgBdVhDQtamIlBoBkMHfAQskDVWmcuipyYoKZ2W6PhaF5Iw9hTy44lgMYLQukkE4C31sJhidez
u+9MVWsa0m2lsLTWQHhNWuR33fnSP3jBJJljGU+YbvdU+LXidqe/rJyCrOcFy6Yc697IP9pSLFUg
5XL8tu3ts3Hy5AbVX8LAKZGk8R6DwEv9DjgcyCpnlzNjz/D2gj81cvFwFNfkSYSufTS3i+ySkiov
E/zFdfAcl+aJKZqhEHXl2XTn4cMAFPxL4s8gb3wCgxRpAS9WIa8z/zpHxr1wAoz7sITX+pmvhJ0l
8jcBLzqu7TLrtZ3Xt53oKr9tAWX9wOYa+AsxSoG8tBJd2xCXb9UGLVuVpaBPvav0ho6gS0Islo2g
EK5OpMnIC5DCoZ9SiFbgl/mH7FRwFgrkyoGAxYjqpndzIUVLMW8wXm43r+7BkurlfvoWoWkmk2zR
1pxE0ecnkRTcjDmvdry5YP5R9HK0cwI+SCHWYnAVjc9EvCkL/aKls+Ud7scHvedLOQJN7YPjY328
u7V7EDh1Qt1FH+2qJpidIC51bUlx0xGCaP+Wpl/BGiUbkamp+8APN/UW71gAWEGlS21VPnWwVmOv
/zeslLsRZVbMK6W/4oJEpedqAF330REPCSlkpI0CPdtObtJt4mTaiWfFTZjmv1k9f9Pfkhr4eYVo
OEtRQDTOTVdsdsh/K5X/sTOEiZg7r0D4aLcRW+3Q1O4LeHi7e3oqHKQauHHz4Sn5LOgoyUmVuJnp
sGxdaHK7DlTZvFVPwKxYx3OO7W6AoamLuzo+I6QQ+WJ3x7ejslHGdgxxdXO/k2c7SANFVJZcm0xi
Pl400QP7lTLXcKlXpUsfj2NT8mr4mplqa/OXjqJJDojGRr8B7niKfiAR9JYhlpzOxNa4AmLOh8RA
YJlyyty3QyUmrBmHnbon0MNjsBKYgUfc7vJgZ2l/K/V0heLgAZU9JFpRJPd10M6D3UVwjVcHoRPM
+1VTQy0T8LzSFe1PRvecUuu4D5mg28WUpupI9XHBcqYG/mvuxmEJPRmomls81rUE5XYGN0qYUrVj
QQvHq2oxREV6/k283j1tPI93DD+ekCl1GCOQHoTeagtpH/YpeiuWlSHKpfWJTCdHFh5OaFfgEWFe
XCrrWJokz37v7+mvL+Nmo71biPrtpsHwiOSPtrkufJzGm9dfJwrQ6m+ZmkTp1oTytL1x3BF3q4Hx
DJxzUsJjz4OY/tpYLZEeYprPelGGoUKK7MORW0PY9blGaoMbPmBEqeF9yzNPWR8vS9oBrTcURz9A
dxF0DYpkFyB1jEInXPvkvNcPGiOKKJMnYfZS75OVMR5fE5jYhPGC+adTi3DEraXFa4qnpvaXuXF/
6B/NzbXlUzuE4peFxzoX4staRZI78ieVRfUtC1XD4svU7pfGVT9AAEqo/zoa1DQpDtI8zxKR6s7+
eQDSO9mE6lV73SM4gll0tPTKW6/F3MyS5yX72Jk9SCIfsNZfNlYpF5pk6uQTabVJDLSXStyrLQay
bmv+2Q58nI12nNfAAQfH/sP4uIIYIqpDGp/4hJDcwYPecYPMSpJvm/xISdJdcEeiWxleaMFKo7j0
QEvt5q2V7TXG5U2AOn7mgyyQh/oqXb7upcdCMNPwafEE/GXVEAhrOYhuMD/rwBq6oYDIy59q+Wzu
m+8qHhrPK1AY34HTKk5oD1Tkw8BVPkg1jvrfrTANFET5jtKO/toqPG8j+xuUlVd6CRboL/eG6/mL
wA0nek12ix35nQhTFZtrYpHzkiDYuJP1K9RBj8NsSP3xLF8sZjAH/vxhNCZJIW0HBsqfWSOsxblM
SGpUjfIo65G2pYtG1jip8PcByRoig9rSglPYAsQzQT63V57L9f66XkXChW0FdatdcU64l2yJqDsr
72ekmDX8qLp8mBr1ZSiQHCnss5zHKO8mfMGBkzWKXsaAUSZtVEqyVJTPNzce5S4Tl9orgo1+CiFb
ctBmOadbSTsyGIeTgWhHPYQ/JoLAokHg/aLDOPLHAR+m2l3MWkQlw9xdGGcsftfftrhxv4VnJ1SP
tfTCgs/IJ1NTORlp6qogK7JZViDch8v6s/of/WR2jBTaFmsCJ8m4R9vc6crYpGKeV049ny1mDx7k
A4JSSRqj/ghmkI+WcO9TdZ/kdnii9yujBx4o1UEKnm+FacEUN2giQJGqe+A1+ywgsLMYRxYxR4Gt
jEra6FpGSzqUfs84B0aDrviQ52SJtObG7ryprW3QEB1+Nmebn1MxXd9EkPdJo3kglmOoP6freHlR
SkuZZO9krqvdYJQxw0Xp5azV0wAMTWuBd7jIyaAxu9fBRzEbAIn2Q4iG3y+xJPdtraQEKdJL70+x
vdKUGWXRhoNsiCiAMv+j7kbthywOqo2jSYZwppf6+LT0XPRU1vskvNgqza9nBq4m6+8i/AKuMbkh
vrEbsof0S//ofBWts1AqDaC/rZRvYm9eHjzndbmKJ4srt+XaQivqRpuwamFeDbvhQ6uxSSri2YuA
z2SlhtZAqG+el7qMGNsnR6h/Z9ejGouLJw4M6WycDH+ouR6yz8jEW3BHOHnGqeql1yETqWNjDF4V
7OnKJFuDKr+iO1KK+HvRiGCyBUE6uGI5aH9QOPtW5HCOdOD04UuyG5bDpF0sEpnhAODXNikvlJFV
+1kWvXO+snkrFsLvl3+JkPhH8pxDe5U7a8Kbs3h4Oa4XlSHCwZe6EXbHA+u8SGa/BPS9DbfO3XSu
LysmrZIvvo/Fk8xh64jI/Ilt+YrS7c04ARbf4WVYgzgpTRxAn2toJtoPlh3ZsH9b3k5qE03QIbok
k+cgyP9H9NiWp8CVQTsAMlXZPQnOj5oDuDLzCbhP+gHA0uFIQ+WlfTeIoo1JclWo/q6Ljx/y+065
tZDig+MlerMNl5uuHIj4f9s6uV96iSSoKFfAbgfeipDFbFya+qJv2UKFMyc0RCA3/n8UrMBrMYKJ
wyGkRCcqrvwClg8RwBl0ipuLTu2xsVGwejYdKikGxhZElojcTr4V2nHK5nTpkavVr/10yEiypSPH
N8eKCXDrnLoiqPggl0Abz0H5hvMIwpt1Kis6XwCoU3F8E8r+STh2/uCX4JUNT1yVKCDTCy5CTo/a
G39d3pOGYdu6OAdr1qJecJiXQgR9uR9sEDMPaEMgE9V3RsUs9fjZIPppDSrvJOLqPOawMKoLXoFN
QHS2FKhR25E7MQQMSSxVsH+pyj1y/mBguAggntQE60+zgl3E/yxhzkIkknsyBDTa7ZuXFV8SBen3
YaBUZrOdKQSu2gbFUXu1LbxAghHdWBJDRpBzsTPg6GoEgrC3ydc8GE9ZjlznScrxhdgUDUgS/Ayq
ZsrQyXHby/QeiiJGwLxl4AwhBJEpnRSFbkgB6hnnlUhwzy2gpAxhPnnlzo4xQWQRlJ2RvSbPHm38
M1qQRzy2tj3gnVlF8srcCjyktblqW72dMg6ONN1cDVu6QsGQ/hxyUrz0kAQeyOspqqGg1sOXFn9P
hgZ+FeeEjHJI9Cid3iiT5eklVeTP58V3kVFXyNl856owvwrVfzVNX0mccB1ztZtOYDeac4iCqis+
o9eVnLTrV0ahisL7fIdnnw9MX/+FkIj0vwEqKBfz9h8HfhpT2VOYGyz/tU9Qi+v+Etrt8K/5AK0q
EL/PLEqyZ/gb0rWIrDq9WXqlmPmcV2oyw1CyVgf4MrAQ1zaJ76NmHmuZnUZ9kWROqptu/j4e22xo
c5pHMFqHQI3tlh6piersFCOEcL24R4okPeh8C6t7bSIONLF6TTQcS4A8aPiInO66DZm85TqRroGB
zYs2TbmG18HCEfBxxe9eUFJy8K6g3Kp2f8fhd72CCBlWYWSUI3Or4elQw6IPqLO18uiUfoB/x/OX
8JZeL3c6CwYr8sDHFAmFQAYw5LiMpETCSvy5S6X37W2Z3mhyPoXaxrlfnTYTuTKluKOxjlPZyNUM
4JxmlM2gxcHELkNLZHnOYPTVAmh9FjxLJsj1JeYrF/wviLjIGdpRQE1xm8FNb1V9HaH1UkOL3mjr
+kBAfVHjrqJJeDZhaOvY/BYxPtcVNWZkzMFkZxReTy1lus3oIjKgvhf/KlcAq1x1agifsNAsTrkF
iu+MAJtYsUKpdRIcxLYvQPk/HzI8qR7UJsh3R1EYmh6/edsx7Erq+SPLfXrHzjtvO2wFRGr1X+y1
2JjcNXyuiVsKCF2G+5FdTLi/jX+7QTvkfoE+aMpnW0ycd+KZ8p3IbmYxW8IQsQ9/RfElC9X1o5xL
hPnLhNFP3oJaNgobIf9BLVLYmu3TW4+Lf0IKORvBTqTvmWsk3UWlEeIcNDDnoeGHCjk5n3hzzEpm
NmZIZHlLmFg0cQ2V1FEYeTLpi8FsovMffXAkyop8+0nr65Q=
`pragma protect end_protected
