`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
GtonvLyRIHa0BG5ascvXN09MZ3qOiFCm0qhQWasCekdFVRCizFoeirO1cOSD3S/L7XBtqzCllo4q
Q7pZwE0bdQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NcAWItlcyJiW5iNdkc1sQhABTpjXqZkOrg1X+Tcfgn7grREOKMnmze0hKfPSK2fx03p+1DXa9nI9
aDMO4y3pcvrSQRCRWXgMFS2qba1ARCCZEOEfr1i6f6+Nx8FGN5X5I1YnoGroW/YZxqunrLG+EqYi
XcxUyjBIkX9CxLSivhQ=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LPH3S1XGG8M+74c5vorJTX4Jd0Q7p5hXR2nHLPyVATbLKyNyCj3u2979H/5+r0KMFY+Eci03CiNr
huLATC3oqO+Ri3s+z9ShUHH0kb+eyBSFWWv4Vz/y3dKeMo7xd/qiF6cFD/jwZmVC699OpPLFZ+//
+v9QSba8dbzt+SXEN/jt0+eliBPMdqYocom4RnNiRzWVLRpczdP8jPK0iZ0dswvulkciexDQ2OOo
AH7xVOxZOGncQh6Vnj6rFermvVKMjP+f3wo5tFO3kt6qIlYJvlMl4+beZEF1FvA7E6pKL2F1zinI
FTyZEqwMwZWW/ux/d9gBr39V6BUQmOQXaUku1w==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XhsVvFI9R4kEmwKEMm1/ve3kzL6X2enhhJxnoXVsTfGBwYA297bpytmIip5AhwFQisRjBoqJ0K8l
8Pn3j20/SKo4hFrQQGF0dNNW6natF+zLk6mmfJ9vN5kjz0dnY6GDFbN+3VxaI7EfmTameGip8Srg
gxxI126PbwVBsgU+CTpGeuVit895aMS8BmBuDurrl1wtMGtV+dEhJIRJc0Aq1Wrns6Y56i0yfgPm
51nrGVg0WniIJHCwCd1amAGBP8K+XEMqgFg7Ax6FDLMI9fkEMpr36t/NLdEvEWInQ+uThyiFxWQr
JKb25unvEuv/D0FeWrozh8XdjpoKLAw1GPNMVg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
W3obImnatzWtWQxjvGXfWFuKaXr5FfPdOSZAbNOW8Mwmo4wQnwYiA7HkLDXfdrmslndHMaUxH/ah
zQFKiuR+SbrPT7aIULBLqqh72i8AksoYWph5t+HS6djOrRH3vsKtdR3ywmgroEjQ2QUcAo6U9K34
zqxoj8P9N8GP6+jAQYo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
p5NJqyb9TdyH8yE0AGM2W7x67vL0sjxs/jTTPTMrKPRWFxxZNuqsL6RAPf/W7gzVERxAO3iFqJD+
UoyFnOxci4budxkwr1k61TSgdoxD0V3HQjFvRukqTPnveyj/ep+eTC4LGfMpV/TPdXASgmKbIegz
1MyLz2/mIQLVdf6YMINHpls+EKIpYMQZpwK/hPkYr3E3OOOvzvQxNC9VDhaDMvYytD0fGysZMNYl
wnQ2rJfehLe6ywYzM95pSaORaRL+1Yx2J5fIpMdmGCqTlIRPg/vBGdEvfU7LTH681IczR8haG53W
YAR00ATaZUq26o3QwofFA/jZlZZYcN6rMAOtfQ==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OsRx87MiUvQMyOGPSETijoG08vE4+CeK9YRUiBEhaa6o5uSa2mSyUldHexlwxMR1rBWiQ6uyqUCt
nOrLjKhAiPGydi/JTIixYfKsNMv/tZTwiL+UoHRiZBVFKKOx3LAC8mgFXdUdYGwZnPhPVBIrRJxE
Rc1n40BeUgXQa/BvVgZFq1WN5zlUWx0e+VzL4EHCQl8ppq0b9oCO2dY5tSR8oDlWW/ZOlS5/u72T
OBDaxVQ+J7PWFUnUbY29E2dI2dNIjwjCjYqO+AssBOBH6HZcymhsJOjXSsS6xO1jpNeJMejZ9zqd
GqVBeDYMHSNvyuKhK1iLew/SAb/tdD8vIj8Gsg==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AYMh8vGmPAmkV/4T9vXCAbcwNUQ/U5Uw5Swerl5fs3AFaCZc0Qd8qyJ+58+zr5M2R7LYmJxqm46e
wTkAaUYx5X+VmZ+SG/c+BTOKZ03KypVWl/ISK1LXC/o7S+auCccud+8zMCxRUsKHuKYyIw/9r4Xo
hq9KP5hjv/dyE2FloIaus9WXSRmy3BsOrnOz34Y21Q3ThEHJzIUzPC9BzWKJqAiXhmZqFyQNpIPt
k/qfbsSvBqSTLaJSexAjyCb6KJ+cjdu04kb0KxNQHwNLCdnF8ejcSevf63EwGkmE+UzodGVDp+ZB
5rDYdmQGjq0EQCsB9QHiQJ9xNvYS9co+5Ki68Q==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ft/0b3HbGm8+/u8rq/UN1q9QtlQ7ydmhNvkUH1HFaaEw8IoZqW/LGV+djzXBf+a0L7Lslm4B8/ds
ZIPflSuox2viiVlo6Gu/oLKkTEg1tP9VJQ0SBlLuKdd+1Wtm5pN17pffr2TMr03eYDI2Wj8CqIF+
sz9vF9ralD5iy24MBrbk7D1MMaUjK1iYLEbGPul5XaMw+wCbhmYkQz1aq+m95hJ31EOKL5VFcBvw
0G1ICvealfGN8TBm1MOsgcXCDnEIfZlhrRoDLXx1+eTwJ9G46IioWqKUIgceTRCiJ0HPDdCrElbb
sSVKrR1ThH2yUQnQwI9fGdD6wpMKCSYrtlh7xw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 44400)
`pragma protect data_block
ewowGykr0Xg9OiH+t3U9Uv9yEPftrL5c8Jw1+OUcF1HoBW+M3kb3SwHnOMrwUUx50zqjrWRFafSA
ZwpCFwispzRv9DNRaiYWYKQuTKnjVWQ5pq9KmPKEKNnpQpSFcA/vrTNn2mP62c82D4Zv7noJ0nld
OYZUv7oc3WfsBc0DIBnYf1xMwBvk9PHHSVdFiszqRsSid4fCOIs0iE3JNpW0tQw6tJH+TY6ap/Pl
CSwcnRnyq0fjXjYpLUDgNCGnUR0cbv/yvDoVLhdmv+xcae5+0SkvFJN/eij7aWB982fomlQcMBU4
A3kOz5YRBFxgBYP99rWnBdVE4khwye6kxqPUQ8DPn3l44mvxz8VSjuMMuJXy4AugE1AVL/rZDXj/
kPq8MmQ/SzU5D6/lx2SdVxcXuC6qzY2kfueabDgcjOUbIjvDnlSYQ76/U7JL1YQN0mzNCm1HvnUd
bAbyBORKw1dvjNxbQSQHDydKQKwJpu37auif07dakPGeR7/AdW4fAeNMDLXE2NR6dRVK1hUFER8l
6MM0ApmM+KRzOhXC90ypeqzPZMCwfricO8fMBsN1EnxpEbkXi36B38HZf2mAyyKhsf/bgkmNDL+y
9KZN7ZoLq7fbSHuX0zyUB1S5N5plXdAdcDwaA9gldDVoL4pPEw+9XzmeuZzT4Nu+157CVm/j1Fev
GO7pHdA3nfdvD1rkPt0o4SSEXnrIJvpQT3iUECvDRc/Io0/7DG5O4Te4TPF0M1yRScQfUO8AZJRs
eixIzLT4JoEsNDcfd6zg5JgOb++x6WxlIdPgnwAZgZwP8RG4r/IW/9KFgVee4cGH1YiImXs8R6Nf
rx9VmSxe9d5L4NG3JXjnOkILKwdHR1ZPrru9BrUnS1QC3N27nbOyrBDDTy63hTkZUXvYAjzPqx4p
TfXQNoKC1ACr80H2/C7/3MOHnSng9a6dMJEFUy7VtgHnCOLawJ2XlnOSqL82E733Av4cvZA/YilH
p94cTex74nKgtLy3Pd1muX1ttODk8CO72k/7t+TMcXO3WFEe2nFMWPIeBsLLqIiJ6nCY3CNega4/
RW7hE+EZ3wQADeutPUUYDGjsRJp9S+GPwnsaurrWtqAY02O2GmmU+9lMbAW5TXaOvrfhKDnF10bx
dG8NDccTq3VsLYwnby+77W+9fsfkVqKdzQa3S8T+ciDi0e8okSnFNX+sMQgOBXI8dYP47HTawsqe
qx43atay7OrlN0hn+VSL+qI23/E40ye8Rlgc2i+zvJhQmkjMF/4mRsngQf67ALvDrsq5oZm4uYtg
nTwX2vj/+6ZxoNBqgYecZUzwos2hOJhxCNsP9SPxLanU4cIjkQFOMPhrtP/GoObS7zTCX58N9sGc
+AJZ+l+K0eDPY7/s/XPN34chdDO6RlT2MUq5v0mxsZjps1AmtvudtEgQhzzo1WKGt0trFH5NSy90
9F4DGI64PISSqF37MjxTIdMKpGJQPUojw8RER79jWjnXGwBi71F/x6XeL2ydhMXGAAlIVpbydISV
VZCzZqVE7vzwiA8gVwWK5hOcsoOlVIhDpFNZiCIa8h3Ssl/sT227BuKiih8/ZQ577Mp3B+pbCbfC
ujK11WghO6YOHIMbXcJBGwdcClYtCdBbiW3fpVCT6EqgC3hLP7VQRM0F48Xqpc9PHJdoctUqhT5Y
RBtEC3OTpjB5AOnmUyr+H/0+jeb3+R/dhWLg6A3AP6X8hAtm6HbZCHp+NFAD/ZuFdCSps1BZ1Amc
iTWbLkWk9nm6rn0l7qamQPiQWTJuiSpSzAuSJeDv/t9zMa0I3CHGeDcupL/sMKBPsb7yd0J3/wD/
vUrMPX0NYcMfVV8hRvnsQkuIzz58KTYvn6p2qTrEECAdYkA2V2xVPid+3aJvaS5wbsiafeOr9GBC
PGn5bgRfLzJPJeeRxckY+AZ45sMx0ZQ8Sp3oFc6sNDyLsGnE7618Sv2XOwNI6Ar8Fjcg22kYwm2Q
AH8L3SrWdXNWbA7E0GwfuTF7ewQYytOfZcBokX+cSoHFz2hrTss09cRbXF1QnU36+nnubKh6dvLr
VJtTLbTsRnTcw2IiqtMdodHZxODj1i9kCAbbsZ2iq1sZ1n/ykzzf/UW0wcCX4Dvj3TyJ6t4FJ9I9
NKq0qGUTjG6/WUiLHWhqq8sXTWmGrPr+cla3fWdtEUOBxu00BcZalhJqKN5C6+nbqO0ksw8NAYD8
ZBcacSaQ3/K4jOnFWF969OZ1UXBi+MeW8n6WAV1F4VZqGk7e+rvA++JcNj2WUh2mE7agaFPKrP+x
s0uuEqqwBX0K/QsNPdu8N8gZBAISPQIrx4sp0Mad9Az0Fx20xZtiQkwgmQFiO2sZbd6wL2lavw5L
KE26T5zDPkmsvcZkzGM9P4Wl7Zb8CP6dgB69CgENK7Yg2vYDyzCD8AiFCwtLtoG/iVBNPBP6DyQ0
0PUSTs3HO8gz5asSwZ3MVf1Xi/Muz6bQe5SgM6ZxFP/0+vvtKRHneEl/7vvoAcXpSQPRcCtUPjb+
F3fORCwWnnFR2W4And9bYoXMYG8OFN1G/46Y8Pt2+r83W9lLCeqBT3GMTU8gtuFxB1MFq05SOWLs
bm3yAAcstTNBqNe5gk+cXRGzNgkU3RaU4g3ZY7JGuL0UCY2yP/HUiJpiWs6A3h2SFhMbTkcbWVq1
vHSGSwuTgkw8ReVv0a5AhQftfO3VQfdKn4jy/xsmxrTM2zHCwvo7f2L88w+yrv1vJHQJSL/RFudC
1yFm9xlAYjAtY4d5xc5GK5BPDbgGT+B6d7ZAHtCW/Tb67uGnAFWksgXD923dG0KG9ssRIX2goN//
Layn0wCpwAlSjtDkfOzZg+UrulGYvqTk9jKad17tUBlntrzaEXDzz2iLIVMY+HUjF1EGz9Sof3x6
YfYuM3Ehd/T2ioFvfTZV+0Do44o/l2fs21vYjhNmKeqhwUAd9Y0XyiuuFrFBh833gs9EDkhoiT8S
bwm+oPPD3lqZGp6wC8myCcVpPEK1dPiKYh1lJN5y9kq3hsWTKzGIU1wNA2aRMNVpCuL2/x6aN2dz
nNo6t6Zj0KBq7AlnMRnYh46JA6IhiJPP+0FCsgLPdKg08mSlkPRzvpPrGN8Oo/TMxPZyQerBidMO
8WuQ19utEY3ttV6xX3eEsoibf1ksISWRcL4dYgi3Uh9eV58qdfegfEwB8Pg09fVGXvEMaeVG/NL4
PoKA+A4b0kZ1D7b0Z6mucuKJ4sclQL3nsunCFKrWp9v47NFjOkwVlAM0lHIviwg61+xwGc79y2ix
zUEwwgDIUUBqi/fP0yApPGXXX1NWa4UVxwENSrtpm62YJmSJHPzFkFhRSkrDaXlUbX9HFRbeeqzO
l8zHCB9PA99mL/eQF40qftPELR7dV7Py9auRpDHVbusX075GyLY9kWeTp/thPlYDiJ95bL5bFD1E
BkI3ELIZDdAkRBfJCZ9dQW77/62c/L124iJSnnk2/jHpm8gnae1IGUn5FrO6rXdLXaVDP5U1fGWM
eaCWd1DiThyfkp0tEp+m4zw5iP72xqvLJjmu8jERPpbVkW07I1u/xX24//WwpFLvs4/OPki/O6z+
aSypG91Siao3HQ7u/kQ+clAc07RLChxjxAoZz+eXx24t/Hnad7NAuAsyFmoFaIasChiB0J4Z2EF1
aS1NhOAbyNUI7bQjeEFHhqxd4AB+Qfr7usxE5GZ1z6aMx+0NN+ONoetDtlyGdeldFSVf/2wYeQI5
te50SiV6PYsL2REOC8Ha0G+L1NYf3jInCRmEr5gi1T66Jav+O1selg2Ge6Y7rmNtS86LiW20J/nI
no3XifMsalVJHyC87SuHPtIDn+kCaPOKxPDZZ2Xg+zyQq8sOYkqF2+Tomfp5FM/KKIV0YGJfqZOc
UI6yr8u9RpJS98kMT4KEgSdu7l8KVR1zMcOW4k/8BtXU/5yVoRNcHI6vbNRLoaceoy/aao+xfI4u
8/CnzOdqwWHKg00PsvPdPWN2HRqua2I0ok6OM9ArdVh7zsn/zCGeDT9TLtdXq+RQmF2s/OOWf4OK
GO998Y1ReUqU1CisxBRYc+nPGvXa2r4EDn68n6ZITPkdAqEH8h4Wo0H2qMBxXlNwuPVLDL6GYtDY
Opeqtdn3J8WORTjilR/20Xka+G+baqSJaEBcu8p0r5FzGE5SYkT3re9c4ytihTu8C943/0rNaGht
1iAFzvbZsCbdBHLpZQdwr4rjxIcWCv1Fz2wzrQuPfR6dCJk8Y342+F3LSVcq5SGWTd0vYwgx1R0r
OvxnFGZP809Cu6qWPCZ9u7XxjeH/zeUyS2LZmFIpF6snqfG3PIJ3aAGl3uLBypYf0YciaKpp/9R7
1jdxPUGICmJ0yR2/uHlOoGIpRptD57D+Q+He4EpSZCpaY1F9SZ/ifO0uwSIXToWF6wqY87lZ5o44
Wcck2tyJ0U1pe33fuPmNeQqQN77OqKkzTwj3r/SVYcB7aYRcnjBWFNAIFQNSwTz/RmkaCBISBPys
p/cO9kDXf6c7/CNbI0Xdm1OOejgnJoQ18idgzcWTLTGo8s7XUxgmTCm2STRfzXzLCk5zpSMoVnBZ
rNLUnew1xtNfaYQZfnOnav4yjdAzW5BcL8xpQzj8+Kx868c7m3L32x3ntK9aBqf5pATvzb5knpXg
FuUkB9yvRm+wmp9PGWSUKX2Cvw6B44F/y1QXVVyzOcQkF3fCAuzbVxNMvWm4hqswoBGvpjeM5RiI
cYm2IUEb9Lia8OWGbZsmZT4kZk53/ofQSUb2Fk0SDLWA8952CmJ7fWkAHQYDzV/XiUOVZyu+Rlfb
HmPYXFDprGS1jL3Qt7u8vDRY+9mKVY76h43YpwdzdTzLUJLZFqDrzG1U/zL3MdemE397nyc/OC0u
hrY38gutCnrHoGW7t68B+zptax3thKVUBq3fUadvjyKWda3FGv9eUGJutO9yVyeV7bc6WRoFb9pg
vdaQ8gwrsS18E79dq/F43QDzJXBJXzOMTBrr1BXJgKgcjO3KnyfPb294FG7XTdlcAzYMsRWK28oP
XTHKdbPJRkQkRLFJrYdnPIDvGxTytYVMWbAe3E2JA2ZzXdQK1DHnI5+1koU0XZWLJO1HhDvyBvUK
kawrZkwc77aByv3s5QTkEgtW+rbFY3lznpM7cI9QmZVsuxkviSAZZrLV9kXrXVj/jZksrOOBtiCd
HREro7zYV1CnZXpgjPVz+4cBc5nvzfIkf5Iw+lo5B3EYBM3ZNdZ/qAHX0kszrSng3331BpKitkwg
sumyZTga6LJzlqxPysciMMfSaG4sdyJ9Q0LQJMf+04ShqgfhDQsnZLvQz5VDCVp/8ps7sOhp9mlA
3pQ3wzv//eXqGSNZdF6++RVRMVOACs2AiXmj6dXQMEKGHDmO6Pw0/PGDAjWuGQabFbdNFzkDXz8L
AwxMvYnAIK37lp9mQxh1fsJbzpCWMEPRToaS3uKWJD4+E8oB/u0FZ9ac9EZfvnxapfUgyPaF3+uz
czT25HMTT/H7JSmxaWLmsZr1NdZeMJ/aR2ZSNUZJVfnAQZ9q+00Dt1MO6NKemkMEtrOgxZ8HDUhN
pxu+6zBqjgcqQg1j8ORedtvnoU66PIuBIG8iz5jOZFvHX/PUfj+eZVZnK2PSzHnuonoPGK9DHbj1
XyPL4r42J0tZGwsY7g8DFYOXz4veBUBHNxRcTvdXRjkrVGy3RiWG77Lp+r/+HTOqu4CBCEm8Pjqd
DIQKZbeK6wciW2c1xBDRMNNBdDvNPm7syj1IcfqztXs3F+r9mj2Qw59SeDGcv1IjW4DPBrFduwAJ
eGUlbfN22l5vpQGfv/RDx0Vx28HeevIUbad3GyaUO6zmt9615BstRQYjXyqeKARWLcmP8I2RFBab
RPLF8Iyx7DRVoHkZ0J15+u1wimZIMeJ14OTUqJ4m92Q+ycRKMFJN0gb0mSTzA7uoM9B9ndlq6qA/
Ko8dT+nmLwYb5dnWsFHUtJWIxg+AdVUvLoafRwBXM+mGT8MpWzPNQBNMC+xc9kZOFn8/VOGUIC7M
xnL1OklV8a4/hAExNsrb6bBeSmhlUiAN1pHO8jj+VqcQUCVXsQ388dFIK/1YxMMBpPZg8IcajlmY
FT8KpxuSomnTDwG+fGUrpUavUabVAYAHjibK9fQHXfsW3oUv2cr0CGnpB0AMMH5V6uT1Xqa+OL8F
oE2ST6/1WhGUSE76qWp1/g2FYWXaEmKGNVqll63i+YBib4pXh6RpYpQIJOMBdD6Ea8UTL/qa+wGs
Mnuau1VyhzL3paVEC2lbok8K2uDuGySeKeGT/4ANGFKvjnmllGUjJrxLByCodvhbD7EfsbGoGbZH
35GYC/zBfY7oztM11IW8JfFsClcjAwp9uiVuCHYT2MxXABQs+6MOFPfiy0XEvAasPfBbirt6r0l0
4xdt/q+i7jqKhSq/FoHhRdPJ24nMvQ0zaQHzB9LGbBK4efkSdfPSDveQwbOBWV18R70GyMjC0ZaJ
A4QZd0Nrw5TVVXVkWDfanbyJkAhhbMHwtQXebY0cEV6sot6MGYXRkcjypOevTEpEAa/1H0r4zk40
rKrlRB/9pvXRVqvyLmeOAzHlaaFPh92fKtQ/IAaPXP3N0OAhdINPL6KPsh84mK94rLYPrdy+XS7n
KjhQHoE+DJxxPAWgLiiCSqwRZESLG6BBjG1MTn3SEXpO0bpP5WOn2rfgrWFeBzYDrXwZ94f8up6V
mYtX5a6hpWKusLeWlTsLHk3AmT38GOZw2ugVa80b5thsJ98kqHjM0+yodh0jb8Uw9HN3Nld8gUNK
MrI1uw0Dkp2trUkidbMfMpJUrXDOTtRf6wmVVGmCZ96xGFdXLj8zen9sj6EllPRjx9NFGM33l/Za
78atYcPSpNAspwLOUmeC4f4+ts5qwT3QWxp1A2ssNVCijY+ZcAfdHm1X5p4kp+2iOvkyQB+gXOA2
dKGIk0Oo9aght0hpxvfDxnbtPByunAyjJ1rkUrtnu265nAFXwIqllkSf/mKmN+t9TJlMQDpkhWMv
fu1K0vc6Ywsf7cCuEZyfa39s4/rgxkFJqSBLVp1kRAmoXY/2czEdf+thb4t1y2WEE9VVYtxYPRvJ
nRuDTKntkqk0TkaA6DBw49ZE88FENkRhr42T6r8e0CrgIhD3CgOtTCNfbaDPsi9XSketCizj+kJp
9dUAid8N1W4AgQki6SHv4hPZr9tzh0N1EelSkdexWj/HoSkjcBgJdWNwp5DuheKTMUxfcjJyLVG3
fJ9z0ZnmOtaSNgBRv2GTd9o0BhZ11BzNZhAQ0Gg01qkNiuV5K3bUTZWseytwT2LHnjqWO234e7+d
lb+5PiBJf6dREY6Wan4RuM76JJYvzOTZZlOqG7zlEP5eAzFpqputOMmP64yBEPfS2ZIZUmdTWnZu
ZVqWF+AjAKmmT9dpRup1NSoCIAHVSzXw7lbRVuaWiw1e2gM1d/yAOJMyihVHDDLGBu/bFo22Gkzn
9jtE93T1OnUC8SUH9MMV1VBzED1DYWK8ozo+Rgw+WX+cWYwTaUC7LoJi9zVVLa35icrFhhvYa3PU
yV9AzjANRkyrreDVR3PmMieeBZvoUvuxRMWuWacp56ws6ZIdueiFxM193bQ4PymO8IdMwzegWd7v
AjtKquNMTWPzaa5uzl+Oxnr9YseHxWjJ1iX3YK6GpyQ+Z5SfglRXAGPxi4dHNwDJsGzgYF8JSHOZ
p3Z71aUTYBoGJA4pOESCdslxDtEhq2KHVWYgBZYOYal7Hznk5YG7Vt5S7mNIma5siLRmqOtECWXQ
MI65CMRgq344LTqMHtFohV30qer1rcqoFuc7L3dw89P2iAmsnHDrL63ulPucJMC5fzOvtAl9+dDv
3Jgkd61flE7j8yUTzXNDxVjA5HvI6mSOIxQvtlsEF8I0X62uKEf5N0Z6GbAGqaUqw5ut6AMxoB6+
adchUapoWEow5zTWIm49dsTEqxjhxQ/6itMIir9mnHD7hXg7Dix6hn1JmsOD3XJYCDh6/0d1nPvS
A6TWaF7MZpPlatf5/rLV9PCgyZlMp/eQSfBjZXj8oWmfmWfBJiZYJDKNORBFWGVseDCzu0ailcAV
c+D+cce+E/aYWtk57OKmHMB/DaHNZj8VRR7JwJ8zC+D31sY434yCVNO14f2jnFGwuQIqZlobNitP
fVjoDpDGafJsY9GRHmslZP6ToClAYFZ8c5hw4GRC23mkr02fV0vaJ1Lh3KTypZCq6CVxJlkFvdH7
iCjRBAMuLtYtrCLVjzxzkENIArR9LSChjnvqojenG2zOte4Q4tFnKHbtuSn6SHN0/Cyc8S1chVV8
TILuMAN3d3oTKP9b1q7GZVozakUcNy/lFeW/fJMDjmENdao/re1Dm3xGXpK92VW1X3xG1VaA3M9l
2v7Kz7+XoxIQn7BwotDGjSK3LjA8NXBfyEDc/WeYfSnoGKekp8njgPVV3V1bSNi+GzJQA8kA3u4c
ZAWtYOsx4uZzJSRd8X720xwGiMnlU+ExQTVznUpetihDugUzNXrHTaGf0jy8b/bjLcJ3Hw1froax
C9sPtiIaH0JXMCWv0q6KkndWAjPOnt0CZAQ1PMctbNGDj2vvue+QmVyN/N44/8PwWBKmz71O6RMT
PBeBrHhG/Bywez16ASI6YkA67ePnpczInK5jSd9jK7EUiHF1KiobLG9IYnYuQxklRDrsxnZMeEwL
2LoGageMdzJxVeSXhJIdn+jjlVebWGNguaL/G2lv169p8C1Vx+JkxhhpeJnI/9ZsnZw05Yj79PcD
LxTgMXabHB1FmWGWxhcd3YGS1Df5S1IJjtsap6qlMl2nu7Yo6NDUU5AShGNzPaZWbRZZHAhhwCOz
7eqwSfZosMjQJjKF/aXCxcznDN7aio05Ii8//7G6OHeJ/ICk4kHCsEjBPsvW2exSnnhAx6S1qMNW
b1yuln9FhNKSyza73HYqjchEAY+E/YY3vHUHpoJpnbdBl7cc8yx48p/LYFoLh/Y7Il5QIT2Lkct/
c2BZGiW5PgzTkUr4iRP22uXluWmeLw2qiqhy0T/pOK/504bHXwXfSUGtt2OmDW+PGf/x0h923eWt
HftB4fdEn6zy8600gMIOI3WL+LPZcr3Uj4IFfkdejRXvw/ydkpAAhbbEh7dEumxB2rvOH8BsXx9T
i7thoy6R3ZJ0zT/EM1H0tB4n3Fw/BPNY3DUBqwzAQhnnxnv7LzBb4H0fDJ8DLi3RkzjMnDBKCKxL
MJhLrT8cmkJgLycWXmY8+MGirJZigK1cwhKsN2l1A4q6M8QLqNab76XRVs2AC7CqmmfmeJsd6bHu
oDWDl3idpzRf28HESl2SSvDnyEmlhp1kqLjuOzAusbQcNiHXJ5/GDfNiqCD+nVP1HgGaS2tzVmc8
yD+kEr7l2qNDK0gHpyoQ0Y1mFR1Hb48paML62xrcxI7q4kXa23J5kGdBFgbMbv3WSz0y8lpiPf3e
z/1wFtmLUJzXDxUp2OmtXN340erjYmC7JPme3FB5r5LGqsaYuLZqXi+o73Dtv2leXMgT8c/rrQbA
x7EPcKj9oczGVg8Uggj+sAlqCRzNHrSFTny4PoSf0pAMgzd3qFcqZxS/YXWWqtJqODcPFB6Fbp1s
6vQP7bjahFmkLTT+5+1tSounNQxQJ3LIMc0/ujlv3ISMYuW4GIdOzZOztPaLt4S1/dhQq3x6kDfL
j4lccmT/ftNwBiSlwbxLZDcYEfSU1jVMRHxH9IaGn9MZYLcYZhqRtSmwBn4V9IeV66bBdanlkefk
KozcOUgnPjeeeJqivG1XyJ8WxBt3M2A6pUgXhi908vIZcDGCSu/as4ULEDZqyjypBdi3/RJmxjAj
GNcTncu6zpfFFNYFe8cWp7hzp1WFziGh6Fi9hqcaYamrGLGQ9Rhh9xNiIi2ED9lF6nHnuzbPMia0
9mJR+E0+ChA3RrMtHYj49fLOoWVyQ1+/AUkIkdNqv4E5G1DdH5tsXdpPxxbXa7EBTJYvUCTADAmb
33vtFanWGoZq5mSY9Ezob3SwXExR+BuFzVYDPi0shAtcKrMJclvpTwejMSVEMcOabztvyVA/Fkb5
sxuVrEmSrz+cIngmFIjVLMqqfYAgqfXqO6/40aISE2OwbdqeJZ4zxXuc7GbX1eU8OfGcLUFAAQLq
ijRAbID1eY0/Z7LIqlT/vtzmqBMBRJjQCAAUGvE9SAubF714gIJgKT7oG6vB9vu1UxbaU0TawxdD
pIYSLcL8WWCfQ69+RhRpvPKPC/uKy//lpvzzGBeewqPTfpPk552vfU7L1dYIjl/UQimkQcffLL5K
tqV9OY0sR5w0+orwbK2YJg6n20wVYhRsVzT//qRTSCquXLCysXQ0eFUcvljuPCwabKfbmQK7JQkM
StVmbfnb/Jgh+Vf/lRVic6F3uqpIGhAHDzXxh6g9jxUT+ap0DV4R7jifFb/tIsBI7AfBS0vwTOTE
7yPPQzoJQXWKG+tkig3v8ovTo6Uakq2hug/3rZzhFizESWChQ9kvA4T00GfDRJsB3GNUMH+23oQx
NG0OAbnA+hdVKG+MzokI5EhI33wwNH7XKb+NvruGRXhXar4x0mQAfCG/LOEHPqT+m+pexcxSlJwp
CXOC1wMQ/m2w6NRS2J3lRXxLdttwfkYoxvBfXLtapFZME9qXe/o87aTMtj8sz6QKrJXBFTkUwCQd
lm8ZGpJhSlBz7qpGAHw8oAxzES7pTR64VY5xYiDyB32Xh1KpPidIh2ldVlAdISmFz5dSHOgBFYZm
e9/tXSuOfja+vKupErjsd6+8HtHyUM+RkZqHHla/4L9N+c+BXJVm5ZgrWlZx+xrD2sjOxQ9GQzTY
YVS283n48yAuIaHeZDT5ml0WYwMKraANeJ0RREyjO4aSF20GIV3eeD2oEQS8dEuPG8t9zr278Y63
CGyvshGw0r4U90oPB04k8oDbvMemw9z1vSOcx2IAwgen0l8GNcL5SHTII+MlQ/CrUkbF2TJEI2Gv
OkgTjENkK09SD2t+sBmwjmVnqxLvW6qVw3/ktC6QY3pROgtbMOcHtlrHv5DjgPY3n1FLjCobdPgt
fRT+jeQrClamCN4hvFRvBXhrbIYez2ffriCxoY1LcjJFXKn4H6D6MIgUAbnsBrso+vOI8CE+tCvA
VXf5VI143XIlMoEBiiSPK32xPTz0hKPdtjXcKk2x7izr0FIUN1op0ow8NnC5VBj6454OuP2h7yos
OaR6T+BAibbSi5Kd41QF+piy9iD2m91KQZHVHnW+AJ3oHm34KXjjwjTUAQzQEqe5bVGkRe/wQ0Y/
1MxziRKXu0O04ExNa2ReXaznA74QGsl95srjNFc8FxBONmcZwPuMLK2H5x53CiFzrpWCdOVueoIO
RxK51GuWrUT4YzxfqUm8ZZMCTn3q0ygWpAJ5rrucDWRbeWm7cEFzt+6PMNX3jiV0eCKy9nEii1tG
9yy5jSoGR0lUAHzBZyVJyoMM6dcAenv/8VhOJLPP4Yr94/2TKRVFeQJiJAUicJFackh3jrZ+FaHG
1Q3kILruzP/QrizcYJIQImQi9Dq9yQjvVAAIfOX5dvYOhnVh9UWDvnOZnCXaOyHRF4nomSZYOFob
UlAVLOKZ77I9cMRPKzvamu6B4QviBilNKiVv5fZ0WWHyNG0rANT4IhqcTucM3cQB0eXQDCK11Hjf
6Jy1XQEoQRpGMeexGL2QsXmnGpK36NVit+lj2EHUktpCuJzw3pao77csXLMcgjBcCvHu3+WCJvA/
JyNLa6ZD9dA+plxBJo4ogfCzUOo42QMcXMo3cXP/wcybUvMis91FVEmvMcQD1hvP8ml6iKzQtL8j
Jv9c+PX96MlM/ln8d0x87kwVyydFweQSZYYK40zSLW3HmLDa3Mke7SXNaO/zGe+UysRRUPEYEkR1
tunSchnIxgMNNVLRLKV9Aw7YkQOOWZchY0AESJ7ao1iEv5hVng2k6U/dkb4wV2oi38u1y1ve6lYn
6oh6+Rg8g6I9V84wvPhqM6e6C82FxDGjiZ9iGFFRZmmvQ6TgP0NGx+JScO1p6NI+Kx0Y3no6g9RK
u7eT/AMlMTsEl0T0/CrEfqu+tZOZF+cq+EowVNkc9MQTNzwh4IkHzG8X4fhdcPKot/cBi97gbGcd
nFaJAaNjAtVlW9Glb35alSrihIfraHp/ZEQaP+3gMHiFFwiU1aGfA+E6ZSP5ki3nwslrRzmeZMlk
X6OdYHjzn1/QHaBWpaT2LBM+qpY//QQZNkToTQTtBNTY4aNqpYsfBF9ACIdz5Ki/vsF06KBrzPIH
3mxD3vWWO9b8fjSk/NZc/TLKajATYoWfqFRG9vWT4s55M1uRnFnYW+gYmMN0S63YWLY6wiADWlFC
NnoY41cL5Y0iI9HzI3KMhnxg+JGT8TP72WqxSZDQTHLPcP5G9SAcIk+Z+CMUS6k3W4SfigrHLg42
LWFwApEtyY1anUaAQMGH1kFJZo46JSCifes+xG3zWrU+FeM9DtU093CF75aWCvJbhqH+nm8nj+vH
pwhjPEVhYmO5f7JtWszXQmsIJ+af3NYtIwJth8AkFlHMi3OpU+1EhVTJtZBhkWnxl7o04/QwkuYi
5csdPNr3/k2cUTPfK5LI8oeAx1BuTyDBV+jNr6XNKUGxRANBupOOvlE0sIgaL70cEql/w0xTQVaK
02pLOy7VZVrGj4Yl5e7EBwtbTN2hNs5Zpv3iADlDSqhDQtH7iYqVw6OJWMyIA/DVAS2yzttTjn5M
5QJl9Gg37cY0RkIHAi66DPkTtEZwZTMckZyxsJWgHGUBZqQKLJCZOqLRREl/leWPXPVlrLgl7kmR
bTcbSzjdFMzjkS6vODdcxYawUvJ7s1dL8ehAd4TAKMwfVjk+pBanT9FiopImvB0Cx7phCULJYCUN
cQvAaR3vm5tGxPfDukEDeZflQyBbc2c/frG2Unr2HcyUm7HQVL7VWccIQQgwLiW7HUjk+vCj5eim
9CySpH3x40iMnNgVtwxt2tu9OcjjB5PRF2rETVSDG2haGj11Qzf3VRCjGKBlj/wOdQz3Ps0tNrYO
wqccGcfgnM7tdWdjhG561U7Y7nmS5nvf+YssSHFqJ33SUI8/dhFdEdd+3DV/a1JZ0zL24VYjizQJ
gel4KBOAI/qY0E7j/iNyGWqZBCkzTlO535KEo3HpK6YzdQcGjHoSEXjWXHrvMZ6cUD2MTDvCmhzm
ynTRHiQYTKRyCSPQOVCDpNhwDUvXBKUIsaQEst+wHWCgN17vWInMTpKD8nT4LnDEw7X/PqfR+5SA
cUIGQat40Yz3szgTqVv7py3A0srdQfj+4NJcl0jCr2IuwrSS20//LoEPFTpGkgbYjU4/nBKKQUzX
5eC4H1ZrQ5WEXzPSMt0gLIP7ZOvyCupln0ViO8PfCzi10Am0yEcGqeNsBjep9jd4tIsOAtTXaNFs
ufzJ7RTolBk/Yv4k8a0RGDu1n6kqGvhE4iVZ51ClWkEGPX+M6RT8N+symmCio0MX4/YWnAJnbslE
fK2yqqrz+jUmmm01UJ/rF40R7wC8ZB9/JmTyb4+YN5TvkPPhrubpLbjDnX2G+ogByXTmWGZyy5BR
0LunqUHQxixd6rydoypSG9pcZ4EIuN+bPnuhTtubcBxg+myvcCo3E1SUrIAjTnFlKLLT232Cazb4
VFlE/du9OUeF51Frk+OKDaTfJ52o7R5Hzgh/sG622uCNa9co+ynN20bzbjXys8xj/BSreHV2HgiU
8MXESh+7bXx+eFv5/oDmkfcXQcOeNGyz+sHEMxaood9ODWFon31xPfNTcjYIZiycRlcWz/XW1BY4
9C8ptf+nTO6RyfAtCf60rUhXPWFOD6snUHsllwQgWGAvuYuemIidK90/YwA1MMDeddLoRjtDtmVZ
Iel65MOEBki1p7BBxlWdlVKY59x6cAerO/YDsYQY1KaMVIefLXOFV0w0Mfx0hz8edq/5D8VKPDym
AOWlaAnjLq/e1NPoFz7yb8aUn6TU4ZvsPo9lHe/VLsekCknt2yNOL2Frs2Q2QQpAx3MsgEQwrq3V
vw6BsQUdIsC9iX5G0QO/GclYhSJHgm/vvkXLDS/tAHPCnvPD0mzCJDZ/we8xTilYM3WS4lVQ1Qx3
8iXXs9ulaPH0fuZwvHGvSS9VEOq2F4nUavy4y3BBEeIHPwCnba4FixtjAebcqnXeN8ztO/V/Ja8d
KdgxjTE2lsoqaC+E/OW3bA6oSPOymFG3P8lPiaPSa3d5hmvzFNFlvxD1ThT9kINhF2cjUBVwyAf1
8OmXi4kPH+9wd+uE+9t9L+PauWcLEOYt4hgWe6J2pPa8MxUmM6iLoiNC8548FQAKTVW9nXFeJgNM
Ujx5t00AwkLvZSfXkErB1J5VjzyCC20htXE4QX4CujjZ1Gnk8kVkYClv4eq4pRxFFfYkQLBL3Ju4
IaCZxHMqHR9wOuxfwfFEUesuwYT2ncquSJ7ZhLt8+f1AkjX/StQ/v9WazmS/DWhoXZe/fj+iOJy0
esgGGqYZF35qta8nO2qS/2elzHuHwT35yhxKJb9QlM2Y9K6HexqlF4c8e1iNnyJN4EEhEevgb4Vz
MueVdbIwTCWbZDAKUVNMjTuSKamfhvveYfYdCQgtTuRLMPTGOfyz2y+BAQ1Z8yQfEhUflfk+Ggdn
fESCsdTuAyPwNLZdq0jpU07SB6vA06xth+rUSd3e0Ty97ia0b7CSfVqpoFPzUzto9yPYstGo21c1
Eqr2+ZpJaQQdeNdP6odC1XZL6c+fBi1CrG6NY5xUEJv/NReATCp2seof6wSzf6Mwp68bRL4dGwDV
QSsiORY3lIyEv9ueVM9hN9tdSEJ45hnso6m9iB+LRNjeFljpJ2FHOstAHrsB4rQFCvECbV8NAO62
fDNmtWANvLRGSsxPIBbK5V0UG+aN7nse0u8nEhB746cFyC7fMwVRM6ALPV6Wez3vW8rkH76dvMos
rEexTUmvWtMFLBB7ay6+/pRv6vt98N+xQYJJHquhQqkMnRcxlcIQQcn7Ou111c1gF3fRgKZCBl0/
scM/PNvFbJ2ec1/mISCrAAXnttsibIBMf3E46eeoYWmZqqNveM60BdIks0HzDsCoXHGrGhY+xEkz
d1+0FVshymlyI1cQL2aZ55wKSBlOcPF2fntZTylkgp6LA9ven2qFd1waETkx6Jmx1Sdd6rgCuo1/
w/pgL62qgZpeIU+9Bw8v+i1cPIBo4RHuEvAC4/r+87pQHiY1SYHoqENULWs9ptz7DedIyA4fBPJC
oSEE8hZhIAoYAkvKslueZY7ENsOPlHGioBvE77Ij501hFhHrYxDpPyu1zHKcAqxMCsBh360jDYCd
zVc6JL7mPR/46gJEavFx40ONAdGsNwCjIUtpWoHMcBvMgYJa9emBEycorZTQaAFVDabHOEamwMYF
UFqnmPo63UaMUIEsvrEN9vVKSQFOlCSiOWRv/0tCf+K4ecuwYc1h67mNPFcLJv0nhChlNgLY3/t1
6ovXqU9wWPaSRpTS/tiljTG1Q0bN9ceUVvpRdeo5BlWhNfS0ZU86UPEAHmx+m0z788+MnRqIPnW6
/C5DPUHP38g29MgKV3F4qXjEAKGMpPCjZMaTI98cHfW5jW7aRK5rypYRK0WWnxvDuPMcqj59mYTb
vTCJF6dlmdDiWAwBq4cK4fHoueZ+ekd31vlXoiOfOmwgqClajlrVCaG774R1Bugcp5gxTAP5aODl
U7AWDOdjowxc1EVLP3P79sQC6svvhTX3ONx1P31cohPzy7DNKT41Dx9wI1qSXfzZU77a9fIrk6R5
3+eINb2q6lJDVb7CAFEG4CknnGTSs3Bx5ktluqT/2w9d0C4EIXmwO4zZkaaKraz970Ds/U717RaC
dDJCFzs/3o3ce/HML3gqOn4dV3iqJYPVRZqO2Pk7yudlqIK3lU8ZwJvTTCa4LPo+pLHpkSzMDb1S
tSIIGz2VAnqgHymWNZBudimcgH0YIErsL0zBGgNdYwVyzdy/sUEPXGSDt6U2glZQVPW6UXTGdYLY
noKIyXi0xgr9ugL/KzF2FiVIvAcpiLaCCQq7BtL8b57wKWw8wSQa2YRImLFBGQ+jYZa4ZZWsl9TE
NYwKHOBqE7xXaHjyeL/xSKl8E2xRh2hEe35l9PxdCUMHjhByw2Dmsa19M4+QXqjiU+8VEHez8rjn
XAyVNfaFKAfsFXRs9sRU55LEfqFfmYBA8jJvrQ4knUPocilzGb3S7+/LnlwpShZSFbgw+87ku23t
LQJqeeDUOW3CvyuG6iSeBmiDwRIVp94ERrW6kLt3NXRg4WfE67LzA9zKhmAeo7HoMhThkagI2lOj
d0kVuPkIly+eGr6BcAzRniiM7tvzG5Ch4jCEqxAoXOATTYsVoWGLQydHEcUpSqQw9RjKk0MjLsK1
vYbIA1cKtWqk84uLCO8afAyDk4VczcxZZrHc5npMcriY24t4FyrfBz5Cb0UeASWV5Dmd/y4010eq
xiCHS69CG0M4V74oYbXH6STEndalUKY4VMyWyM9FmaSEivYodgUDkgJ2/S3BkhithkpKeNkxuvcY
4g/1ZRHzkBzyehKJRjGsqDvS98bH4bojiHFEVLRKI5lp+W3ZwzB3wHw60UxiyQSYQo5+oyYknIm9
VJEOHlEkJekDY6UD5jtyiZX7DIrwm+S3RRl7TYe7zpSSIMyQkFJRH7j1nRXA92q7eWeHA1BgoieF
w52Byq/JVpdGvvaUbmxKPPIgHhnFG7JsUK6vhUk+wMM0MHo6IX3tg58M6z6yc3uj0U0AsDlHpuR2
0Iw0Ts+nTtmyQxpWSsBIXMsLnXhp+Gin4OIlK+W33AXB9472ShvNHIguncc38xNoiad2qEeolQvi
fYHQAYbmuZBWfde0wBGFJMUZSn7b70te10URxYQbSflCMYBnrADsDroWuYg1XQN3sIVD+dsd13JM
HZ44FT+MseodVoLdOv32NK6oqC0iBaD7gz4S+gs6Mpr70SUF00KnS9yQ/LHU160+ms7cK7kw2iTT
jM56wUQAJywjs5XTcGnhG04+LBYz3HAzivLmn80RQ48+e0fWp7tbGP/noz21AxeXmfvGzkW5TG7z
YK4zc7EmvlEU6cy5BUuzk/6BnJQwHVj1OwRYtelaKe2ld0763jsvFeQsW8F+CqS5Vss8Wuz7q/mO
dpji6nmMjtB3AiKDc4i0oMMPKv1eIUetqFhWG8nSLZLAIn3jUIUee/sf74X+7/gXakgyPGUj3gh6
rccc5lMdnEtnfsM/3FqcGWFkh5dz/jzDePS6WYvEisvxX4pbdzJZHjogFqR6KRt7uoW0RyNnH2bz
RE8olcbEPBg92sBYE1eXAXcf6vpOAY+qbDDhL5TyB/jp+01rAOunWuX9+m7FkCIE6nCdmHpmOTRd
aedVbUSsu3Y90SHNsTqvbyfBXTqpcO6L/AqYMneSN40NGE22Ab4qQvD34i281Lq/pSju4qZlB19H
/0StDn4x3kySr/5gvXeuApsOA8WNlN44pAjanxk8HVd3KFY7aIloHY4MD0na9ad6OLiRpRXGe47z
dBBkNYiAZRC0XDg6+sNRgm6Ohlzd9uX26fdjcIbbTXlQ83u2GKaqyLxDTjkdErGmV83gg2cQoSSX
FQyvCzUPFS8VSk5tR6yF7zz9VBoWdgocp7JFwL9pCt93IkKFvZsEgGnOsMGruMCfZ3ojyAdAUF2j
Gtd5eWy0HX73LyXekuMmjGHgQlpueFYDC38mYwSy6ENjNuyG5kXFqLqfR1G9T0eF+vKSwaoxIkPh
eh1JkDr8DD9XBuTk1YvnsnvbWFV+9/sFI7rkpW1Mht573HEtUVD81kKcMQ2fuBkiAy1nV2+Booi4
OoPObXqC+vabegLhbBQwIAN9lnn2rUWbOxWoaEzBnnSmlztkTHETPW3fElHukRdMtzKbs3oP5loY
5WylGhXcpfykMTuU8M62Xe5tVSjHNdMvrtGO8Ti80+oVDSVmXy0LGFyKzcag6pdfWT8YVsgKIi3a
XNZF7/ruTxMj4J9dWn4SUIjNAcbtyXLpGullKwCo0k0lFgGaJUCt4HJJjD9TrSwOUtdEx1X/MOFc
9KL2pXuvZPwY612+tpz1nXWl/IFevAE+T8WaCV/tg58XCgmdTXHo+auCCMajnrCz3r+7+97gmhpG
NJcqqGy4Bnb+12EDbVMv/SQUXoUtjOQ6xP57uimdudmkJcG6pqRUdAzC3NK7EoM48ASDsHOzHKbS
wOp6tOBvS1NGr4jZLH+bHxkFHXe6SC+MGclyInBpqOASrIhdYK+ti43KU2u3UMIFg3qwubxcyz8e
mYyzCCvCWW8rDnZ/4O5m2d6bLC/PU8D/1UMgMyxY5xWNqCF2d5huIGTWt7gd6qGzrmMg902NMkLe
zFgeuRFVwBmqptMWy47EAowJ9hKUpM7pS2bbmhzHIXyaz2quWZK7gcvM2gJ/h5TdrYuL+gqw0w4N
ar1A+Qd2x54Dbt7mvoCgRb4qxCiB+xcGQBGKK/vB81O0u/LwojTHRPHpTxCfIE5vJvi3+LuWCR9c
mMDn/ot3KZP/p8H7hQEG/K71rsXi7ESXaFzjDEj2PZsifOsFZqfRSmGl5CJVwa/Zo11o3H7dxHY3
EAe3MC7dVcI+IjgcB/jqU8R8GdSpQi2Q/Z8acH6WCXAw8ucEwqviF2sov8o61uB4SX375hlbX8gW
wcd6DaT0QUTS0Qyu3LfMDyJliHFPwASxGb2Ltd2ulumoTKa8WAnzj+RUnZaMvmZkcXxrCS5nqn6x
xyuXkgrPfkJSmRLML4P2jBv5nfQ8PeAYkf8VONiqknFBreh85dnJjv5QYc+UUq6RG5oiS/rF0zcp
VxwMCj8Y8l7qPbxguhiQ25ZT6uSvP4ieftsBoGnu6+Ra7pVDiukggSXTk9BrQ/+QeyLy7m47jsOQ
18YGoLX+7GZrtnKQtM+q2zkAXnU0QqokTUMSuo6vBQadLUNLLzVVZ7hAtJvQeZtxPYElmSllyI3q
o+ud05hzc0UuL55ixNZLfnfbJ0vrLq+jwkOsMMgoBhmGRw7++TdW0+994dhKttkiHv4chPlBNj+h
+csBq37llsPTOwH/P8dpHGCD69dBsQ3xSO0FXSPx7p9Bt8ZsggkA238m7dfwPHNLA/39TCx/Ocun
1vikww1DnpGwhqyvl5S5FTXK0utc2VpgiG8cV9wg+Nl2DDMfD2fNqjU/RXQb1dAPZhVSg7nuTjiv
bY1FjuW32ayzdQe6B3EkBRggevl4n5VWf0rs0+PLaF8yAiviBwZ/dr/YOQJyz/IY0/KdnS3wT5a1
WIYhTKaYuRzQeJaSQXafg8BzZpUkuo53Hg0eYdDIj6Hgu1Mv03Z8RkzmmR+TjIHN9EFcletZoQfa
Li6l1nP68A2fnPT1rMnfUt84jlGw6bcF2qhLWQTDtzJmBY4xFKpKDQpvYHLz5KGi6PichmhBMy4m
1Enc51Y5tTVka+bSoF1O+DxNg5Ty6OAvqWou6M1FuwL1g2xPOWDo37ENFmnDjXcx9M5peW5K88qW
ZygcwEkL8c7AxCt9b8D6m7ZU73daeZLiBaZr8XUGL4q26mynZGa30zzVQNoM5LoOraa9zX4qajJA
A5NOeGD9yTjiBbk77ZuC/P7Sgk4XFzzigrncerDyNcr42TyzhKeUGV0BFGUiTKOPNarybTCA4Zoq
7HdoPpYRjd4x+lSVYgXwzwVwwKLZ8wOs00RZuw+8zUcRiF7z57Ys76kHP8mUDvi3hHaqXU5efEeb
qjQIywq2nIBUg3jmSZfYgEoOeoQRKjIkkCxPgGZ4iu7mzlReN7//DMVCveeYAnqCkwOnytfNqk2k
UbIYVw268egGYOdHcx9qcs1uRqnQJDwkbI4Yl9t1gvAXQufF0Z4UC1FK7/ZDam1hDEqJmlrK1Chm
/OInkV4YHprjFyXjeectT0TMUw3zC9sl51MSgSSe4AfJzHQQKa6kPFNQ/Xf8E4Oax64H6YoUWR5n
u/Hk/cGFq64WviI/73jfbK8hxdnuFaVs+oqEGZCaxT67Sxoc5f57Q5nPhJ5ZNnrmzkAtmDhqF6/p
ErZWXH1Cvly/DHkujPUi5MZn1j/bJ2YRM4XRXR4xI1a2CCM6e5nZFJP3mm5PO87cemKAFePAEtPW
hKlIaKTzOEj1HSnv9EkgZG8zybXzD3DqC8a9DVOrSy3KJrTOTLG0E+zHW9kFeDzpj0WKMCXSmct/
HGZmcH4wzUz4AnoROyYSo4aNHhBOTF5+6tNq1Ona+uD0/ZC6fuHFEPTbdCg+wOaII3bdopSr1K0a
wrzqPNYAAGRT/FQGNl7HRt59hxBLxhCl8zEvv5z7sJgATp0IjethGnU7Pcc5yU2GF2yopama3Hd4
f+QfgzKvR7ZxMBT6eYnbow94ETWkrZD7LZL45UjcARyR1x7KiMi0pkx/G/sFxBiS4zbRGPxfV59L
WwUrzqaihTr9gY2VmO/ZxIivHlyNA9vfAKP5lmoQPSRl4qH6ePxJqUW1WskNdraLwFs3QtxFrjH1
CYy0faR8vVGg9M4NodZFXX0r5n/kWiKZmLj+4HhHmdYpGXdanjoIyDIq4mOobh2YG2aNRct8YbLt
XShSvSN4USRnpzTDBIwy1d9kHP2zlxbeul77sAPgJB3Sj0UOJkVxFH72qkYj8IxH9QpWAZ7Alq82
uehtRmKPujrrSkHCGL3235PIfnFFCc+jO4uuxQV1QEQjHRb4THFQ6BN4Jr9C/B2vko9/jyt7kPce
/7KC4d4nuteJL//wCVpQ9NmPOkvNSIDE+9ngjDb3ivSDzBcSiOXkjC2JgTqgAX09BzCU4ZBlTqeq
56oxit7kgSOuWrKiopy/8WvcmAFurzf5OpEhDbdobXS2FemRdqGo5nG7Ip84IcLgF5Yom8hvPAFs
vPWBSyDufL8yuPkMA884Z/DgdrnVYmfUC0c7/Sqr98fAfT8+TzI1KzRFeSF5QqCEXMEOieQhIF9B
jZaw8WZdz2qePsWxApecZuDXvaoJOiir6juoK3/RgAl2U6U9jWfZKQA9kKlFB/Mdm1d5Pr3kTmLQ
uomVak8i3vtu4qlV+iBYuGt0V2TTAQFs8B8IJsvWMQKW/SHEvbPgM5P7h7LkEWi6zwyPYXcOTlql
lG4kCc1ApLv3cfO7l35JnDs/lBb/JddnyQPvJhx5GJCabrV4s4uEIojN3jzNDA/d6ddVpcj74UWv
w4+fhLihBK3S8yiawsTHCehiNWfXXl7YcCKTiYYzvVsKLkOXRk0ybGidpyboJ9kf6t9N0bum94sq
Y2nUP+X4Gvkg0v43tRZ/Rk6RYRyzRMm9ozMEy3C/zaA9/G84C70O4yKKoyflkhdurjQqmyXvZarH
njsirTP+GDKWyyxFu7zvakM9dnIBrj1f1mFYi29viAP7bf3/VjlD6Iws07pNL4VBLkDbUPBRXf+D
YfSrWwyDzwNtZT1lQqdjD+OWW5SOVJYWW29YIcywcMCZCkabHwdMSdvtjWBgnSxgMXYQ6wysLs1M
vMcGUT06n7cyli7LzjEnm0hVZT4VpJl0kn3AU7vzCZ23ShtTzxPptOmIAbliZ2CJTNrVNyMjBGpf
KXQ9fdFYxu6OgAltM1i1XI0+CKG1Cg3SGutgMVW+e4ofJFawZXvqiPcKeVVi0x0HMh1Mp1H9FapF
NUV06LQ22ul8LjIToBDRq4+QK2yUYwy690UoVZ/64ZLeKx4zGHyEeWW1uAparV//ENg1aXZhSBgm
lC5mcBXh1S9jhYyIH3BXNZHpwy+m3Aira1AReMcbraOt8PwpRWL4EsozMwZgz3h/jpRLCFwIfHTt
2Y8QeMroMbr+V8aEENMwp3K9mq5EO3s38hMwHjVcWNM4uQeyEXhy4VoEWj9YFik2NlAF5MNAD4o6
VoGa4SnLA4dWOtZ5H5ziFg/MTeqE98JIFDpGBTJZwM5QcMxgqfR5xOJnDerAGKBsfCccEYMenrt0
skMmB+TVV23Cnq8rHtZyqivry4PQzMOsBeKKm+VwYNOaE7ENoQB7KI368k4PnMv57qoBYwPJdV4p
YMoedWzwJ40EpOGWZR7lJjTpmKYfmqHyigPXD38mZ0llxbz1KEJkfn9hYWOUQ7cJcgKrHPcdvWdx
0ERntu5BjsOQ0Useqc/l+64u4gfix73YkmO7IzQ3seXNAm3bPZE3h7kwrjCahv0htSmawlCUEN6M
Wy4P3fvdNmrrbSuvuB1s50bdwpWcR+MQ5m5XRiypz1PVvfsDbGmCNsPierZu4uifmDzh32kATF4h
xFGo0Nn4KBZuUFfnNyOalfXkMniDyhPV1eVWlVZYpUrMxli3aq1ji2IWWK0KhH+vQ/yDKRQsC3C1
sE916YTnIG7q4MFoumBBozF9SkmjGkE7yxI+2t4k82lWfGuAcMoqHi7JULJOLeD1VZw0rvYZtAAD
kbymK13Mh+6otjQqUzQH4f8nbPNvSeAkdFRa9O4aFDZ2AFcEUAvW9Y4hiC4wx4sCip66Stina+Ia
P4OTQyt0PNbADNyKWEB/TK82XLpp9WVy+ExbZ9ls5dLuh606r8cpoYSFuQpAlYSYQPhW3S9A2sPm
3ml88/KIcvl0cXDnp2Qsuuolsp0B5Ctc4wu5tTrXX7eqWxp5IvZRU/Jqu44Ec3y0tijA/Ab1llH+
4nZ1O976RsHr22ClKPf6PCf3tW8ReYR9JJ38Vh1TkbOB88vbusBwa5lPc733zPK+ampzZ+AFSJNa
eaHGUxz4Z+jaDtbAQBl3kNysGh0RTtmP1WxOJbjSU7+tl9aa0H2/IJHyc/BUbOnVYgoOaiLmuQKt
r0qXtrhIe/NAf6KZ0w/xVmDBu0pMtyaR3948fnWjZt2baFPaOmy26JIb4ReY262o3OSfcSIocQge
Z6x75K52YZSM87wgYyJJ15rpk+b8wsMdMlJNewC7o+LsxUEDCG647QVWJBbkQw9Dn7faXcZGoH7j
VXtsXgSyl1Ou808VrjynInEC0tb7UREPLDHK7jdTVGkUXpo/NT+w2Yp5fEKRGbbau6c7YJf8qW7/
4T8RkvG9lGAL0/IT6U5To99Gxf0Xe8ylnTx75N0DmDTPLCT81a/AsmKEplFWVVohfEwvd4N7046q
T9VisfsfV/P4COb3h+5mxc2CqQDQ+UukmBCo4mEh03usYZJxVcIf2RQkJjnv+o4WvYwk7dg7CFpm
s6U8H9h6UemvRz1gFBU6LJwQdpaykIe4NMZ2cCn3t8JyonuR45luO61vBxdaXMAEAOrye0RRynFf
Rm7RBcHJzmD0l2J+ML4bb5Lcr9YSJ/arSQ5q/fQ0gaUsAQI2sSjPD2C6FggodLisTJpnO2DgIGQx
v2d0ZKlU5hpngvNIAxlaQkNPLNOUdCxR8tyyXxqOWvR0YqRE1ApW0ZjYLx7ZXAcJTVMDr5e/Gglf
6bEdke+J0kzu88WfXXsVrm/Hul3XxO4XAPbmxZUXFVqAPhz9YFm7pLMN7XoUtq96YWyi0Sopz1qv
9V9pd33sfZfn4T0TT+TBEL/RVWIYgsP4O1ctx6GEoot5eidwFCuJD/cF0/nVS0Gt7EywmyRoO+6y
+u3zQEV66IT316Ka6ZhUvxcFQy6guIZzcjDxdBS5zyXfAZmF3SrKJhOKf3MAJefj7XjnTgbgORPn
xnyu8rFAtEV9Tz4R4jW8M3zKcfDLu7mlaPQtKSij0C3rB6Br7uP4t+3l2FO9zhXwlQyaQozjL8rJ
v7Aqc/UHPZGqSuUHHZEdNFWDCoV7VsQLced32g2+ElR4iqnsu0VyRMaKEnMg1glW0wWmRrDoshgj
mJZut3u1NlLbYxue+2WTNhsAYYfzQ7Yd4IDN32NMfqFwN58olsi75GZPuWb+SocRWF4X1jWjzs37
N31dRPlAjBlj16gtrY6SWNl7lkDfWizEtFMOfjyec4eHKkSdB88O9Uze/PqBwNOQDHq884aU9Rcm
BKO/vjSIC9aKGg0UZd56xnDEik5rmPw0z6ftShPmk0tEPOESLx7S9AD6VwYNdRc6XQdvv0ctnGZc
i3nGBwSzy0X+5qtGZGTBa/iuZwUhnaYu+GbOUGuuqbG50r28x3NYh8oFb87ZlmNrMBwqYK8jw1Zr
jeLZKOBXDCAgsBoBdHbeyoSFIgnYjKVGCrugHY0F18O17O6MWdPUhCjtKlukpFJvefhvqHGUnNri
y3ocH4BzD/sTyMZWBIIdYO2OGzFlOCfAFiX6vQEyqPtit5uuf4GP1gEFxsTX/lPPjmZDAFwc8mNG
21lKNWWe2SfIxyZBKQzWzY7e2KoWParrrAys8TOv9j5BBu0d5Jf13M+KldkW1ASJj58I8jn48nnR
/fry9GzoCmXbL7ZMSwETVBXAKeGHFHihiFygO5F/m6aLGJT9g6qzZS1CMFwAFM3vLVrYC8Y19UkC
WLwKhcy0FUGtsDV50IJ++Tg5s7T2QS69hwlR9ZYZ11jl1akiTk5vs0Jak/Ud9Jo5GmH2QvF0EiKe
GHLeC8VqIWtcdE4bJReuAU2eobVhHJcoOlqQRmbsNIxLn2fh0InXvX7IBPS7rXM/E0H2ivYqc60W
BDTktLx7OtFXRp9QwzThCdwl1eJh2iOV0zS5AfFUXvg4khqzteDz7EU2V64eAEGL+T+SIE93F4nU
GyL6NvZgNTndH1BzZQN+XfHy2Fz0MoaxQ6RaXevmInrT8gV7eywSVyVqQKA2Yy4NXEEMzeyYV5zw
/05vSA13Cguap0UEwPaErUQvOyEnUgTRzSOPpyphjafaZvSDn5Lyz/iSI/RQG0cp/ZcOa5bs/4pb
9lUi9FsDAhUBtg9tnR1N+Ki+f60wgFMyuCYGRrO5cB3s4NxAsVa9EsbqozzIH2/YC4PXqIQWkD2n
yWv3GE5WjTWRFT3j/mEOWe8oZ8WtyxyHVeh+qzRt2VGHxjn4XwhcDYiE8P7UD5MkRZYNSckAH2OZ
7h2/qLkj+d8QdGp4qlF7ZoUPbYCQ9dNlIMwfqUqJ2TOsjUE4roK8FsbbBSGD74AxizfnIHI+B0mc
9dMnG+V5rYxTjjeEhCnCDhVTc353j1at8YHkTZyTZIKKmR69Erx964os2CuZCJOtmY/pN6TPwI1V
e7oyX71aoPWdccLP8HuEuzq+NX4p3HTS4wKLsmh0rDF+j3FO+SkPB9gyZdZUJzX9hyAO6D5+IqsD
VwpJxF6ZoUob45kfkqm6SvlWyGiQFN5zzXuiIChdn5ijKHXohdzlT8xjC7FR3McXEBENjiUaxpPY
vjZFXl9jrFJqr4wl1dHiwVJ5KuarKp0IeLLmBQoR+IJnTJxtKRCQwAi4seMTozkX9htA7RqIx1kv
62g7jL/Q+ZDxXhnrplYp1o7qobGiT54sV/23eZNQ6u5rdWtN0mZd3IZYKLjzGF/FYVHPGfIYpODp
D7EOP61cC8OR96pXQEMH68uUU3SX7VMG8Y90suDA1ZjJ4uhGSa/3Wii8yDtP/KmaBUXL6ZOScu2X
DSo6v3K4boAfwwx3rSgwbCgB+BLb6zNrCo2KCpWQBlFlPkmekC3ANAwjSyzx7jUHzCCz9fc8ZvVe
93PGdyLRM1a4uLRunCbIGv3xc62hznAar5WQRVhGVc17t3ta8fkqg28mcoy2ANXPK+twVdQ6JPD+
nmQn9r0yUe+NW6ki4n49m7g1kyPNAI2RBDpLKyCrxjJ184ZMjfFdRD2Aa/PPZxQxavLgovyu5ouZ
8pbk59+ys8fygA2G2+PjYCjgNSIOVerQMhABGIvHzCG+i+sfR3/jTr0B6/QpsJU2riHX90qk5m0T
6Ol5pa0T+jsVqFOkKrlvv95wP7nimBoeiRvlkkWg/aRfV4Pbnzgcsui1fyDtk9bBli6jHemHlhNt
xLAMOwZlqwV1D3FsGR8r3NHQGHqkOcoAK6geLvixfPxwbh4PXSidZXKT0wt5yWcNmLHZqN7/Drcw
KbZMaZOBmmudZOQQJrgdglzZkV/Kma4hqRcIphAGxikOiGr1c2B+uCCVZpQpl5wsUIAyh8EqNDxr
OBhQjWAEbEt+vWbxv5G5Kpyr9n3C1EzbvjspbBrlEZYs+A2Z09NE5v8S3c4LeYhby3bqBDzBKlX3
zhpbxFju+kuVBbmgQTTNbpq1ZN51t40OSpyq9TV3RL+V8qoR9HExJOY+TkLhlv1Sf3Jggv95vYwf
et09Cq2fLMl06UnhRfT4/d2ybCIO6w+OdOU+axUXGUGkex11l0EsCN9LJQ2GR3L00QfVcNqmQRGh
4cCp+iT7vO6djFf+VX2DhHVudTbXppIapbdWd8J8Cs4BosnYCi6rnI0CxM48qcG9tjd3scLFd8lT
OLGKgFmZzcRvKCcBjS9bAA/I716p7hDSE1NNZlVlK+f541QDdsQSLBIv/Z4O2b2UwALvXWlRZynI
OA7Qys/+lEBiya7hzoawrxL+PSWB/16vIXN5Skr4Qxv2dZA9EGnm30fCz16Wtqo6GUf64cTYzzpQ
5endmohAqwhCby8DxMDeVQRbj9KjS7bq63ebf1PpIZ13gp7OAtFEOI1GiK3f0visfiRQWrHdL/v3
BaphhYP6gzgTLjjWJqS9E5qT8X5h3l640KtoV5ttuQKZdlSVB48V1mCTWyNi1nbxon7BXPPUWsq1
ts6o63u1f9SXL13WZDydWuGu+Uy+NZVF255XU9Rx5cEW320WjmXqO8TUBQ43syvxMKbISxdEKCMz
Tlwj2mE5vHejuH4PI9kzI2LMCAeFVtBm1hNCHN6p4M2ycdzhomoIAyJEg/dKRbYM+cR3Ye33pzh7
b5OVXMeKNK804HHVkbilOCgJlkzB6sdxX8JxDOc4xwqSKkVquG8Ecydsi80EVojUNrBbDMkC8a/S
ZbXBGuN+bkw0nZDnM8/hY5Tlr/IrObLSH8+9nr+InRmkpvnF6gkm6ihzqnmuEyKK+K+KKnko4Gum
HoTXIpk8Zth/DG/QG3en1NahEGNigp/y4K/o+tSe5y9xN6QVyAxclBZi6BND8NT9l3lRBFqYMmf6
LZefRR8nQx61JGJHp2+nYsJn3DfecONm+SksTYgyO3x5BuJ3tAqFWEidVBgRm+LnGkRdmt4/rBMs
OVYTk58WIXXQwHks1d7hFS57NVndzppwY/FRZF73ucOI2mI+NhHSLUbVZWdG/l2+krxNRtxwt5Gp
Kehs40gM/pVJwD5+SuWXHMK1Jjm1AVVtMaty1Uvyxl7YBGhvMKw3Gp2azX5T6DSaxQXFeI6toDxk
LYftduAkA+exVkPGFxev9Fbsbvie3a1dMTe5QcaHr+cPxsbhC0/Fx0Vy+AmVa31+8GW/2LajAkZP
L/iCl1NGvf0JUc3nKZf5+EmsT60SwvTizmt8OflnkzkHJM5GLdwKALQ+fZNSpDJUeKslQLsYZ/rX
qITvmP/d2iF4dZvl/9ynrml4M1Hfc6vp3ND0hfapzsqY2WRWIUj79FYEcXwOn+jiWFqjOmAOIFS/
C2Y4PKZSsjv69xGEtM55BsYD9/7QlttmAe11iTghQRoRH7K8yEZvJmLCyCNkjaLvzOD4MBB3o3tj
dTJXsk5KrNkzKWow44WdOjVIv5Cy7lKriZYvwmCu+KOV1Ti2ePwjxKWJxtl4+pX6sNLgYB0R/T5+
IfA5qb+Ok+uEtZpMeUVpoXHozdRSZbfRmyL4pl8gTqrlS1PQ1mB7tZqsRCEEZBM3csGMIb/yI+jn
av6h5DHy4P+zch8XZUNoTwO8KaY1qTV2F0E99mOCeXy9D3CEAY/azRp72tsStwWlM26VHwlHXgPH
6Dg+GTE3lHJvvhKDcj7Yij8yvuQzYyoJBp19rwpm/K6Qk3C3MnXs6W/hEJTTs8gWbceMYR5awhtD
ICawQFcQ0la7H6s+gXmS0p8BO72r+Xx4YAfsmKpcwKlPtnEvBOfeW2G7l3FbOAs0093A+/s5Fgwn
lXhhb0BSOAT+WE+vKI+bYobqInV5DF8RdbBQ+VcdYpllDPuInhOgYW63awWZ5rigZGEf+XgI6zru
feXEw+HyAIxNzyhoZhK6B6U+WtpL6hl5Zh7nNT5MtY8S8ytzfpR21LRT5xzXekj8N8SIPCWwGn3e
b7ECyeE/SvK+ZS6iMnWXdsw1D9SVSRAgNp604VWclma1R7A1zO7UxhXi+FDslPtdnPYn98gRpgq5
WpNinXoHnFqOnZFh4kFRf5LADPEjDrrjhRWqLT+tIb56LNJV01Ud0JU9UkfT9BtiABE06mt1e0D0
K31VcpIOQoA/DDPugZuUOpEWokDrRbKbZpWC/ryJUI4k6RPK3Ewt6yZKRH8IJFmRkKnqblXA+DXl
p32crTCWZNK/3clswNB7UtUrEpD37LPZZTuvxMYEPt9L0owx3i7W5eK6U06AOhdCwKuv48mTldb0
s87rrs0sQThMfelNJv8Nk7pKiSIl/AayGrY87XBgoJ1qobguBXh4ldf3udGVETef8jKKIv8S6D7x
8PAanQ+C7dk0d7eupe2BcqsYC+pcPUX7spXEwaKmSsH6ZJrqnGe9pegDHCDOGRd2tPYX0TEUjPis
nKOZGJHm2kCYUKfcqURUsS/vNC6PBZTOAeQJLHLn4232tCDbKbA7VM/r6cnLsgfNDvtPUqmVz+ED
YDvFqPiqe41YCqVKHZtnGFUJxYIIE//nbvHA/dEGdHmFL6wOHPMOPokeQMsgfICRI17pkP0NhdLZ
YEqXi2hfHGUVm91Usd/C6Vo3EXq4vtvWzQiTnMx5owzPwfWLgZoA3FU7vXJJlsgCSCHJe5OIg2x1
kU2hV4r9UeGNdGzoUbRgN+nXuFWig36cNBtWT2ueC8BGtP3AOeVQfiIC04bGVwT2p6LIjtch1Cj4
jTxzOzH72R4EabzH8yGEgDwOruQmp9jD8/9Jwyqb231UiuJEQuIg1QhbDy0rxqFBqoejbAfYJUV9
0UWVpXNXo5FtnaJHg1fAN2urFu81usWdhHAlJSrCiQjMlQwUWqA+BvnbVEvtC+lCAk5u76VJe7oq
XcJROvsa6/CnetESCkDDLIqbL46676Z56bjMRSUxUPNrh53joN1FnDgYc2YNp3GEYiVXwOnDULGs
vHweJ2BNqf2tuC+VoqKUAUfRI4GlLAsdLWJALLnI0mAymOuJOR0sJIIw19nwTScLBjecqBxV6abo
5FNwDu8b5VR8pagVmCuPLLrdARCp6nUK09wufTA3l2Al73/13C/G8+iaF/QOL5koKUcZNXy1PsPr
gTwLylGxUeRnjDuaCVcQ+GVLNyy/gdn7ud2lQfqOvzFLneKz5gU88vRDXSfEkDxxveTpBKlCSzUZ
VixeqsQaaHtZ7b1jIgkfDV/WG+JrIzvbF5HcRbAtComHkYak6N9IsKgeW/T2GMVj1Ca/wsurN3xE
Tg8vsVegbvEgmssGFwcLUk+girdphBG9YkAldFes7Ch36C1C0g9N7wdILG1b6esAQ7KcCT7oPloP
8H4pa30vqqZeEc/6y2TwEf/vdUGZXAoVZCtOwnUg5TemFqaWphipHGY+e1cbChczN/t2USsonPEL
izGwuiugLAB6xulFjSMDkWUT7BIb6rD0v2w9jgUWfSE/bKR3RDsDTm8Kkbh1+g5eNkfaSqUp1iKn
JilKypgDWodRvTXQ2FDaNid0I45Y8rLhQLsxiy6i2fLlw5/SolI7SOQRjnWOva/4sCTZwI99QoFg
hVHO3OpmbPcqpUR652qwTHgVCY110NKkRt/7s/WNm4UPUDQiz4xxa/wDsi22ixhM0yKcPyfjcMIa
4CGZvsNLSXc0bO/z3ueJhgYn0sxyIYQqYrAxGCQDxVOX85gBhoOtcoiTkvt2oMH1Oco6rGBTgWsz
GuSVw6a81Rgjq7UqfhI48BsCG5Wd377EOw5jCYFq4kR1pFtQ4uqpmEwn21V866WdBmVAk32s2XFH
xdtUeMDYNCI+BKCOAXrJghvJjKp0zlo0uZLmmtJlVQFdKoN3Y7r9/qoJUdgPdzorqslNJ+vRY5sq
arR5csJd4h6LYTM/iyY94sf9gUntn4fslBqqiY2L2qpcxlcHbzlphmDOTf8KcXsqj9gBMzIIUUph
j+88BPnhvaFu706RGMCqXe4Yc4ozAES4JKj3fHyKcsjW8ZjMkcJIKku08CBOpXeV+zntGzIe56Fs
P/kyfMIzmKwGLislIkg2r/auhqE4ylyvV/Nz6U/0DAWuCc95REVZXDfWxHJr0ioqyep4uDs8DYMu
NzE7Rd/7bE5YFBuAtyTr844w81T584EUTe2nGCUT9QBs0GJNPHdWJl0/iygQ9qcpglIS+ZDswJJR
OvW0UHPp9neXVqYpf7KM9jFIvUf34M5bbWswtJTifGZ/V+hCH7OVtgaOfDShrEbKtr89LFQ9ciCp
B9Q8qNR59VzSYO4Cwz/Ky4EvQR9rpzyCzII66PWvfXNBCS92Cf96HBcyKYEfNiE+SB1kDtGAawpM
4a0vbliBxhCF6IHVduXriRf0pAooa+xGw3j0FPiE2psFzx669FDX9oi1kdiI26U/3y3jiqnW3RyL
VKW6oIlmU0sYvs5QEmUp++YZFLl/pPio6WPNn01i/AN6SnhwIo1aJvBDT3/1MzBzfS2RoLjXpXXi
IazRm12NAtRvAS2w8cXsrDjvIgdrD2k6ea5n2qdEAlPbFpyZmGdnATo4G07bscDKQBSrtyU0SeM2
yZVN0wsmy1uwV87UxGl6wjO3yAQJOccN1f+0dIJQiFEu3u2PL60AYvXRT110M4/Skd6aajj3BSvm
SSNkp3WZJiDqKTQXHnW8lbKKbusBxclF9F6q5lU+9WdZcK/UQbf4hOFwBKUujVPCgop65GPqtgyy
kD0cXIgJMNsENEftbOLJ37ZziD/W74jbVQUMU0AAIVX9B66Wtp79lM72lHSZQ808SZ2njcfwLIi0
ZH49yqKckKthFGaVyZvRb3M9OgfNL8af92B8JjdNJhfvr+9WKlwpLe1F8k6s6qjbWdnRI8jfC6KL
jmPg2vAnE1lmeh8M/8Yui70slDjBWUOoLeoK3f8Hqg2YDONpk8Ll147f0l1KivL7cm2zWea3mmfx
0JpLq7p2cYEHwVyLyCOQsE76MbmeJ6LU0Ki3Eq6rAoI9s0/TAYK07j1u46v4zcp1nHjbL8fjIr0G
4hNwtQmlpumQmWaYQa44CaXoPMmRVhRUpTHD3d7TYTV6QN7mmnAx5Byhewr4MpWuvA1FEQ6LYKG2
qNrl1CB8jpG1FuBk6vJeRBST1aXRCKdW1dv361XgAHl2n/1nA2T/1UMUgSHk20nJxRZ66+TXo1JX
N5rY1o9hJ1q/d+lUfH0BcYXEquTDhvDtliskdgYTWeV1SpCb0QWKeOSJ/TOqIWPCZTbXyNuKduDU
+hzPIA6FqlMKKJF7ocoU7xoiWP/N9rwDjymaVhnfWJvUjs+sas46NcokT5dDojc6sZ9mk4UQ4MK1
DZPUpkcKRVQVNrJhG7E8R+o4Ej4gsGktYWNa7zjjSlcDBjnONfq92qGZZMNOxFrow2kXlS4ABaaQ
0Iycft5AfZ0vcWXnlyBaSJ41l+wrIAVtQWclVHTuIdTQudHh0RSlxq23v83EUoOGLVfVL7oBMEWW
eEcSPM4XYANxKaCNDjREFKKg5fmYJu2d+IMc0LWF89zqeeNkue6UJ6M9GyUD3JHINX6seDwhCCem
CY2QRxA//LShG5lBRYC2MFsPPo/Qut7Hheg8RY9E7yyD4GqxQOF+cIsr9z0kvdv/3fNgvQE0OXrt
Qgi+IFEXLJupho+v4KUJx9hA5UAx7UtRP3TmmpezMqBgxBH54jw2zGr5yUoW8raKUkMdTZz49Lyz
DWbIh445u1Q88o6iiEAlxTWrwhSZrE5TCljmdBRq3PrzoLrhMRAnWMi0S87rRAXpPpbJKh19N/mI
+sZ+LTJ4sCOPNWtb42HL8xXHDXVyXHvgXdN4JvV3FC+QQZEwDthd8nBCiJ/ENjOr3HsV2kGchQPr
2U/bsH9zMFuMJkeuVI0Cl7RqeOj+/Izl+tHySXXQDnKZkpJ6aH57lXSWuR9CUIQXq5JXK8X4vIpv
tbRnIZR6oUGjqwfLWhss+M4c4AQPfuoQZmME83rP7oS39NQgkKrvblWx16BYyuJV4Q4Xv33rGyw6
6YdrMxbqghazAUxO/ZSiPPPZSp5WgGBZLHhCOsdKRpKYVT7Ed+KQytsF5fSSMk8EQiJMHnPAUu2R
YGnMjkPs9RuzVr5Oi/laa2P7CWS0+o56xUaMENg7g1pjiTL+pZrbObs94jHT6O+K+bAh9f9uOw69
sQXDZHpKIIqFksnNWQHITODQAqmfJbZI1ocjTT76bcelmix18IIZ/KBl/KVU9EFHz42bEwh8dMKB
Z6VqU436uW0z1hk+szGc/6OJDC95HosNBSPO0UCnCl18ctJQFLtr9w7o1Lbn8ObwqAKja1kzO0VY
MpN8xSWxq206LbH7AJBs90P46ZHrQwDcXBRrvKFgxX4MsHyZKT9u9vW62DX/y0llSrx1W6JBT8ic
kXMVaRJuy3Y5JahUo8iP23lemeeIeTR7W8Rwnh+WaRSysdE+z/FmiKB3iXrg/Txrl13bsfwKC6CW
Z7xFXWlHeuY6YwxpipgTLIfUSLypRBUcKqwWe6nT2RTfiR3I8RXRslfvaXo5ZZOyoR3SzeHh1d1e
kyy6ZRHw9d5dzGXkWW9bQ5cxUqtv8qLFLm7Gu0jNRg7P29mIuT3Cvuoat2w3sbx4ZPBGxvrC5ODj
Rir+U9kR3sUMQ9fzx9/trwEXxSL4wIsz9OsslITqzl05mRTq6+EjlTeLmhIVB4rJKMUQ6aN/sfUS
+AH8SxvHyh0NP/e1G8ZJLMLncAcYYIxQqPoHZLFzJL0aVEKk9c8/UojIrtYcStoyzmjM+L0TYXW9
dfsVxzuvn6TPb5snK3Qo/Puxx2EKfIdJQxQuJYwUG/HwWnyFyIfXXQjJEVDeN31hs70mq2e06AUW
X/LIO4BBlb4Xc0WffwxvbnfETY2CUuYmhPH05USHUeKXK6ZM5yV9dGN4pLzlE3IVWXPDUnhA6Jg/
skIZ2Uk0uavsqSinpA9RLD73vAIIjqMONAJOAckd+4I3/Im3k+BrM8Y4XfjJAZAKM8tmmQlu85Q9
sxkFqJQ95Fxp01fUm1v4WCgjDH83yBdPp2S2yFBuEBDghr+lQLYAx3Io/3qfMp8iL2/TMw/4H3ZK
5w16TgZG9qenuj2QpnNFZrxSZ+aYN3Gqr9MG6bKDXfCtvyWxIu9FqoTRcj8ZskjhL5/uqJw9u7md
RN7CuSRHtLUSPTh8KLTiH5U+A1P8ocw1nPAFwBOft0BluMdyTF3SD+878spgLuJSyURc6Cci6UJK
FPciIw/u3bjTzrB8AVqQGMKLkyblS/fUhV1kUr4au71Ne7b/unWJAuWQZVd7dPdgsWMC1uiQwvqX
6UYBhBb0OgL1oRWGjhUdBp7di6QHpFGOuF64P0mZCYGfRogA+3KGnGtld/1FWSPHdEoWFQkXaEDi
CS6OJ/B01E4gNoyhqFfT3O0VfWkadBmi2e59KmO+b+/o701OPh67LeX8ODX4uuv1mJJFyLwNk79Y
iAVUckGIDW97WCS5WmXNaEGWjJlU/a+qkXIYaxCZRyTFcW5JlJPFb12ocw2Z+TbTB55Ip7BR0U3/
mvVhsk/rr11eyo4J4nioXs5h0994xaVaZnbbWEUE0hYRVeJjmyEsfhf4rSFTJRiPBouWG8uBYJe6
ql2CQ71frCu7EVbWfeeIeRPoOcwcq7QkhElrYI5ifgHvfKGt+B9RHm9dA/hZ5QlUxZGxgmwXjjDQ
Ae0tdEG8VJBPRRM8o1MGsmEHfeapPodncFU+QYIu7f2xLEbj9bUAX4Rb1w7z7p7yQXCU95C+EVxF
3hiYj8ph2RK7tChj83z2sJEVxRnXu+ULnj7TdDUwMw/aQ37V465e8cD9KVeyv+f1iw8bNBz2lv13
4zzBV/KUEX7uL4IVvns4LTGdQdHkjIL7WSGuVugxC/xbaszUHpYu24rB6/H/nNwCHGDiaUZJZtQE
RR8+HYXP10oFe+B7CfFh3yskyhJ9OfvkpD05X6vp/m1/ISPUU4xpEjH2Xb+5LJNDp+IGfyIMJ9nT
YOzRgbVUUZY8jq9qd86maKH58bYJSNPh7Xz6sNt4LJ0aVqkGUFgKcVEOG5kaoqOCGjU4vQwQCCRy
lqlJIyl/SkhjUSQrcXy6TRfcOQ/WetKeyXgXKZgQYJ/ioI5SnQLVc/LHucY9PmgNtF76TnXg8xOn
aCStiY+mZPJ+FVm4LmIARtLIw1WtMIR8NfFdWVd7w5VffodDGe2l9sap86xmJRdAVE4WLOcVZyKA
ErLTN/eBnpxHd2xHcIXABSkgmjQr0nO9JyXu046L1hAk40jp5NAum5rhW9/gXSKZHZBeWtFx6rma
w6GjeCvjrCsLKUD26M4Bo4HmDg50PMUKV3pxMz1lv1eqg9yJsofF+6NSIPDOMR/RaygsmSQsKhq0
FdR3y/xob5NnFvBVCDK3XsUTd9xJNZdj2l+AgM8FwzySpfEzuM2SctpWwRL4mY5TLSaOUvyUzOLq
A4znsKRe+sm+p6Bw4XnPT46gDskDdnva9ajA3mvmN+w/2myL9a2M+ZGqSxUr2I+7qZglm0dLe7Cf
fa8EcJgri9LoCC1SX6Sehg556BwbtuIrCxkvFzYra6hZf4H+Sd5zn4wL89jC41NlSTjd1b9kcS8t
+xbQm9pashET04pwzVv7z4m60klL5G9MrBcVlLvDzRKFugCAE4DtSKM6ew/HCt9FZoeETl5Aar+9
7d6Ll/qYLZRlZVg06vTbzBKUwTJY6FBet9vxEYx7IjkqJaFNVrwAnbU991IYGrd2UIjsFvI22ArF
ItKEdxqzP1UIcLuNktEOhNCyD1A+B0g7ZeER3AKAM/LTtxzPmwzWlclbHB1qEcYofLdb6GfgQBQj
5S9ldSNNAnmDxcvLFQoOq9tQdactiUCuL/tXNQQ0eWnGc/XDo4grczoVu+QmIV2Gl6GUE4Ani3rV
9HfACaqh9O/qGr/eI+4kYVE8PlfZdNcW4v4/RKWhZJVUK70YbGs8cNH51IpU09m1DsRmHHlWcvpB
AEXNoaaM303mhUAogQpa4r5mJ8th4zmZG32hqPUtHCUsf7a5UiQOqjy5A6t70l7IGVTHzze/SjbY
kx78E7VGj2jRcyi6YmWNjID6jdVqorndsKwLTrgM76eKe0IRr/sEKCJ8ldS4yJeWfacWe4x9r645
OQqC3YRBHzDOIwOjiLIvS7FQP4/kR5Tty54HMRTEPEOWlWcVzh9zLUfziJ3q9EwkRRDR51+hBSSL
mUKdmrklt6FcOEjfsnQeMoRmLPA9v+cCoMhcR8qQleNklRhLZnn5hXdhDN3HbK2MLZ/46XNcfhz+
ksCCD4jgXvml/1TTx3UPlBWwaML2EYwcyQpLh9gmRi8BY3keEssX9kEh2Y3KNcUkpmx+slpIYfX6
STqAWta9pJHK/CSjderqfp6wT9AkmhUQ0FoFz4C7F14Q7W9X8nCVySNGhoHUAEVXCvGNM8TErRlq
XJJbqrT8HAevLEbUI2BJhdgdIm7TGc34xlZkUz/gArzQXYcbX4dnX3ac5kUdWOliw3KX73behDNH
sWDh4IwVpA9L4FsiqUtpCxxlsYqzAe23EwA6aMSPwN4lqA2XIo/rsHk+sCb883vO7m4JtVwTov4j
/SsiTO+5WjNEy/5/Hvyvr4rvg5GXeSIpWSzdaBUGfFQEnYYh+vzrdbDVKGpi90LHkKS/SA72+3tq
IVHONP03EEvvuBSDV7DOps1gRyHj+f6bgea8M0Mu88IyVO3eBCzZXJKD1a95Jw+nH84CRK58Pxmh
g+qIEfR5g7/rX6PjYfeCeYAJZdyLUT4sFIfhcUXAloE/v2sgOFQASldXKsFlEZH5vX4XTbgG9g7O
bk0Y5MAxJKNEps+WxiMOLsadp+XzHXvYSZT2vgpO/FNGUSRalAJ3Ww8pr99L2wrHfZPXnE5fohl5
MQyc3Dy5R7CZLedJABH4VI/wB3I1m+SpYNRPlDebcN+rcOnqL+Lplu4tNA74UOel38pczvsa0//p
QbG40/e9+GoH4UTbjU/hUESx+9GPRw0beAvKT0YP3IbwgdCpiE75tYJ9ANmFFvO+9NLY/JYzjpB7
VvaGAQMeicXDCfAhr934FeawnXirnfcBJDqwd6fAbodOPYUJPcHh9/f6dLVLfHollVw4lX91CS29
o3P+Rr9ZhuunlkygpRCEnyFJjtslWBHTr8YXilUN6FOcoHrGiez/XzepNwYLbTv0jFqP1nshHSqG
5jitcEDyrd/QQpMKF/IX84i6IZOL+uNCm9ojoYE5RXiPtGMs/ZPA/SetPVkkMZ5Ob38zfPHDiUnm
YTsNgHjghP0QcPjJ4/QzqK6NTywfx7CES3vX/VbBQ2XG0X5UqV6gkLMnzh+UjpwhmUfC4BVeKZiD
OBTjZ9cgAerKcE3vlP7H2mw70QplFmhZ0WEjkix7ZrXoj0f4GkQnYTPR7DrC41WNcUkAD1f08HsH
te7Mp2oDBAKV/8ouBKUo4yL8M+T3rU5ICVJeS0gIzoz2gyklI+bJZrYj6AiGVBilFgBbWB/nrwD1
w9aZgURs/iyiXR187pMzNymnXcknx8wpyqBcvpnauLv7zj5gQ2CPPnqU79+ccHWXODhjopxaiRpV
r+vW5oSnh4I3Y9istHbIESk12Hoa+D5z2QV8igQbZ+EgqUaphc0kfov2Nw3va8geRbBP2nsQuay6
k2NHVY0IuShJV5rFpe/2EZHOX5wPgcMODNO6XdG5v+6QQpdT3ggtgpvqyQXuIZVagg1W+fS5UHl/
O4oyVEbGH5CvcqhDr7b2auFs2WZL/Li/v1faR70X8XZ8ZT7kgjZPYKzmjzaX5v200Us7g8vvYNUW
Flqhk+kr3RO3FXGM53h1YWi4rCccTXz0Z14D9FsgHaAGkD+Mn4brPHp5KvbRYhjgYyWrYcitKLBE
G4KRk1x2pxtA/nPSkHc9Ljyi6EOaoTi7yuk4B2y2qBHKdxk2GTPMQwcmaJ3pvnlmzSDvqse5pH6B
jS9JkGwL3xZ8kV/ed/q2G4ltCIGIk2WRq0/uDYSSMhksp0ZNMDYaaUzFetPRJ3Y3TdGtl6OyZ7Io
C0pTUQnlSN2k77vJI+vfwg5bkFcz25uxZvq1W+NDFlrljrwBx8AZnbweOJRf5nrxgBH+m/iMAZBR
Crhb1lNunCsyo4Qbk2ARq2awluOE0sbHZhFbTisyyGo5aQfVEIu75SnSUzwENwGsJCXW6O9E6DuP
D/VDz2YkHKPk7gU7H5j+jOe225e06xqLKXI/1JB3YJLvXb/fVdRESOjPFPK6gcWnjfBdAfNC3CWi
K1AMjsRRUbEnLH85ig/MOU5cD/7g8YhbISvGBNwogiVa7dtKZdPlFhqneaGTqcowBdX+tJ48d1Ik
t+yfU9b7SWsNFpUrKkcDNNHy9g7oAHh4L3YhXf+utXWOUxuQO+wbDc5XYM3uvEKKMP/ciTpzE6iJ
YdbLmQ/dHOGDf3xYMIPHP4iUZIAHwPSFXtiL99WdDBkjwAQXHKyOamtCgXGcUp+S7XDUsEdQ+bip
HD3tTBWkJV2jyZqI7ByuYeTm5l6719M6NKy1l6UJ8tIxesar35hjBqRfWEcrF8qt5PDN25Lfg/ur
ofh6nxS1vcSWM0bSnp6F3PZ5/kMG1EyDkA7B1QdkUx2vJRTZHpTO67Y/XWvFM0NHLgnOT30cDlPX
FkAhCPYDz9YoV3Yta0wirk1ZD5UU5tz+gG9lgX8Abv9SSffZ5zXepyMNdg4ucO8MPiI24P70bGL+
5VKSEteJZlYY3azdqzT3Ux1vgApKVz3+0/6jPk+GdEktJuoljIvauyH2uQQt4oWkhap19OzFPsCJ
FuZpNKmDIw07OITHsx+XB3mbTgHmrJfTHPmY1/dcTGtWpZzrw5xAN5W1dIA4kJr88xyo2sRskveA
yT9lQeFPgj07iPf/jkvCUnrW6S4DQsvttzCn/lgQ7Z2rWn286TtB/U5Y0633QtajAoOdUZw7Z86B
oIr82xiBrNcqGt6OSq8U0fBtj5SuAgdFstBBRK8/cm2iPh9eFeihWXd1Q/3XQA/Iuz2wgkWNJs7V
GFSNcZTBPWi+Vgp4MFZuaY6m6Dll+voavpUr/PBWtsSPRoxQ/G92RaeX1+rJDO/7jgY4iLN96N/Y
LY4amNjC/GnTTJheW1t7sqRW2KSkrGAkK7bPyIC+bht6Aui7OwZMhGL7T7YG6s4F1NbRenLXYL+L
NbYyKZ1bbSp9lxyhDQwOKWGRNIbnEYMhvWzdJ27hgphNYNscMaYISQVIURl/ngO4hIR5R2m/YTYl
dStAmv0WPYOrupVTKC9UdaUhK6ClMWhE9XSLgBaOCUU1gJcZAQ56/jU6mHNPDASMM5q4vXSMbW3t
Juo9maXpE1RPXw24EzQPv+sOF2vhujkU8H3gmOqflhxp9Pa9thxjek0mSiiOBgODKls/MZyo2jYr
aH1+Mo/kh/rZs9xhFrQKdEgj1T9Fz7MR7Q4NGhCA+RAKHzYXnp7dp1hmEbHZ3PuBBQb5rjN5ogKp
VvG+cgAxtIlcvJLcfAx9Yl0RtpNhxawnuuOAlKUfI06hetBD+9jjc7av5UrRJCnbBGrFoR8986S9
ZmlFNIMALWx89HGxCiS0z1vYLpDBTnCD3HZWOHbwCRCZ5duSlQoeuCHkdbszXcHofG/7k7nVERdT
RO+yLDE2k2qcyFYX7thmTLgvwTn882bjnYsz7+E+KlpU3X78J/SjD55nZfbGN3MqakrroTQyPD1n
/+W+5F/oq/tu8KRHlCnN3CEDbHW92UtrmrZIgnKBEd/d3RyRzKGAMWKIZODsYVpT3PhUdleCwujU
YGyVcC/U1yCq0mDuHc9Qc2yX7QY+rYPFkyvBHGI4Uqfx6muJSrwH7bl5swtef6bXKW3fqV1Bd9xm
doPyAY/eskAggn7UlsD03JE2vFFQ/48pTHp5hmjMxCBZpHcAqfnLfV9u1kkgG9Z/zk3Nmc5wZAFP
wV3d/r8FfL95YOXd0fApX8BOm83WB5Jd+m0budPWNfbX0iuyR8vtixg2nO30yoxusrtNtA1oKIyi
bqF4R8w+N/qKWhGrJVGskBsk0c/bTWXDijfk3T2i9dCj6wwYhmLFuk09m4A+/Kpa0cgdknpgWG3S
VOEO7PJFcJD/EvJQx5OFrfjfJBFXG2AbshyTHvdepVxwW6NbR7wNRuOj6ih3G5AGvGU7Uw2VUbRM
VWKqplAn5McyZvJTIsTpL22onOvnDMvbyGkuxhtEkmSMRZBLNQdLyixT/wAsNDIm9mMe0poKlr76
LbtVlmDTy2OsfIS5mDeZqYEbIqdVoWm+TZt71qgoYRA4CtyqBwSP8ETB6KZ5wwbGg3JuBlnszsnG
g1mmoNbvnhrc/JKEBRSYeqczBpSB80gWdg7sXMPOa0ow8eeFfim3MW2OU4id53S/WpvBQ2Av/uaU
72THz/nxJUslHsuBk7lVbZUNcQ/9c9TElbX3q0OfNy6i8wno3KKeuXJro6j+me+b9RpMRzwNKzbg
mg5OnMnvMzDTiepOcJ7Z1d4bPzp5mBWJtYJSlm+S1aZ/WLgdcvumybn9Lo55x2j+gsk4h1zKpmHQ
FoS1KNJ2U5DwTmrzTqdCvMSdXs0l0WL66V+ES9pJQUZtxdQbc4lZln4a/xrEYkNbnPFmIskLNTNG
Xq6VVSq8RDP1/ER9lzdcI8HaKoOkdMU3e1WUexuvw6lm1lrcHvgfDty+7XR4ce37qy6o3pksRJGJ
f1fMezR4G3H4MOUSF7toxeflvBjPaIIsFrbVeEeJPwVdHHbK73hpNg9+j6cKCvsaIQsvmouoj2/j
lfieQZINm+VskV9gXF4usO0mquW1vgXDuZHLLb/W3P0bkVAC6ZYIBZgMyBbfQdm0pVmMHRGkLIma
NISz9D+geP89vmrqRpICjFVEXjlruWya5YMT528LJf8JWk+LE7XXmIKnk3/tmhmUzS9ezj6ME5oP
W+wS3iscal8BpW++GZAbcMiLfYHhG/rM8sBphVvpDTlJqIu0zxcR5k24UngzvC990ZVklCjVkG7W
cN7uPxJiQWWjEN471VRYaITp/OmFMgoVRLSrmp/G7WnSK+EEuPBDt9rt86HxvB3v1zisSwu6LHj/
OUXT8yieYNViKHi9TNMa/p0drodByznaEiRbYcSIB/pxmucT5DKCNT5Zr90W2skEJ4R4VonmcxjF
bAhhyap8jkVFWD4zmlgDqFh496tFaGG+Z/mrkU9+NS0g7zLYAOoPKen3248ezzAbV9c7eSZNI4KD
aeQwctR2hNtxb3nJB8Pk8j8QDf3q2OCztVmvvcxnqO4xfwkJq6P+uLJpU4gceIZuK6XSu2hABUAe
541L98c1HoltWM1ID3NBoBV6SKScArdpTfUu4xPOr5/WrSrrYrhUdRI3Ov4zMhLNL9NZk3UQKkXi
fwn9p6DQzKXWWBZ8tUwu41DFYNJb08d3gnb0fVyf8YeoT9lZDU57BsteFqgxz+5AlQ+YAvODYKZN
ljsApLYfjFc8z5U481vz6nyYznM6JTOhFpJuqHqqrKygi5/Wk1E18vwy61yCNpTiceTa3CHul2bl
KlyROrCNZZcNqJKiRnxvh7On68/jzETe3FVllW1qcgU+UurX1R7YiPeMFTUBoUYjVQJMbueUPcOP
bfi972IoI9gRyT2HIYBUSPSPr3cBysQB0mfZP0sfEzJ7Xaj5A9Y3RZgG2J8lmVoEV8HAB9Jqug+u
/vehR3hEsNg3V2nteeK5WSfYkBCnaWiNm2hZ3q8AsLUUsSb6oy1kIoQ8aN/6xkh7ENvIMJO3yMT0
+nI7VVV7xecHCR29yPT9SSrHIuuil4P8uSiIPmBr2g6VrMbcsCYc62XomOmeJ0E+gJ7//gKIBY1D
MrqsuKTZGniO/W8GyCrtXj+pM/BFVQ2RYHXqQtYV2TOghjSTc7HH3wc4MRvS/RrUAjvBw7OR6Ygn
n7DJWCkLwRMMPOUUgYgsif8Zze1+zxaYQjLtpIn6H7wLRuIn/uWxMvP5RoSE+QmCymglBNI3r7uv
Wci8dmmtszoBRQBz50SzTwtVzmznyXBpUxb7b2UiERBadYQaTiwC2LB+HKgl6zvhCFHPGf0y/aSX
aLWU0nxS25+/+IdvWOh9TVgY5hhuHKGhzQwCHGVExUWgf+iVjKwfZUfiV6sFVAZ0TFmH8X2NjWBJ
xv4qhwTRUTLpo+bDN4lr5HeTto2zNaOtaezSrFjGEedNzu7pf9h6VlPvBXY+dNNtH+cB7vA34IQp
gZ3he+0UG/SUMoR1sd5WB+3lhTozrpR78gDrHUVwv7iY8w/34e5ICjmoI4LqXzxOgIxASdWKjnX4
0IBAmzVz/sTweJVrArvUDNYMwt5OIjUt0ErqhSg0BhhCeFqtAm10IqKectY5DD+8fITPpSo268N7
sf0h+I2z9HH/By2zEp1sx/xN/8syHArBeJ9W7XM/a3KHy6tCBErsou9/1cNboFXjQ8OLBcUrUpDK
RrjcO8B67Sor9o58paks77DhE0XyL6ahKLEOE/EoOxj222KWBbxIIm99dwMmIoCl3OdSyygU7iV+
lU3ycFTSq2nhcnwMKs4fXED0QaRXVd2hBwpz2AVdPzmE2jHjLBHSaYoiG65tSExyfbPouCw16oVD
fZ3bYcAsFMMxtY/fVpIh/nFy+kw8AQi603Y5Wr7y/Hg5Y7IPiI3ToHxrfum7UfWH2r9pYsAtNYBq
QC1SORLKcQYh/2EsbD8LU2fDzZ7yYLn23vlXBrJDvTDDR4vuMiIDcLMCoruoCGSbFB/ldq7lxxxS
WFN+xY4nH9LHcZjWaUq9jWGcRR6C+hr36/8H6+UJ8LFOtFHt4/JLK6V2lpQKGxytxrwZjKM+b2tg
uaVow3wFAjdBKWuYnLZPHQwPPVKTSGUTAAbwovxtOCBuvC+hJrvxE0Dj+B4FL12eQ47D4q7TSsIQ
lhAqq7W7W5P3mVI9nf7D+4DEL2osdsh6FwZ6LkLR7i3F68MrAdQdTJLMHuU40f2m+fLWwuz+sCwM
hAtFneb5l5z931QZiLmdcyZjPgOiS/LbnrmomTRhStrMGNWYz0mhSiQ25KfQC6uTisvbhFRimh/H
0Drai5I/oTbjXCRgJb2Rv/myjIXj6gdDwx35MInih0WRDTpSLT562gZMhnV2cmmjniD8cSFaM1XH
Hi1D5hYPptrZsRBBsVop/Yj6PY9tK9/s7vB1uSvsfj993Hp7y3JOlNkkDIO24Q5DrdDYV3pwZFOg
3Dv4scVIygdtN+W1cvHBStPsJ5MRZHGmHb/vfsYeXin95gAukk2EdXFGx5hpn2gvO6VZA67aRd0+
L153/kTXi9FLpMWNidR3iCazN16bOG7leDMRaRiASIQ/ZBKXIz8Mlukti6ZlaeEAbl3AZWm7tEjL
MKOgGAqtKtUd8hTzYdN6D2iwnxmLlbabUD0NtRv/MBsKsUVlZYCgTYAeYOlVnCQS8SF7Y6PCrNnW
AExkZZkYdbtJW5ee0/MhB2bna6SSiVQanwKknrWyPibWDOCbB4XEynCNEKN2oGmtEFDYvvE4uDVp
kKG5aLMtyGjgyEhSuIDCBsU0dtf2CDBIZqlsjnRMHMnjheu87FUw4oK9PEoSfLJcSjwTKrchSJ/t
FG20E16MmBCkf+2NEKbBmOEmz/i1CVUVcRhksUu+Z3khkh/2B1tfTffM2EkBuZujBcer/6qpVLHJ
Z10gQ6c7f/XnGIvAGJjSubaC2EM0IA30PBMiM5P0ATYyod3Tx2yyjGZgmJP8DW5y/Q6rHUYTSbQM
QkVWcaxyfnSQ4pwViZsSkm7pUlFDDZDC441rVYmnvwcA+Mt5lPRwqTOUtq5G9ZyHO/sUNpwbeJxq
q0GkjL59bhxWY9mOT9x1Z9W0HJzO4qTJOdzyAa+i+Eq7Qpu2LAsBEweM+KrE7LNgVq/BJGzPMQeX
qdhNhKB96ElYyTBmzrEDbyLOqye4redxw81w2Ls1l5ruwc8IUlzvV+KVwpawm+RwqhTOBo0sWBXJ
FZOX4sasqzQ/NJ1CsSl9RGbrlCDzGl+ZPRytNytCnsHhiJrAcfqbp6EKvGYhZHvClsKKvL+p3whr
eVD78RUKtI7kQ1WD1kmhoqNxXKSpPP33383fVo0KXI2qvtbq8I70lqY5wOrMAWq+YWm+C5Q19Ju4
hd6ZuP/YcnUYsJjTciKZ2TiX+etY5G25fm+tFPJOs9wiclXWhIHcT57YBtWNks+en9DbVaiVCSiv
cKP8tgs1t93RT1fTBD2UxMrAy9/c1D/sFa1fRO5mmRlx0khiQqivl3UZl4y4fFkwuukRdDRUuKI7
MYOWVUM5JGIC5Z057ATubLz0WwHqJpXfgtECYFWKx6cAQvR+jR0zJsepuQiK33uP5Hu/l4FM9xWl
g3vuCyO6ZaK50o7epopO/UszCJiOL03LICYSd1KBSx1Pmq/ARlvBKxaaN5pA7ScBbbwuLpmAxjcj
qsj/YsV8wZAYaIjDgUJ9QV/HnoXbGoTmzAlzWSp15xg3qt3QHH46W8whyJ+CFrqf7Mhja0pbqjDT
O/7sy33kjYCzxXk8J4bhjSCAzfXOWtF3XYZxPhO7r6eM75mZxApr89KJAlv241FpaI60qO+UAV0P
Xlj5SKdVetUgjpVn7udOYwm7mgItW1y0rfONoDWNs0ixZ99eS9odR+JCxFpwHoIHuz3WBFyo1GmI
Q3M+7iSJkaWENV9+NUjlY8EeCHWstChf4yNwzs0cgDvpiuu/VKR13fWmmniclSSoqI5d7K50BXFc
wkGpqi03NTC6dhwR1yW3HUO/Z+UC5oUv6JO2KiF6FyTVf4p3NG+/WinUhr5OfK8W7B5NtNEz4gAK
hAynIHHdapz+twePZ2u9mlDcKo6wbGbbxqw00ZYpFJLqTdUKuFRSj1mkyhv2mJQtXLmOcyr8MDUO
XA9Xd37OVzYcVfYwefqal8fs99UOq+pKoaEzohKjVjXbcV8Yl6wGhJEyjmkNFzUOrSLwyYnncf2M
dwdTRy0iTB6RMcAoSGSUDX2bBdVqbRT1nfGePE6oGDb1V585vr3h0emSPDXUGQ+ZttDFZ3aD+cUs
RXwRFTdpm38EMHMW9xs9KMoq/DTWZhuJxN12YSiJi/ZGdejGtEVEYjbW2biXLYtSysKO1tWriePC
Zxoa6xWOxGnoZNbDEaTl7tgjztbEIeqxhZJC29/mjcrOC33nuV8PkrQj3QnsXCgmYfI/JQwDtZko
abPnyRfqtPUn8+d9ycodz0d79m8xykx4ID2zNBF6AdTQdnIdGmBVGhj+EoHeL0QKSuBq0BYMoYgs
9HjsOrEvZmXxB5fsLNvClt7jvdJdb5VB8Xp5psT7oDWPKVZumDiDuaiI8rxWwto60rz2EurHH6LD
l+hqhhW5Wl3RObhNgJQjpIhLm7l9LS8SAshWktopaQtyqnz1Pr2O0z7ja0Y1tZtHImnrZ1b5RRaE
WnfIaEk3yUIoU2y3zFLuMaFfDkWeMmr6tnQd5ATvTQKLisT/cseioFNp7bpQ13YnRwMRs+59t/91
sjn393/kKaLEh1yynOU5rqJo81rJUhJPwHDLYMwMNktzwx48JOMXni5AjbQXL9UkQs6Pppy6+iTg
vRs3RO82bFJN+BPbaK2V38ElOVI+TrQAgj69Zz1S7V16D78ec3ZqKKJt0BkE0R4BU8GUjbhLF8pi
DFITAUHchgXcUAwCMn8qB1iNVTYmi3NaB1SyBlAWt7+DJGlEx5rG4qmlsjYMojliyoa152ssJPAM
O3MXolYQDhJICJdQ8dAmkq3ASIWWhMatiHSTJwvaxzGWN01FRyFePHwDfnmWJ56iMpxiMbe2RLoX
EkfoEdszF7elT0j9HXDD+amsWm/YdhaR0qmCwpEEcY6OlbDJlZ5ly9x5gFQ1Wo286C1tcAyhAgQq
jdJVG6C0yo5zzYxEfhYY0QXVpP0fk/ATfGA5UizTylgzteaTdQEkG5ChvM0JlUphL3hpGwOcw2Bo
gF477/7e0A2rI/IcafEnaesHY/cIfKH1Xx2xNFFmU/q7jWLFFJK/bcens3zFPX0NoPDAk/vEHlSd
GQUahX5FWRvAttJb7d1vW57QI3P4ujknBzlMDoKptRI1BeCSE0oYvA9utE18XeOYh411cPuXP/pd
JrcoxIyZTM9iuZht5w3Syj0wu1+xHdxJJIg5bQeQf6e/2QjX0SmB3NIY13o67LImsYq7Rhh6YXSx
HroAZbgDIQreO7Tk29z4sca/TePjOqAoTDCf4HIuX78K+DkeCb1ebXZmZ3YGWBwNBShcoyDSLxD9
G9BXuGRBk5P/A9Uu9CkyeGsymGhSYb/qUIqkgj8Pd+Go0JAcqkciJUuMj+/zDWlxEND71LzfetCj
leTdfuHC1r1QTc223lvGNTRuv6A0Tn8y5fhSTh4c1Mt+GPBMT8AA2OGUR1hVYS7UL5WhxaHPh3ry
I04pSbKw8Py+LOesolHZBGfYrM9XM6PG5mUXT1LmhV7IyxTj6nPxkfDZpnPYaUhqxuj0bV7zK9JE
670ptN5wBLjpYGfp8hJ7h8sD4QB1XOr8elGepce0fDB7WxUlp28RttAhLdbzO/bpPLDQ2N3S9zU9
GzChrk018/mNWOe2vFJY7ktiyc68Umuq0EzpCZd/FHPI4iy/CDi8rx5+gqi7NJEJ1X2DbIszoNLq
CCrKVtvVOiImVGiWaSksImYuLCRQS25HUmVS+rB0f/i57dVQeYKUhOJTKVPJOnMaZ6kucDAkiNlW
Y6DHBoMmfzfQYZLIoOstrUJh6Pup+ZwOths7P/BK0sJKLzNMqwKcBTZBsOImBEqy0fkdHqUoFP3a
IGYQmVmlJ4RuN/LHPdq2wp9SIaaKmsyiU6zs7O6WwpokgcJI5z8Q99Vv09bLiLoCGALTzzfKbVj7
VYH074e9XBvzBeun92qTG12Tb9cZu9z6yJL9TJx1lgVpgWYsAgy9UzamoQ9M7ww6CAcyCSqqUWyV
ykhck7hBwptsSIXS0d0mkeP3q85GaeL2WaZ5GzUtXo/rWUxQLd+Ml3Osspx0IKw/lvFJyVtLgl6S
pLzaxhJ8ZK5KV4jFGVyeWyZPqFC/Xhe0SMbQuRjrzwROQThR5LeJCH6AwhQIQ+EZCY8Wgzfrc+mX
TtyIe30ByhHO8nZBYcPMRt1z35/wL/5rIekuDCe0hoSWacA6H0VoQthD+5wE6tIkFZf5XjQ/TrqE
i4d1bbuSlnZ7gtcjhIXlkgGQz2UliJVAAtrsJmFulBNRaVLng3shHYWVemP3ObneUX2geoofwHVS
9qafOZdYqCoMlziooBJHdsk6dFszllPFZwlnUudo9Zm4tl0uP6BkTCxVd0P7qdveSVCi+26mq0zM
YySOCaLDT3HxQdjjtdmgZvh8Meofqd/ATyiY2VDxmM5azyL7MypzDRmTTQg3PVNzHWErnZuaNSap
DglFm4TM4crP1PQDLy8wmjLao313C0mL4eSa4dvuKEpyCgNWCjv/iLLoQqA7YNAeEkGroTbd2bd0
jHC86Q0TSLkEyqWX6laXJJ9inOUQAoZyqH0y14ZCMXezMVnuJI7s9z55b90RqXZ2AXFSH1P3ccdX
0oUb2NZevkcB4ptrSBmMwOzRlFUhcvZhrM4GK0th8YM8qAhzbX5UV7CRdnViq8KGvVOCG9UJyKAO
1nSkiHaCWam35SDJJV6GIhGZrJie35zC6h+wdT/ORmqQAbB5oDZSzU7y3j+E7rsbnk4y7I/dIXT5
byKUR705d+sH/5CsBTujMcgU8wK2BrDV0jbdFaQq+60cKR27ny0XSOcPSk/qN07HK4vWku1Gesqg
rY+VRZJq/BUMvRaeI2f00ofEfzPMHwS6kz9ddpwZvMBD9XBOIjHLgIHQNYydwQOr1pIFG3IJrE4A
MIKKQ86yfp3gUhjofEwx469mdfUwVvtvB3gaPGcPIfWhiFLhZrPZ1XsgW7Wj4HjoQUwn2l6nxZ22
PSacIGpVUTdFP9bnWU16SqtUlNJvE2BohfYLx0M/2rqjahctS9RFBBGIHTmVYaSIXrtfmCUQOJf1
mN49VCUqRGZCtu+GFS0Y5WqZ3fmbxiOZNI4QwACezi3SzNeIjs/7VbQDN6Qf8J7/8s4N0y6NXPRW
V3B//aUTr1miW7zh0jMbCbT45XBwmBtagwHwb/bQYqYjKsYMXxlVv/xbmnhZSJDKnNRUKpridFSy
NtRizJSyZ2u1hN1KmuKbc713b6ul61zLFNPfahpok6T2Up4N0wT3Vw6gAmLGozBoodabc6h48uYs
MX3Kr87B7LmDH2cB/X0wMntxRyxqpb984tGQg3Ic81dvUPyFM4bUN7/AJy46inDAEwZ2A/Im4i5i
eTj/R3Lq9Lt+7+x9l5B+EMuVUD+TEczEqKdYAMQpsV5rho8VG+q9FUZojzaSwNrratiwezt2vEW4
3o5/qbPmwb6GzUMYEjG32f5318qb/Bww+NkX0Y4jFgCdg5TapqSMrh4hMqMjwV/MBJY3ZHqQOeeh
j/1MsYScMvvWQoUtdGLA8xH27XmXK1+4e88hT0Y0nl/5acls/gifXz7fuBKO2nlT1heA0L4E8cYy
DP3V1/TgP42d4dIpbF9ArKzTtPiAvauWnQY9TQJechFh33ESEPOd20nnxkELFNEpBsuKao5gA49R
Hkeo/RnKj9s/pbO+r0odhNtg6enqrb3CKZhAUDm/uFu/JkgIOPZ8XnvLYfe5jtBkHYPaVygcbbkc
BJbvpIzTz4s4s7sLSMK9hEziGhCLcISWNkPksn5sZzBaVEAgs/L8dEjkW1FrCR0k8XmhnwYedKP+
L1GDdSy8gPEQIpgs6IUvOEqJPMupEFZEc00Qt1pVCxLTfcb3W24MjvgKtTtfcGa8QL8Bui+rdOBU
yWS/q35hO3FYFZZYJMAeaI5ytp0Cxv/esLftwvn6dvKCl+STUOV2dagqOERnJl1/AliqxQglZgLh
/3WEnTYygMf5xT0MGzlOW2VMPP92E3F0RlxeQ5F/RBXdMgcKIkJJlQWdFJNF3GHdUm0OOHBh/7G9
pSy3qcUj5PpdC9E22ZTGEtzb3uuaN+VphBjWf9zEt1uiCovZIxF2AC6ToXKIZhcuT4rp5rqpewf7
AbKhlp59ZAz63DeQ6GRYMwFlc9/hHSIHl6rujjyTrq3tGq5vnJuXL6FELHARhmSfc38aKsYe6cRw
XVF23Ciu/11xdvLni3t/mXcBDhXdZKj3OuPdglM6olPQixAjxi8HZPx0dlj30yRgG5J3MYujlmgq
DB5rSHB2VogHxLUmnhNaXPYdP8m27NXOvfL9Dni0Ejx+F+DPApmJW9IMqiyp6HjYjaFrnMtk0Fln
2Gw7KKCdISlTP8sWCuM9Nx42t5sncuCkWZUKNPMPulJpsf1Z3WvtLKAtVFvYuWx817/iuk+lO5Fz
EoEAB4NCJoEio2msxdRCYHfs8ovFf4+HVJ9EZzKcD5c4ZFyp74RIG/HJV8qeNEDcDtrBq/BhwiET
RWLF7/NkrBr6igndWQze57H+rY6Y+gH9DLvvX3NFwuQKgRM+02gJ8v9TYdKdy3mCkwhUYOYErjnZ
Hj9+XT89KeQ+XW3Lp1yxl142ABDt9O7FvCQUc9dZLcMuHVF4UndM+Gd2F5B7Y+eV3QYbFdCVlM1D
OwhgR7+/z8bNxp7IfjHg/9h2JHa3KBvWokaw/wvIY79NiKhaIdgwxJEIQC7jJt4NVVZHa+Yv73ak
qzLl7ax4suRinPJSkEJ1LEvOVHGDyCzwCk8YyKSvZ1yJt8dWH2QwVc8760hXcm2xwHDRW6dsh1LA
OpdNAETgX52+3KNFsJ3ANrGgAjrcvkWksJS2kbxHrgWhNp1TXfWHcfHRhJFm3kEK0qwNSFZNLA5+
Pq7xXO0MCLmG9rCNtLQEYNLFxttu3WDXbQddxMmPV3nzDS9TwFwqS9ugLzAShkxMO9Sfold1jAgL
tKYFaJdNdQjFgfX064GlULkYAACVRXeOnFh+EDiiLEuQPBgfXkSuWywoI4DDcdH7DHvYwXzw5CPo
Ae90yp3/U/GKeaoo1+vB9UHlbX2vhHjt9PATlhfMjKhism6czpvQAZ83HQaSQZnqJoQY2p2nlMDh
8Z60tcgLxr6kpQr8v8s++KZV0yUbx7eIajUgz5l+MXC5uInxlp+/MCx7f4aM894IQeG/ZXR+N8nk
yrRhvv93U+6uFqjhy8+5zgWkYB7Y3FJ4T1wm9Nl7L2Oknq5oQnROy+hemRfls/qKG6xRG1MTAEyU
wRhXf+Qbtyc6T+o2pj7bCZlUjqtgaAEaTBAmLZDYTwKh6jpB86dIrbfdcvwwtg1wH0gviPE2/Fbr
ORH8HrJ9cf5qhNMDHr83l4cP8ZgKNTRG2tHZZZCusyZCip9KwyyMsRxWk1qnh+vjTYeUwTE2DjIa
Yw54u3dvU7d+tygIBpxhDOteKemRSJfwtWzSCdr8g3ko0n+vv689xspqmeZLiB624P8GFOMgSn1j
qtBRyM7gM/X4ikef5+/rl4baSlfYhpIys4tWgSInaR0KSEOsDcbZ8TwhWYKa+3WM/WXCEvbdv+br
2xQ5ZjkBViZv6w+WGwAM50PyMTwSP8/oej8MRKM1Tku0L5f6x3mIdur222X3PjX7ikjGVC77Q7A0
vgSBR6YuS2UCJlyMhoEoibAVMXtT97krP2aAnHObGw13ASnw7v3TyQXUjiUTBGY8zAFd4ngWaNHL
n1j9L35OJxDDT5p73QPvgUmXMjmKjgzmOd0HASAukYaXyiwNG71Ypg0mpYls2bnzge2/qLXiYuTP
UeZKTe3lJb0jJo/fReLuNoBPRqCJxdqQf8F85aM+3PKy/UWNjKAB7OMi8Canw/fx0/CmL+Pu+q4L
Eo/cp0grlsS9OPJpez7QAKJId6QpblPj0+g7QWvITu+N1IKK23QjpKhv2EUH0Q+IrBAv+7d5isue
cJCkNMoCURWP62ePe41QzAB70TjozJ6/3/hZ/DcEFR5wQvCEHU8kLd2a/lq86YAi15UbHO1ZwSg5
KPM4ceCPo2gsThr8mWXZHX5n/+Lqy21QswP4R88rDoqdXiIaSav7e8JQu6y3tS3t6quztTv+Hc6P
HS4CS9FkZWCJjfOW+EeWxVaHHcwTsquKwYfuZJ0I7ujxNI6et0OR06b/G58cvW18Mazagk2O4epm
WMzNTv7hcJ/4qYrSHAJwH2sNEtWvzdEfzK6uMl2rRHVjnUOJ/ryO9Kurqb3CB7pd6onrodl6znft
R2u68kVbl6cd9pCRPXl7wQ8MWVWyTFxCLQunG8AAQ4kMtmAON/BoT/+nuDLJnmjGY82reCRkjGEh
8kdPeP9a02BaEYrRxbltya6bIBlTYPEsrA0Kajm1LjMlKqrRRMVTHaWmfcqxpe5+1VMAZU/jVpJA
ZpP7eJrLKfWPAhn3olJgHiFUrFbwZH7uEAQe8wP4mXp8yEn2Ue7t5rIEq/2dvdMsVGXeq/cWWgCu
NNFv1D9TfeQgUSb2UCyy4YoBTwnE9NMDkX02oPpqOkoZoZtkryehdEKiEUXJ+hNpuwO3Jx0fKCRc
r+cm1M53/FbxtB3HeLIFeEpqf9458yh1KoyAjysefd9AqPUEaSv0kWX/ZJUhKD5SIvsPbsz/mY0H
AoaiJgSzIXwf2wEzBpCsVtn2SSflSOqGcXF5PjdemyCrzTv1E5lhJH1ivvS3bCYpnM4HWhsIVlwI
t5bHZgE3iQ1Db4l/sYSgDDsaY+ALFOKIGoVpON7CmSmhUSKLjG2X3OttDx0+KiXB2wtwtc9TRBu9
VgDAcyd/CeVN1sFQ4LIwEdAtZjdLMUszofTiIJQe1GCEu9LH51JF+t3WmpqPrwZd2Bx9+KbBjp6O
C9NiWpC116oVlvOhrfE17F5cjZMFM24dbht8AE4N4ChAQgkqs3DhIpHxbslWW5Se61FLDKh4iPcg
BBTxnXUx2Y0hlXOFEqBHXWY3QZTGbmkVs+7TBgRu2bEz+0jVg2lzkfiNHXbjrvS1HT72TKJgTVPe
DA+pKW7890sJ2aCObdB7Yd9MmeTno0o4h1uGeXd65+gHI4asw/4nbxfFRL/cMb+XQzC0CTSSEffY
x7zri6TUt4L/hwNPhikczt4OllLlsyScoY0eM/A8PxOusqL1wx0VJC6BM2z4S0q021MnSBuLrQ+x
BzF8s3d7iiRU5KVDhRXQAR8bz2XiG0gx1UQG53vUr3InkKhEmcoBSPPg3jlk1S4O5pM86Osd4EYg
OGv7BngZ/5BjRd0YzPJg3mkYRZEjoNWVUMLEiAq9Z3p6iJqu5tBBz36ZkyeA/x8mzVG5tUMba/bq
TnE4FBFt9LxTSyVoQAUMVg6IgEIFnOjiqfmMfGIOI80Oe/r+5hr6DLos5ZbGkCavN+54lqMGp4Qr
a94JHNUYjr97gn3EAtQSB43AkYlaBcDWHncExfeTpNy1ZDyuMdLUDIQMsNyf4KUIo3sues0P1a5j
es4hfdvH/fa+2ddu0Z2bSCGe/pF9tNSpQP4TiJlBO5e/K9tEudkK7pJW3b9l1PHSBWIoTp8tSWHD
Rm/bi9w2eXod1DLLo1yq01m8fkWlyFuyeHcJcDIy6GTuZcwhE1WeuUO8Pd7VYD0mtO6ZhVf0HElS
XVH3G7/oWKxiV6Kz3wBS4huNCL0W0vLpXHxX7xgvBa8uidNsBA8WcDvw0Ffsk0acdDFxcrCu831x
mE/cMymz4NH1kRqLvSDEqvW1ds0iY8wkvMcn83G5ekYxQ4wBu2w/VkaPYDwY8g747uydAv2IgSY+
oWr/yx0U9tNnKfZvLXogK+1LIZnYYhYzZ+ljItIFsQnoczaQzbG6nMrrTIQum3MH5bSgNk2m5boP
vyYGhjMDMRaUFEWJRp4yW4QZwZTQAQqHRKQ+km0pB2opnIBgdtdUl1PoS2aYgqcO9XYvzM5pm1Je
bgpzhUhOLz8d5GyVztX1uYGTwAeClu9mQfbSuH9XFKFZ7R16h53nnaeXu7J2hl6MWp2GBWIpE1vP
FEZaZIA2/JP4iIfiGseCK+69e88AR0BEFgBenejDqsJiNyvyP+ZUHCb5S1i5ha7AxsBpwbGloUsw
Oag4q2q/cjMjVO+Mf+3Cxb25XLzC693hzc6UF4nrbVNc8KPw4Nr6W/DbOJLXUJyy0PLRi8TBZxmi
xhTk881NUfcqKuvP1EbkRrgqkdilc2xZ0F9mr+CVvBVIAchEaiE+UkxRLQxb/oM3xUrLD1gd/nHj
6lJ6rQsOnsrq3q1RGcww4g95nRlIN4nBVKKdlsbvpjJv89o6/pH2MELaBatAuDERWOGqqXVw2+ZF
USOSImnSkV5xdOu0DwlIIIRcDd0zwE3GJVMfqYXmiGyDGUJXf6Tl4xAvY4MvRioPHrYa/FR3nrHs
qo613UjbV04SXSloxbvp2EDnNxrJrHd1DXv7kLIcjaacND4NCtR6ZZ95bajZ2F7GP7+G0FuNMM8R
o+39k7MRQpkMjzVmqCVQd4EqhOWALxBP4kMLMAvpFc11VeA+3QBnAn/n7Rl05zwnTDG4oBxVhcmu
2f/Qzg8uCl91ag8hgLV6+Y8vdFIDVDYz6JSW4+NQVX+vf/6abyUafUE/wen6FtnXSPs6k/9tuMgZ
ThzZMhE8EM0aUxVPnaMng8chFOev2a7M9DjnLk2tQET9ASyLl3LOz+hMSUylyCdEEA2YXqKSajD4
pGhVBwaQ9GkB8foafY0UdYo9MxHARX3oC/boQ5s/YTy24gzXwcIQF5P+5rSj0uoTrTj7behmExak
a+2F+siXus8Aq8qqaUZa5RMZHdTlNNj6n45SaP7twFlO1qmaUiXAdmltQu2u2VJDTMiwTwtDgM96
Eho7N8YIc9WkdcmpYMdKnj96rJ/1aCnothMwfV9OAfpgolWmyprTfMx5OgEb1QqIwfLyeNkBZVCn
+uXWTbz3HuQC2K5GErxVwJeRMe68SxQ35SXHvhHFto/rT9hw1+4aBsRR6qAKPfQUFsWWZpxmNvDM
QW1HbObusgujhH9vEntIzxJsiO+WdIgoZ4nNm+vHVNw+WzJs9HXW9FwB0CKNHGMa7Ek38zvVADSd
vRJoq+41zn4QVNT7/flYuMO2QR+/6mXZ7xtuPy4SA4jW7s6ITeX5zRlDV71UsJUn+Sma77me2qRl
/BKFMRTwokFJdS+vjUHtMKDWAi12mz9RZ6MncZ1Wc+sM4gGwVoxOHxvqY0RTjwPb+9EWzbEuAN7f
2imO3tlWbq/41EmXEnrszcp63dcMsX+8PlIHiQwMp2V8F+Xw4Bej2kbuqnXL1f5exHH4CTKGfT5b
ky25BvlD4IIHuc6Uy4sMYxwOGMdcJOpr/ZX4xVuMRefSfutMuZZW9+XXdmK2HbrRtWY+AbKXRQyq
/kiiYNEOFYYF0pgNMlikfFhVIs9B8cHITrMcuzZwmaD1v6nO8Q14slxIvcw57H30qcfje2GH2Pqg
sHAQPCzWgtxYRCMK5GZk9q3CGyOC1nxa3Vuqn4yNSYtx0jx2Li6jqHRxNhImABNyXPehYqnsLXiL
ojLy56xaGBLmFMQ/bJggWP45J/cFybof/t9uh/0OQ64elGthDKLabqkVaO+KIEximPgLHD8XdL3/
B84EggkRqTTGa524BpWMbt7Bx/n3Sr/O61clAJIdqTxvlLGdSKHlE2OcU1Nl1zJ6VlYOe1ShkXDF
EYoEbw34l0JFiACawEWzsZ7IGmZrPfg6zTPhiQ0atGzhzV1fJRpI2dFK4k3DWxG7UZ3BHNcnL0Ww
N0D/4e5W9KLYkqzIFB5SbIp93L+PLAeTaHN92E4hxjrTjrbnysc1vsdlyQ91NrFZMWd/E4voLASM
CHaa6lBcOWqZdF7eXrhuw3VipQ5v/hw5iZwe6qtAfEYq44GYTgd57cAg2pqAfz9/VFs10lwjoJSU
PmlopwNIvX9GNPjVBKEqZ9bN/clOTufrPQrq6f4i4G7oNY7dTfspgpfYHK6CO0CS9VZ/eMcROZok
bHK8W7x0O2IjKA3B1J1w5vchjjtywWO99AjyOEA+HxevMrp6e4jcG1XFH1ZqebU2/Eso+Z7u0Dn9
cHThogqekvhWKnR+CH0Hw0GKqE6PKG967mFBTrg5uJJ8oBqYtEzUHnNJlLC5UbKDaaRdEMHB2meV
dfqQedgnYl/Kq+ticVN/D/CojNd+ZtwkRxu2vXTLaVe7EqHmuA1fQXAiQsp076yN7k/Ssl6naNp+
f9w1Q3SBUf2QjcD1qFssR6oP7ikAERRcPiVaf99BC0UIZTU6SjOFyodrq5Mxzm4VaQUEvIe5b3F9
0dyKZhf8FV9yWYjhxGhLwuDVgBysIARccGI1F5qf8lscccX1gCTOE3lNjTeQ3Uy5mVpFSNTdibZy
HDZ6wARNM2+OmKH0iiY6G7lhEn+mkrv5tmt3eM+XCwodkDNGLRY9k4HYN9reztJ1Ciyfi4hcUu8+
EWpQ3ARagIj/T2KztqT84YrdvQLvfWqKn4coFDkX2pIzJmuZEOFW9CzK/M9rxMZFyAUiiX80bzFP
RkVUp2dYqlYE1ERsMWe2jpwXyvfLp+IvoUL2AXWqJPYg+rKuMJVLKZWa0gv2WbIQna5AMILF5TKn
2qkqVfmgZfnzvC6fYPods0j2oz9JODwZ5eAXule6H4tXWhXTiJHq4wkYACFdLTk4LreglYtmE1ZF
2Y6ah2QuovALpWUF2XdZTy0sWdpdZjRSB2XcyabFl22Ozt2Epeapf64Vw5KqOvt/vZ3vhP11iC9Q
tIjvYkHNjoAN7LOXCYWixhd8Ksdzh0RLzLmhZAWGFJ98FyQqiodFMV2WJ2YOxLz3dPsWTOWzVrWy
SJ2l6OIlk1djPxV51o5djH5vQsYT2CvMf6hTsNpyZCLkdMQu5LTWfZNzu0o8RF0iTgdWkgRgbGy5
IH23Y7miiYMlgaORp+zAQ2JyHo/bQvTPGAwV2Q3pReOF6gX1zOIYCVbmONWCC2hZGxaZdO5PwnQs
s57AzOHqqWjt0RrW+JsLX+r+fAEmXZoCjyVbNu2SA1kwdjJBH3arqqSj9vNeob3a9W2o8vBDpxhg
f49xgWhc/FR/vYUtQdprDErsCR2Ori+KdRjOM7+n0G+vDRW6V5++MrLezknDqgjyi90X/heMwnw5
OjubJ+hWZvSq1H2j1rwo1xSirbJdHJ00AxW99FZGNWLWDa+DRrP9ztzMohKJI2Rvc9Mq+oK5MDhP
j9keXN4Sq16IRZk1V/QSvd4s7jo2ZoOShFElm6bTkiC0Y/UYI/PS4YN0LKJkfMZmgo9wEQ1UqIzt
EGxekEXJElmhuZz6A3PsFo8KkKr1Xstp02b6f2m30W4cpPlk+Pju3N5nnqUAxmunDwTCjWS4axI4
K4p3VN+xDL3Qdj/QqXvPBbK2Yb4nO37+EePj5cDMrYzl00sl+8UkaURygnrE8irqbUys8wqvCfiT
K0w6NQYQPjmjES2+ia0uC9OzGhlJK6Qs+Aj2+urbpCPtGSiEXmMaieEHzPnI9DqBjA6BQ5M8vM5Z
7pIMlhC2pCyPQ+zYbsd8MItUCdG0zwZW9VDHKodrCF1rG6EemvAFw49g7PYkXTPtkcHKjur12giW
bJcCCJqwfEWVmKDE9qIR6r0R53ElDnPNXZ0kcG++O6zNb9nb9CrGuxKBryVYii/tQSLEHFVM2JUg
nk0uQz4GUfwA3srLoOfwujvRRRowrocrw2s2Idk4vYTvStXU5ZCNZ9zRlFuXg5Cx0FyDi/XniadT
fw6wTDZcMKu0pixj3Bj3EzejJS3RN2ZGa2v8RCthtlWpJz8R4vhoEjrdmKBU9DSZfUlwXPqsTK2o
Ddkmmuk92UZpk5lSB2yL7L0KbPL4rjmj6dJumskk5Jd0hO/4SDWBXBpyLU3abWgHJs4GRCcu7W8A
SOF5Oi15huDrWxzmHCQ7evb89Nt5iJSU4v9Oqk3lplMkR9YhezQ9Cv/pgVoCBlqzPY8PHfpBIQTO
XNrLX2RyJKoJY9pNTH8Is70pACXi2F4pv19T2KuEZ4Tmc7VRVI0RFkGwl7xxwjsl+lFKO23rVWOe
e+eZ5qDesGY+ZHxRRs9WlzyI+XQtakNE0JEEQcx3CMEzQxZDf7MptRfIRDXwbNvnLMPrabpnmgCw
5P6JHhZ57x9Y1dnQCLx42v/lAbu3qZYa2fClNll0wcLpexTTYc9GoQxRFvDD3p8B+E7chzARR6lg
ZdBEz9L+AE1/AnSzZUtoBQ6p5FaWgD1zr6PxU1WNrrf1GTOeWUYzwDo+17pezsFsUSBqeNVzHxHg
payBPC1Cex8zvpvKPRR71FOmQ+hVw4nMP4ttOqPyeskp0BOLE8xdb6/xYaGpPSvZxAjkQBIrkG5z
EBWgE38pH9OLhLCbypWQv5+IHa6FPYhdKT8XToLtrVpjoAk1ZInylsf7Z7NOMkC9UZSnqMLj/1RB
VaN5Dwl2BeFXT0Md04dAvHP9+O7YlAKg+WXRxq9bvqrUfwKWbQuawf7BDGaIYt+IJ+fWYuA/Akx0
sPeeWy/jI4PBIgl4k0JAEzmj8GN03dzXUPvD/x8CvRjrUTsXnAfL62KJ617TvzlaHAlq7Dyr9gvS
/KL+AQgLwi8tNOWSMpXaPEFKhoNLy21SRMwvWg/icNFU78OcOzkvefJ2E9TOao+m0mhAjMnPfy4B
pMjtODyVl0r1m/GyazSCupJAzLwjl6QIAF0MdudyUTiHkpuyrou1eySpbmGQncLpV1d6QpRc1PzA
2X1JO6sz2Fuk2WC426vbSn4B0vdXLq+vO8PiopWIAJF6D6zEklKKINn+SmAibj1Zv3aE95eUXyUN
GetAt9EurlUZg4fmrKYf2hRPOcL8idESYxV1k+xPNO2oqXwHZc45zXCgkuaVqE87EH28/xLBw4dV
utH/uv0cv/HqZcIphpyjWDypkbDs3IlmjKwyvjaHSbVafcSy1FXWTISL9hddam9VidIrsaapvpZ2
5Y0F4ahApDQNQDRu4Km0GkhZAj76GnTsYLInkNp97oVxyGhZUC51FqT/GXPBarFhs+v2aA9W9L6O
omh+RL7CNL744e9rKRN5fw/GjhG/yzztuVngCEeCafNZl2iG87U1/FTj1uqSEm20koF//fxsZz5I
bByGxdNjUW4Dfa27cQ5oUWj8zJL3E0S7HWZyWG9RyYBX5CGP6S5EM7XCy/8GHEfJ5uYM3l2O4qH9
0QRVpv5uVZ61Rhci1ZQNlwd/aRwOCadd6SBj0membzbAApqslTSysBBJYMDkw2Spg6jO3GkBNhzu
p0szuRn/enyagzocO2+6z58ckmoMNrFqjGzQrjLID0YIAowVji9Z2OadeQJ8/tm+i6Axw3eiFa+O
h5AqkVfX/EkSw2Hd3KESvOYWWdvcQeSVy84fWMCut6nAS6mn3EeIPO5qBax3OXW87DX1I5WQB28J
UKjE8GgiZgCqNcfLFaNz26G1BXNluK7yGMO5EpINRDjIT1vPZvwFXVHohfvLoqZmnraAh9J0+7/I
nvJyWt3Mlb3G64t6txXb9AYlxZ0w/kA1jyc8BU8Xc/1GZ/jyTfG8RRpOJiYMIeo/OQqu2I3C7zl8
T8IzlwKHFwtxxyJ1xLsSlJ1LPH3D2Rs9ROXahJIhhudCZO5rkfmq7phF2UEaZwvnQdUFWPeeZx1r
MAAgMWx3BcrxrCvH119WAXTGsPz5D6GymIE8Ub1uOo2tacuX2naaXmgnluXcEKfWYh+ZbhpcBNEP
pKINogj9lQguPZ6R7miOCNolssPkny/MK9YTpJqw37/FQeZmfnW0JsO+3bvzlDTZHLv38X4MdgP2
yKZ65tTfzzEEBz+RcnUhqH+iUwmhEIRnTY0su2QLv3Rx8D++4GMlk1k1P9RuXLPnBlilgOsni6aH
dcZBvAmO1q14YRugy2wmpJ27i7DIBkNNZoPF7R3wMwrARWq/A+GLqxLR4eo3t4e4YszxenBonxBh
5UAQM9ipGrfxjVbCh4zAmpfnTdhvW2EOCFLNKE3dxWzZ+RLR4m5+wWS7L4nm9DWUABDoOgdQy8gl
CYToYBBsk3HIHsHBHB26MrapJLEy28Rt5tzWe0TJGTlUWJrPCKe/jLlJpqHT9FBY+DgCj2cE6ZsK
zsxUgiUSHChAn+lX9wBJyn3UwaHduRKYoXLHgyT46SE1n9ul4SGAuWezaS/7mhIYm3Ci7jZC9Zc3
EH7c2ueAKCVphkyg1uvesWYQe5tV6FcSqPEqu9hFR8JeJvUmFsTQhaFRPBypwwWNtOrUjwJb7ePJ
tpK7ABTg6FutRGvGlrqEWbIZ4pdE5TwR0zC7OdVaVPm0aYgMSn+gEFCzeYNRkKRTapF4ZRGSoX03
0uuV2lGZSsTStH93RuUbuCDQxz01gquM9/w1YHTybWotJrRPhULOkkidGEFk1/C0AfUG/w5c/ogZ
/nk3CT6iQUwWeviCN5k8VJXktG1cYg/jVEgHR1NXbHeybzybhI0vzwf8r33sv32IyvXU2xAxoTZU
XIdflwlsk0gR2EROD6Z1rLbmFpb34A/pyUh0K1HfjKfkLsOHDQQWJC67mxgmVO3ukwVRQ0lNFBgT
tqdeaWbSPhWzj3X7G4xWDepnBgbSQUnqZtETWvHcKLLvK5e9uKjsYmJMefphKICXjGhI57O5oFaC
zeAzizd3SGsFrB9x6w6e8XJUvsvtVPgE/FRFTdu13dT9YSRyobgt11I6BReJoFqYHdCguHuUzHhY
G2UbhLrVvC84qNbLZXyH+hmx9ahDvBgIF30rzF39e3gcV9D0kdjrp/EA5Ptc12iadejY1p5xYtCE
Yt4mDmPOyI8898lzUT8gDQhnwOZ0bXBCaUV+IkKA4lqYn69fOhZjbEam9owyIQiHX+GKiHURl6F+
YCC+m7GcAuLKHm6vMsF/ro4tSDIw/HFIVXgUwufhj4Z8CTftXk7b3SX8weMaeeNUm73W47gmCgsv
cQjhLLBkryAJjAhJ4wSKLYcURCI2RCjmymYSgShfxhUwMiaZMF7X1OG9pbRN3xh+HXxzkJJcI5fd
87vfLmfywRUhLwXyyo2EdWT0pSM3RXi6DtFh1pHaS+994aKm2W2d6F2k0IgcxyV3HLUfHv94Q4Ym
yKgAS7Eg/w2z+t8FyPy/owGVuJJpbUBiSG8CW3IirFMu8Wop+z4/k9EFbEzJLSRXMwcDpK6VgdEk
61O7vKEEHHpwT+Y6dH+GafkXsfTc+wBtNmfwZswRtNeWY9lXBH7thfZl5x0letwU18EYG14fzo3Z
Yk7IwxVNRw7PtXqlzmw02NzJz1bd4TRlg2UIe6ZYuI3gX32E2HGUlTn0PwEkSX5QXIQoBx+J
`pragma protect end_protected
