`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175296)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCbd/xufmegFFN7ofJ3JnOOEkcYSfefK8dqqsTtJIGMD3GZQJCdB5P2Pl
odMyUPfkuN3+10lT8HI/cGY9nqWqEaXOOkvIOmhMp6LBgMnrGagy+d3JN8abu6Wv0PFg6bgqFgfH
gPwFLBN1NMlrwF+HYR9s0ue0KUcPh8p3cW9wpA1xOxGVlceMpDXcW6+5UZe4I5+/I7UGSVXyr4tc
3h1wJZrHXNFQJjFy3mioR90eRhoxO0734DNOcEcY40dRIsnavv0PMtMmfuFMUwI74pXTogPeWj9E
B5Sg12DHAHINagctpMGoWSN1hSONy+6Pv8PZtKDNho0cpAS0a5XKTGR+pV3+8JJyEIwwNC8rNhjG
z+0XfXhQM1RM8tGG+moq9BoEpi4iOSklGAhlPg/s6zd+zz62OacgkUzby3JfT99hTzbAh39q5s2h
rTNsZr/g9UdXX1sB8u40MnyC7KE4Ykv9mQUr+kZCkwSUyOoHgWzvi8NC497Gm2mNnJh4IJIs7vZw
nxvl13hqOzxUIUOUeuzTQY2nQYHaKOEYGCAtKFUdkBPRX+hIKQL07zZGzi9UgqGUaKSW7+GoRwvc
1SB7+pjV1rcd28yTlBHrahM5G1mUT9cgYIjK8VUIhrx5HOZqtNLcVIJG9uEFQJSyxvWly0DGCyoI
3essxR5P63sCHOSnH6/FiORv+1nmMc3Rhzaqst+j+TLmLU3QvQXO5ftPzJ2MvXzFTYlLW8HeHNKl
ywEqjEgtEYBjUaICZ5/thtjtWhVGTKlAOJDn2pnoczQYtJzWOoOoZ6/sU39D0sVAbN9RY2GZnI0T
bybG7SdaTckQjwQUKN04hngRL1crPUC/Pp7f2Ey+viirf0ogj6zdTZHDhhnL38G4Kb0xSFe/fXSt
RLMpufllEm1qeW5xTNTokfsBq3ixLPwEr7p29saO5Bp+U4kkBUyl5ydKA5x+SggYdKAIGvFLnhbv
vk1piT79vgG5e1IS+6G45rgmeIJvAC5V+e7T+9bpTZ4XRnhxyJ1yHOWDcIKiRuwVwk/P6fi59pkn
iDYLi9Sg3o/BpGGMdCK+7G/KQHrXyUNUrJUeYudoQNHmAz8uipHXXWPNxzpIGHyna51POhh2dZtO
oFE0bwgGyc7uJCNQMB7LC3NrnnAamCFD/JCiKmwb0oReIcB+uXiSauhJCtOV/zBZd+LfpBvi5uAR
rZ+7EV79yKQy3VR98OIfrQ21FubDPQOe87LdGsTEMRjxfxGTXCj4mTqqjCSaHbDjToOR9Tkniu7T
cIcjVq2/hb0TOJpGmZ03sN/36P8gsDvpnz6jOuX1iqWy/cwKSIyKJaJr8/Olp6k/oh1hBY2mB9ri
rq+JHuimYMbuIH+rLVA3+s7L32rCkoeLON6KhTj2SLcPv1IbuZEnloMUOHkaQ4gtBEsbbWSO3oXQ
8RLGdJBlJ2hmGUpbS1bF8YuQh79IhtsG5S2q7mxiEdRXbYoZw9gAMDJJnJll07WPKxEIrk9KLKr7
4K6hh9svjr0pLWcXmOnrYL4ZF/UVh/01LpIvdnsfNe8KXeLrnajvEgr0zEw2y6Id72glYiqs/jP7
2Il6fA38nngpYKdhRqMZ7YFlwX7V4H6WnNY7ZZMNEzcRWTrlfQ7LBW8NbYq885IYl6D9oAC3m+hE
IK2FXKep+RzjPyxnpg7uFUreY2CoDCgHbI9hXjnaLG+AXn4QQUZoqkhVt63YKRBNmrG3gFKKOGw7
Mq3wvUthYqmrxUTJRv0YZhU8+y5Y/FGSiwevYhffL42CHbVmjVE7dgchobyQ/VEjs50jRSE2Jlkc
RIBpohLLvAZ05SwhQGQeiuUFmJB2wSgwSJS5TKz7AtAMYdhWZf+Xr3u1iZe6W3C2TBWJJVYcnaAP
hkTc/AwM/Du2GxB5BDp3EXJSyTXdU+BhsHnIT+xwifSYyul/D8CW3Zzfje0txDjyR+QNROnAaEIr
qoq3D2HVtt5Pf3jaswHktLukBcYmr+GkDsJ4YPROWBxB58oThZDKSd01yHK2FKqankk+pNDKwyMd
hN1OqGT/PfjY2fEbxSlvXdutoYTX7XrzSZS1oX0u5tz7lmwLsYiIIhLNMcQFENeWe5Mzfzf/w6wF
xBDlJEZXLvgVvSugQy9bYIPStl8UxVrna5k8AKSkOaXW7fC/cub4/eReszHCIiNiBWNhhIuwt9cJ
3ZLrfxaWWC0+YrkEwvdT+TjK54E1pq4beOIcMzcozYQ/2vxASPTe0UrmxZldrB5O44g1JaFbRaMJ
mLFQslcnU02WyfyWc2IdTmfZO88d1ZaUge3WYa50LW5ffC/37TEE8yi2acW/5lsbgjbuEd3Xa389
9Z0IXeuTJi3ShUVBUtbB1tT5lemYn7rNcP6VoITg8vC97FV3qNWYzT7NxkXI99uP/22c9I5hvuiD
U7B6kTo9UqnPX0h/XM8a6FZuVxp+H6hkQQOuBwZETcMxQqQ8hK8xfXHkiwSF9xLM6jajKQA2PFvz
w2Deejmua8Mtt5qLbGiqdqIHY0yQhQ/1LlA25Ivv3IWpylJ9zEklERKDxWWF2gpsG4ctSaMxL1zZ
acX+O6maHoAEC5i5yq6ZHg+5SZYgHXQsMRi2Rd1Q7MEhLvsCAfDisJoO6sDLbGCrXM3e0KdTgjP2
AnhYxLl2gvtxvBD43uGMrgtH3cJiqA53kjHvREl6qQuHdNiALzN+vIYhCwLUpoJmLBZrqZCiMRsU
jKGkriyRiKssCj8xbnDucC2HJfhV+SiYSHfJJ6K/xYKCT7nmquqXCzmKOKzaGHgjRKolt8lAv56B
jvXbXee7JJOOJyl9jVfCRRN+b2b08TvfT3KwM4fPfQ8PwcPPpXQBnDmZv0CPmP1W5NE+V0SXF0D4
jwSls9bHpCZRc0eeqCZ06owsI+NhnvEDWOoeqxLzFrd9L9qEhXO3P0ozNSq1pkkJTuhVrevh5wg5
P5S+E9whMVDr/QexoSwxwE+DFFaCIVrxYsdk3QCnhje2jeItysGXK3aZFBBz+LVTzcBJrgoljCR2
FI+7mCkiCDfPE3p6UWEoC62PWLPLSZcf9TdPlNZ6xU9v8O3PFvjz2ZaEEZM3vUyxjzR0BXatVliL
Vo5I+F41RpvraPKAQ4szfkeoyTnvG1NSc4k5sGmt6QMlbuug4hcJNJPMltnpX0RGSNUE1PAb0lp0
StW3TiSoqbv1TxlRVN6Suw5zeBVGYFQezG8cNXJgYxSmp0CEmELIFo7jL8aH/WYuUHT0ybJNn4yf
ZLR15LwZsuHuK+ha3I8IHOyxmv37mslCsIJ+lvmIw50iOl5E30/ulvfTKnypZ4KaJZEcXb9uJlO9
bag46otVD4qSFMH7Vt3w4eg1bU/wVpdCidonpFFhjMt9+SYnBzBhImPM4ZndYSl8yv7x19jwh9Hj
0G1vqqWZgxDYX4qG/g843+RaxoW7IaNvYhOw7EVjeonhI0MxeSPByRVcK3436Xcx2N9J7aN2R43I
a+ENNChll+CXf3uWdoLcaaMl+pZy9Il6gKqF9HbbjUzajFvTA3FD8mRxyrsUjLyAHcPCx/xpO9x7
swvqDUGgtPYujyIGtoW41Mlz9OIPZznZPFvsMgxxAb9f21vFNK3FJtySkM4Qy2Wt6m16EOrIbiNq
Tq2x5fSHcd1IzHqByEjQ1gUGT257x6QUJPCUdmq4Whfuc51XxpcKiUbw5vtBZQm63iqAiMTeL3vE
m4Qrf/wn+P+4PqpQdnDEPNblEUBfJDpoZq9PIjiJ9QRix6i0MuR3yzLhnctZq35NxZRqZjz2KSAT
Opw/Rt/of6+q8LoIXc+wPcGKtCojXCm9BrACEvBhaPj6MQr/B0doODeSD+diiJo22xfwMQmxrfPK
8Vxj/8pQhZzrsdvyg7AFRgR1jIrumYTrlaVKz10wtZqyVXMcKmvmpAUHEYjRABNvQI17bGzCtTP/
Qq8GAF5lQdL68gj3zjcCOjp2VqSDjpYXfESuafaKb+arhNNwTPrwB8Xfyq2A3BzqBAagymSoEqX7
9ZE9Q+XfobjBFHDH/4MIYSMLJ8JbjPvPPiM722qgVOkXfnhI89EKHSxMVc5REZ4ra2Cj3GkLM4Fq
goLR061URo9bq81/cqiXk0igC1QbxrkGY/wtqGFqyKuOVwSSE8f0NRm6NRYhbf2jpNRgrM/wKjRT
VVWUUewCRXVtBFEPBc4/4ghU1il5tXtP+JAeZ6xpwV36ixbWKjJnApCKbRqPoEYKOpXgoW3td6MY
bQjmypeb+65ADKH9Le1tuTuXUNI69R2k5pVt3eh8FZtKbXejf7i22xodZkSZ3nGHFsLud/fe0xCM
xicezhYTDEy2pQ0YOyJ4tnGaU31wPgn05N5yRVzpnqLgJyaHZUTEoy8ufMdPNwu/vgqz2z15SiBK
GOFl+32CeR9CxNpi5RKgTWcQK10HQIldLaOY1GEyGnz32ruooVlNBB/nuHw6EOFHNV0a1j7QXjH5
Chg/5JE625bXV/C7t54uh3oLYZcoU/6ON/rUXrnp+L/Rom2ED06k8CYyxNBOKVwmmj4X+bNSJ2iA
PluJoED8tik2qQpWHIeZHPN1zPMxNEwZ/NR0qS0UKJCIRpM0wzWjYWSwKGTB3iJTU9PU2iSiBuVo
6W9PW2nS9Rg0Zuj0ttv4l6pnuRWU9is10OaAqTUvkbXif++w/V1WWXtMZYVzCOt0PP0VKxFYlemX
IekDzisZdzWFlk/RzoHHGkvUJo23Fx09yZCQPMcmKMhCcpfs48F/j7vLvjxQ4dzVBpz751yA2bKt
NZF9W5uN1B/OsadQo7ISn5bB962+dRvkuHzGN9Fll22wxXwNfZ+TdOBmQ9RVVU54XZJuLERGovks
T0qwmO/+3F3TZy6Zv0ZE8qtW6rqEfsTz0los6xmbIn9f2PXcJuJ0DjLenCBH44uXA9q4trb2a+aJ
AO3JtO0RhX/tl2XbaEsKdO1PSt2WZtplS9aIqq4SSpZk4twRbcYgRpI4B/i1usk+2OgY9cCfrSwG
tIzKkFQjs7pjCOEJBc+N2vxTI5f+AFB6iWzraRmPDAlilg8k8+8e9UYiTWCTDVyhEaYVDNXbA1uA
6VliHpjYBP9yK4kgF17Wfof4bPkw95D26RXiPdi0ezhvrIKc/8SeS9Xl43ZnTBnjzatM1BidHo//
31DgufpsZEmvgw97iSsWSWR3TKSiEiiBL7tiGr06tbrVW+idQu5AKH/CDmovjOKDB/Ws/Aq5sBH2
Ey/2s9xdaouF6HVEqd2pldX6DauXpcBWFQDkg+3A6WYj84r25TDCZbTjID5DMSk3JBr4UAO1nlbK
WW2w8bnYpG/jSI6m/y+3/eODEtuQJ31vXiBQej/DeR0Eg7EP0aixSQ9qcyPzjsdo3RauG0feoOMc
2Fd9zyX08n4kVgBLcCcuUdL2eX/xAQLExhvb46hPahVdA2JHXjRSeRXWt1GngSnD5ay1ImauJQgr
DU3jVsdsygKa5JDtTHwBILh7fCyem8hxc0X3BHiy1b2Qcph29szUyQdMrWq8VA4NmuLIZUFvNt1u
4M/VjuQ1UuGZT1ADFZl2/ViPRJ1s8Ah0SyEdS1hkyXv/O4+d3SrTGWaIlQvC1fLUhRaCC0AGb6+w
vTkbWiWcReLoTAi3dq2kggNsRtO7hKY2AUyzyqYzA+4Ap++Naf22qtkcVmQm1ZR2JDr2ZujD6wV1
L/nHHT+MPXLGdUyNm0/VhbqItmpi7ALLuv6DvpWrgAWZ76ibGVQjk1yK+3bk9AwmdPduvKBL//MO
MsGCTgODfgA27UFUyTSoblkG+Hz6VOVf5vcjUNG09zqM5iICfnvyh5Im4XH9MTsXPUte1qNQSuia
lSI60j+w7HxWHxszj9hGHPegTKLk59JExj6PbrheILnmDxkuVpWvtcnqSsPUM13hHKuXN6GAdQe8
1aPz6WLrNFLq5GzpD7bZI2vWzlwgQZacquTS8TGznVTbumK+R0PIOPCgTTSJHD+CKo7gNYhrQyar
ZqSPOHTCejWrlND7CRF6+GULV9xNTosmWOPXGRRWPEceDCn3B0PmU8kJK/Mu1NU4xObeph8M1S8I
yiAd1nYfhD/HEjNFg0ZrB+8+yTik7Lx6NXZh/bh9q3NQ12Ch2YNzdkIcUYhhABrH+0wPhZfTEKDP
1XnTgz2vwrpSuAlVpWihYepS6Moen0kTKtPpADvojT/Qa0hRXDeHZvZNJKdwHFQ3JSYqsMZ3O+kD
J/wN2S0mWB2MlaWY0DbEPlsn9sWFcBcaOx4QbeBcdOP1D9D0h/fFaa54FTJTP002hEI5Pflo3fOi
ArZxeSzmE1EXELRGGqFk7+hTHKH9Adsny1riOXu5cpuf3uR71owJxreeXLZyMciPTDYotwS0u/Yd
WB84fu4nA/WSEbM6kO7YefugHFGkxjo0cqWenpbSygSEo7XKyoTgc2WkIPlaxIG5RLUHqD1eMmYo
Cxk42tMODYD/SQaIqloVAQ4GA3qzg1lkCGa+yV2P2Zqpl90fdzpFedCDuUkio0UMNr3QBU8UtllJ
KCinCP1Tv4ZjO7eA0sOoycHt8J3dDC4qzQOOKQR+KkL5SDmBaTxj3+ECyHmedkcWT3cpGv2MDaMK
SwYofk7jhxLf4HiF5FEXrBd6Q58yiBgaEmTqs417BmiSoE+dvs3qr1GRpXd+3FZvLJE02kqH40QS
gAAlY5WcrphEea01AvHsTTcnSbCTvfGFS1WZ1qAUi3ZC1JhVRJQBZM1vBqpkZG0RscDgFU33I+E6
5ree3Pu7NIdDWkyVvbWLzH0aKV2YEIOVwbrJb+dW+VOYfR+uzO1o36uKXoB8QYaqqljA+RU1MHMO
rWt+UhGR7FWIq9XAv72gICC6lGIGPNj0NDVxWFkqL3b2MXP1W+K0bvLVcaxNa3oyD3mkIKG6gf9I
vM72DbGwKb6Rw3nw6wuO+UUQmnlUsFcCgPi2wdoEhk21eYyfQkcSktr1fVjWovDqkJamioze2Dmp
vK3I4Fww9AygjW1xyLs+G/oesIGAaZFVKPaqiiEg+6bAS/puMENUC4KR70cg+ZQCS87FS/KbVSFj
CbdtXW0fTCELujEFhNaKEs52Q173z3ip9y827MFPj+7OKMx2nbtFv7XSZzu6fkI/l1TwOBDIH9Xs
4tgJUbV6z414BZpPTxovZcwI6SuG6FTzsrYVQXToBPtgfSEUTSkVjwsZDmy4eLhKzSQfXywRsXJq
2rJuKU9wfw18i//x4XqyV9yR1FHvB4Q0OwWMhW+fVMKTN3ydz6K8O/S7rsD7mBrj5kY28THZH57a
O4NFxVaYLlnkBoI9fMSyXbDuAXU7Anultj5A+J+KrNs62cy7yWRB0TNB+W/nhIQ+73ALOcgEAEAm
mOvr14nGh8rmTrpZFW+8bm2EF+93EJjgCSu3r7dZswho4AWr6ykjK5jxa5JQVnWA+2MUorxBBvzV
3obwFAOROSpU6+fxLuPwiiiHRiLTItFAf51bwbvOl7Ah6seXOJKwkIaBeRiSMYZDIIIH78XNOQ7w
EO28glvVMnSNPeEJ2nXIBlOqcGUgef5dCrRF9AesTe0BxgM/6Eqdj2GZFe3W0pAihuSgf5ZcdTjl
Hl0ycBcw/psSRJ8649pai9tTPvR8cN5+dttlGGQ4H59Pit1dWC2WKugtfJMSkR5/2zFnzYoYxkiE
W0lQ4QeIhVcRIWybntGVg5oYfKY5RDkwl+tRs5dPhUpMsntzfaIkFVQ4qXn0gwuTweuEAoBrWy17
ym9+9iYVgxSkC21JW9MQWitK3VkbqaWkt51lQCO656DAjY0YBDbl+Xz0m20we6X4X5VsoNxsrd79
LPL2UHmmzbMa6sUJOF1TDPD8fANA4C369wmzTmMvwmIQDxwxHM1ZnNDe54vWr0BqxBK0aYlGT0ti
DiZzG5Z7EFL6vMcNOkkfPP3dhdzrlxp0iqtQQhmV91LQwlljbHiIFFk2j/ojeqWLZw4amJi/4onM
Drj2/8hURAae5aFniic3JZMX5cKhu0fHKdq5DZao5ziX6BERvxxUJehhr/SWI74hbmKfByKxwMSM
nT4S1dr9WCvVN7zqJI27u1XdMbUmLqxx05lL8gvw46zBHZhL9fR2KWc7ZZDmv18y/LTWBMFzJI6t
BYcGLEXUwZbgBhiFyvOVC9z+SE0ToQJFeWzUNTqpg5YBw5P5YBTgUS+N7KbJP6xYgXC65sD3rPLL
6BuS+RRcaXTIjOlHyr7zSVyMJ9VFw3dZYE6QXe9X096H4yillSpcknDpPBCvJgTPRe+RpPvwbUbq
cnLvmjJQiYyuDIwi31oqSPveLdBOPYCb+BtwEVu6qEzfexCardMyZrVibjsJOTNCzVvD25fV48IK
i8jMykb0s04AF7n/24uhcX2BUur/IjG4EDwXPQvxniySOezpZR4yqwBqpvLvCf8dAnM3UjFlfjxQ
aXnZ1ASSoIKoPjOjfDe9ZECC1KPP9HOt3AQsDdyqeFT+98w4AFGrxTYMohBZ1Bs4nmKgIfscLTIp
aS/WAD8Qi2FeUZhB5MhCUgWmUOjgG7KpNKQBTszCCPfQbyypH6GzvivtJMx+deUTBUxl/fzGwv1i
x7ARTuaYioxNWCVtl+wsxVa6FMEbzyDBL8H8WhRS5LuRErJAbhrClayX3axrCShfZ+UGx7Uln6E/
z/hTSFSEs8CuyVnWhf1FaBjuWCd+ILmJjN1wgVA4Y5qbX9y/Ui/l1YLPWrQo61yI6x9qPwsrZF5I
P1zcklreKsqfiBZhqdmx5OWwRGMSo4LnN0dkVsZldAhnAcMVU9yFqGMgx9xdURkpAn0TDaQWmCiN
8CV2YusdJx0JdsYX7yYS3HqYSY7Jqtg8vbOz8RQjmi9/jPJrHsiwApyNtcQin1Br1GOxuO50tRmx
QsvkJZBaUsLSeBHYH9V4x5huAY+U9bgyIKYqEdsEZTw+YPzzkKV4qjX2RZp1ugh7DHIZcltvtgxY
VlNrJkJ6XaC9iKCBoBDfM9BplTcxIOEBdPtdy4cuxD/8XzbClGoBTRfY6aoMzD1SB8RjZr2r2feX
fUTJY+ZXX31cR7F0tpI6pMMk62XRD93iPLHFwHHx60NylWRzgnI38UwUudd/pHzMrOBP9tfVM43L
Hh9bvenvXPFuS5Wxp5qehBSBCLDFT0NettwS4sMqSinGXg3XxquxQzEuSmWKeOHt0jxYD3g/HpBs
/Y9WmAUei/FcyB9lSQ4sG0sWYoUKJHIj/N24xX7xl7zkUCfAjXG6/Q4v6t8EhZ829t4Ni30IhBnC
GYSPSBH4FWPw1pnpqcVXJaLskTzeIN2/RvRYxMM7NTOK1OqZW9hvJcPKop00NJa3hIpWYb/pJMR1
O+yhxriFLvqPhpewl1RdPWFrXmWnn6I16aiTv+LXEC/OYs+arPIJs5WP2byGuqanYrgaRI3BYulh
4wUrFnH2WcN0neN9efjUYpstcAg3YUOgUTi9WSKHGIaleQvrJHaHrlp8Sy1DOB3UdtMisvJZdGJB
25KUiSN5Qvp6PnAa9AICmOtQdxxxFugOI6qwlvZAsuUIHiDAgmXTjNXURcpizXt1nTWe6UsaHdUP
qw/BVLv2Z45vTvwcfSQuUdSHijpiARhgbXu0jMms//BdtHvKn1bupG371xv81R6zVVp2Gfn4mlhV
pWx56M+FSrrYAyINQoKblrLdbVHnGCOS/Af9e+xKL4SwsVtDfur7EldMranb9CRlCSfO7W1VweeH
7LU3sAt98ZWaL+FxHHANrONksIaZ8JPP4jOrdMP3OmbUiR8jdxqDwXPj1k/gmMNJ4NSTK0rLp9y2
5NQ/6qtomtv0ufvGpZOEqLksqBbQdqwRCSDREAIkDtDCSmZBgP5HOtwitfSp4PPZV0Ko2M499gqi
HD8zuy+UUUvdAB1Qkw/B4JO7hMo7kpwmeiJG8xD50BFWUOt6iOPOZTmcbqWj/60aHc8ls/1+hhCu
keN1q3ZeX7GXWmS9j7PU2BIot4t4N5rXmdU2Gj6uHeGPa9B61/KFM2SkKgg8W0t5oqmj0ApcehzA
77b07rckkc5Qa7R7+QJQlchN6Lo9Cd1Jl2Alw8RWT4Ta4Yryhd2BNUwgfXPfYouYVkEVM0xnvKcO
FcC/vcsW3AU6ChlS1tCgPX5D73KlbRMjBPviCb+zY8iKamy03Yqy5pD2+6d87KzcHUHQbVGdY4DK
y7lBlCC1NoecNxsWjUKta5ndJ5YiANLEcoqDRX61DExgSMP2ajVJYfFPgr/C9dlf7iWWGJcASLEp
5l0Ft/RLAgr2vsEi10lL6UUnvqyTL7RY8la4SPBe7eBrOvMpo1uFlsV961o9p5ixOPJn8K0a4J4F
OYh6/GhWJvGnxJWpsSyOq8JFTmkgwdvP+J3GaP1bGjz8qSUcHbpAwhyelkNEy0/eOENl6KbSODqd
FMWagGe5+XWJxmQeoi4claw//GQZhMm7VoP9vqtMc9IDQPNarOCAFK++334RyxKTtnigN7qTLMXZ
bwZ6MbZ5NTczqsfiPG7TXsEt16Shz3wNPiHb0I4yTK1896aks0+i6LjCU2LpvpOVIOhu1hDh41NK
GvinzF3DesbdmnrYymRRNNQhzmkYeEMFIkcWzyE81w5doPiLgkS/x0YKKYS4H2vKDYXaF1HY0iD6
FdESnQl4TmUnKl+r04kNFQzCNX0zpKYYXrciLasW9NEKKNQw3xPcPukqwziuU4XqNZo0Z56NN6v2
QEJ60rFitAX2fGa0IRahUK6xBtP/qP/HuudjgVwpJBNyS4wYaJNuUPuLDa0vAJm3iZZdeTRtfAN2
ZRyYkPjC7V+GMBBtWDfP9Y0KeH7rkTESNFGd48HyevptyPk9Hee5xove2NihY08zRtKTxY99SYdj
QnRwCFDE/egx29mIObG+Gu40+9cilXiOJFOvNkbx6UNfWt8xp//aV2zOGjD5Bjc9a50BjTkpyoTy
kD3fj1webOuC2pG03ZyUYb4Lj+MKWcaaLZIRN/wPpuzfXdWo2AQCH8SV3/Uf1CJXGShDvivnPPKR
rAN+yuuCRZpwCaNY2HaQFzdT9kfCTIYyeOA0ja8IPM/jPYG8wb8u3Mpo/ZT0KvbwBfgSP6BCIXpM
z5+J6eYRlxZMYqhacsGjcGTH08AeVTxiF/312f2OBE68EaroNPk26qBMV3DpoEUEhX+yQSIHqMuo
76SRwSSugC4jbWElekYAKktlMZZDCmMYJH/BpJgoTNzNRoE9wQLrOLcUVTqpV/fQdWn6JxXn2/72
xBO8BltUBc84uYusvqhrlqSII2mWaV7/X9Ga0rQibT0DVWc5nlE6P114MYIGkjaOP8XFZkRCeVZe
fMvXA2zcfuKSINKBiuyBz7cSKh8bY1JL1NJEVvOd1RHHr4DOq394na0OAnfasnPHe5Jf5MqIVsbD
ze1T/fHwSsKv+jl0UYDUIAP9WT4zwsbUi+YzRLyEHY6+u0CTAomvR3AHyRM2+KBn+TtnPuI/i7xQ
kuHreidpe9OKeV013yzavMSPBcw626OCxiLkO7vtuKje4MEpz9KWS4g52O0UnNq+O2aYB9Wo44Y5
XPbM124rwqUzrK6uAzSR2IJahOyi3Zat6ghPuqw6QNbXAxCgM7L20bDdDO2NVMf7eE9FTf9Afqel
h1rCHC74ZK1XyAZtxWoOOFRjkgqZx+fy9U1aM9aAVct6L0+tVoENrz6k1kLyTU4iYvAYyeuiOOla
jznBZMgZ6Psv8Fy667UPAbkQnN1OkpO7bq57aIfoQqjepwySSNRflZgZnkiPXTU7/rsnsHgUYywT
UhE59xIqyJsqw2LhuBTS5q3i6fDL6LMeI09PU9+rNRytdMyYgakTTcTDkJyWeNqTsJLBb0c5eki9
Dz0v5cpn9Qf8Grm3geRt/pk4skXwq5Ukw0rtaidMOI0WnCmlbEejlGDVVwkROMKCjJJ88U45FoKa
Sk/3UEtmMb7eEGNcj7I74r0EoDno/xLfFHUyf4Uinaf1JQCTw1h/MOFJlM7iSNTk6AeJkJ9uAKel
tYSC8FzMUpZff48EjUBeW1zBgNJF9gmKAJdmnfMqN+JQdOrRneYpdt/e6ZqTN8Nqkh0X0vWn6Jz/
9Ffgde8hOaJtHRWiTA0QDCJSXIIblcxhzIagKXqCF2xDUhzGty/JUZHRIUuWCfSvRo84xiFOSSbb
pX7BPyVGQKnaW7Z3g3dlDTXsi/4gn/950tadm5gEaf31lHRPBAKcl79rrTUg3oo0k97XeFfQPvuA
CxSsuePeCeSxqvW+f+D2LXPwtnOegNvJBZNpbJM8iEteOigNpvTjzWu4lgAgU2weXgr3D7dP0Q/y
PAXUT66D7kj+EZyqmCe4L7PMFKT2ayKe+CrG3fF85k3p5eq1H/3I/qu3RO5YKGAeHI6mMsNTC9s7
sArmwnt5pMjDwoKTtzCScofttR0LLgLYQ3ZUnn8CZoJ/JyDA4It1pesO9u+YSBtx/bgG6rDs3Va5
I/fTCPxEkm02Uk4NSNj0YeWrXpgauYZHZci9RmZ/9jVKyiUDOjD7zybfWtQVmf0E/pUCrUTd+WTd
N1lyKNfg84qBKFS+EO0xhyWazoenDrJ60rz0dKmIpL6bIc6YQsfgbgdB9KFM9t0OZ0x4Xy95hFI6
+B7xfN6jwjulZPWeYB85IueoV28A9w9tEXT9XIW1Dvvk3Mm6LG3oVqL3HMNg/P9F0oXbvRB/Qaih
PDzwKgvOG5B4SJp4K7pxw6cAM10Sj0lPYeeyaRwsOGXCOzqARrM5Ic6LY3ThRBeIqb/rwzwKC+g/
HierQqgZNZGnCQ6z8wywBni/ocALKJIAMYgY1g7vSNGfZEH/KcV13fF6xigddSNmTjE+/Fp3vaBB
SbLQ/8vE5eUcwIcZ3R3A6TswNgObctCZ1o91hRWsLSbUU1yJv5KkqBFYJxL7INOpWwfM33/nSYf8
O4b6bv06r3rsJrZXOAK2ln2sq6Ip9XwNDmEm4NYF49+Gf4hl+wj8gdY2MppNnkPIg5cGJe+WUyFu
B1oY8o9TXIGFEI08u3gV6vlHjWBxZ5tFLf8zkEP4DwngFdQFhvop3nzv/Emrq3GALkKD8FhNs/Rh
dqgZrUSw/p0vv5DgxYetS1NEOodwCgNph4cIlVXg7ZXCpBGnfViK0QER00arC7+HBQKvB4o8HUT+
xLYWZGiIlmJGs07QZFBVFU09lSN1ey2uvyQtG1DcWDWSnBu2a05GjAwqZYFLHzVeNLwLiz50kgZ5
reyePy69ED3Cbx8WrB31BFX51FY1hxGWYv5lhMJOpDxUck5fkwYwbD3p/1oepw9EkOUZXx/btVzp
qlCul8gjh/afih3cDkmldS2msmmBbmwnw72VGDaILQYFA/UVueqtf+VNeOiOTZEun0Ar4GiXQHSh
dfjRG5FvR9HRSNOcMyPWP30O79Fbj0Jv3nPe0fz6SQBLERo8OVw3nQ4xIDJDLtPipYoxVT3FupyT
4sB59nkm4/0AbiodY0tFCe+W1ygXQh5w5QahSyM1QRCZzit1sAbcW4djdH4OttNDB+2kBBGroydo
yEuFO15ZxQeAvTmUVpQj/x70CQpSSbMkzrVII14HnWbuiE1eAhMj5Eg0BbiNgkAKcH6k8q7bicP4
Vf7BFth63mW+qIAmn5k+nVKcsv4KM7/eVv5bpMSXv9hOWvhstgKgK2vdXIkcdQZqIt40W6RpJ0nr
TwelODIlqvsdZ9GWDEX1Kuk/yREpXB6lZkGEZBwyBd3wsCIKkgdD6VRrsqXIAPn5Z6I2AOy8Dafr
HE4RAj6MizuJCL6Mlbv8p5qrI2vJLGHiPwfN5v0qUmdma3y7kblxvDKEksOaTjdBCE8+Po9opACt
PszrvxbzVh5V2dA3SkPIOJrSl4m6ubrrnMeaLA5fN4cTNcx2xSahFeJBxqujyQgklBUC6KbEn/y/
/nbTbSvLsLyQ1xGmMeQr20kbFKbNXLzVXeY7H87M3H6721s3cBT+L+zGnOwXFZmhKE6mflB2GgwE
KZiWtHVUiWyZVBGFnPVOzCssLJRnXdg+1dC4CPbuWY5SGQ6Ly+j9tOosAIu95O5vh4ECP/EY/UMS
mfnCD8kJJ6ClL2qmGQ3cyPY3qxe/8sNZ2u5/BDNfeMSlzNlu2AOECUBOC1abvy19imPvDXvaZA52
XdtDJghuPQR2H5HDXNvG4ianrVes+k7BzAKvHdZNxDvMUXrhe1e2CkxxEu6+1n5PufKAtMSOpAfQ
jzLowfHePaqsPzgjn9ciAYeEVvJsIpVUCgW4zNoHHXa3WjPXH+81CwvnjufjovjcYLeO8sDoi44n
8Ndx9ho3M6FPvwTqkdPU/j3aSTbtP/02xln9bgJn7Kvj1pPvrIfN+7ih3FRcZFBhPDlDQOHbRO4r
DqbnzOfzPxlJfbU979uHDc6Pl93XTH7abhjPoK1+L44ewZzv/7J2ABpkIgpaiz06pHwhwwCytkBb
Cfj8ZH6Xv6rtxDFlKWZOEBUNR05XxWwRYrg2tx3MafevbeW+OEAh/tT5Bl6uAWWiGd7pGguUUBW1
7B9WiiF1tho2wX7Gy7N/La75harbD0asiQ+s6aB6T0ZnpOd6OmyRr918pIHKWQXB0+5NeRxXS4gN
TH+VcS5luTM6PIGxsjq7PRJ7sjgyLflSfOQ4C9FutgNbGZaSDlvDa/s4hQLf52oNBZUMAfx0aPha
zKDepO3s4t87+kDCdrIvcKWosVqRMcI6VNODfxC1zHimNQmj8YplsG21KA3lj28wl5aFQrZteNu+
/S2PJC/WffijYIFt/lNfWdZXz1mXGLV+5y3qkJKg51UwlV3mUMfQX9NfmTxUF7rtWRnUwwbXnfpz
0NDFbBMLEJpzLCqi7YAfsL4B36H7R0O574UTg5Bzyr+3/ogszvpCd5JxaEHSL17X1Lt9eJ7LlJiU
3Xv3NeVeYuHkhqyuSCteBl+b3i4GzSB5fQMvVg3Uu21T+DumxCZ1fb2n0BUz1N/8D3zogmzVCjkX
fWjfbjFRUVqsOVLTcfNZi58K0jJzaa5YF+K+tJ9weS5KI43f5rYFBCuFSyIe5Xsj/vAUbRqmk9i3
nXXBLYHhKRIFkSDCgdR9nEy89/WnB0MvYOqcXIxFP+7YUL3CVTYCplXKTjPQ06Zz6N0wqpReKW88
diYnpowUqD7vifzfmE0AvD6YRRIGq9XXjZbL85o8D1QFfjPGA8NQHaiYIjerwk3DUxAiXkJbyp6d
/HxE9gPkzyeQuSuJAlmpQ9jUffyMuTU+RYbeRciS7nUpdc5mA3ZP9xrendxgmZpaxCd/3PaZXXnA
3RzqCiGUV5oDRQ1F8RZz6q+sulzU5+//ISwxb9dztUJWN1dm1wVL5gHk8qzA0VEWwd3RWG5BRZb0
ZRjcozwiqzKdnDM5uTD1GcWkPRqfzB6T+qNLQtz62dmXJne+FLYJWr4ZRg02jhSRLMSqclPyEmeO
5DwI1gb8CQYM2r7srBXplVDB0P2H4V9fEqyPOIbWV5b/O5Lq73YwHMJLUHliSIkvJoiJuMqiPk+z
ViQHyBAgQY8w+EQD3O18CLNbgmI3G2YjrF+waPi8QMWVJ0er1Nkx068p+wyaKTTCzmQVJLyd8pHC
TBwtecIs+OGCK7lWYyWObb92gIzqB0sGUmvy98sNWEuL+gm8eROuoaUEyoLp/Xfc4H26rilepAUP
9ZnSpGl1tG2dp7bSlI9Kdtv/lXJW7ZEAR2E89w8TdggrHGApybeZssKvnj73zkawH7KMWw1dD9M8
iagxRhiCc9FKB07VeKug1NCMCpOnluGBIjP5h/pXcgB2xDn/qWe19DJdqUfNIfiDIIsoxzN+r26p
xN7m7qMJo2vRBhWOj0Xm/bS0AHYhl/1U4Z3tK7pnFy7NUtH31p1DZhdtKS3g+b8kk5WXFIaXmqKZ
4m1Q9Q/zymrBSuZbbqRv99H1yoqh6PxA0RmPyxBwOztR4SmtZskEE+Cos2mj8AAjSrvFaupDatji
BVXtRsSd+dS892kI4mZN2sSZze4V/1pFdNhG94NwVpkQK7WmDZAP/GSo9Yq2J8dZsIFIGI2j4qKi
J6cKF7wDIEWTDBuj4TF1Xk43ftZVGol5tz7mjDcN+b/S4KPATZn7UQk3GGhEBfkSgKZx1TUMcWsy
TfxuHp5Ca3TIplgaodGw2tpiQ/Ra/vGrZ5FQQQRxmfXSIjjyrAYmXk+RnYR0bewghPIXpSDU9dvn
R7sixEin3Y2t5ddzh9B904vAV3SpInqVmLnmgLzw6M9DliB5Q+TRfSSFMxLxrdr+ahLYq9qELlXd
hshRivMtfGzNssmcPO5fFHiSeEPXflHnnoym0JmmgSPlHg/SflWLLe6SrisVMC2I9kV6E77+maEc
ZQNFG/9GH0yvI1CSBXhjA98VXHo/2bZ9mOqdRZafFhI3iDqnriYipT2Mu5/XYGaN8/86QDPnC9Wp
VEbbRJnsLkcOBRz29YKCtPk6XVoF261IbhcDT7EhVuzI4SZSFmIi0CXBy/nznfUEk3CsDpG4hq5w
SeRVOjLWJGAaGZ0iLocC6rsASjbvY2DQWKx6MErKL9T7jGNLJTxY8jFvJh0uYsSCZM48zCAqzHYk
ESqDdXB2j37y5dcg5UuKD50y6pgthuqp7/qXQLBQRFQyyPeVjCMW2KVUKf7dTYLf5i5tXJ5MPEcA
N6kt+NXkDA0Jx5ZTQpGy1KTpguy8Ai1OhNmWvSNqnOJ/7wbxEbnAcciFBDKb4wEUWYB61GAud7il
+E9MoDcL83ijgWZuLx+pP9OD3aD6kwpB6lOoGxEPp335oVW51c1zDYUxVYk0n446zWiP7G+6Nexb
87Ayc+sKA/nAlZ9v1qSCAu0/seOXSuQuztet0NscMZRdhuMWAc11jdRcWdKtXIU8mw4Ez4E4bRsx
ZlOgg84K/4cNABihtuYORpXSPKqM6FKr54lYGtmfI763uN/P44dCUp7CbsY39REK59ZHMAtwwzwS
rvZAlmdEFQDzCQ9y14te3fH3ntGxakpzALeIlff03P09ISJngre6KckbsMJ8RNDFMZ1bt50VQbhE
K9XD7+PRI4u7/vkQidYb/xRy+HR37qGPkyQwl62H6fIn17E12TQyVhr6a8AAAQ2DT5VvjvIKET8R
S8yeW3HD3ood73n8KeQjvpDOvSg5Je6cTwI7JdZNk3yXg5A5uKWwXsPoKPZ79D6Au0siL0GfzkJZ
HA0kPGCFx496M/0b4ot1abZOKzu7iiU/ziYA9a7TxjRJvJPudluglWWXZl5hh2yMj8k7kSHa379g
4Kdvu8lCsG6/vQN34o0UIXt99AMX01HxLlsRjHXr3iBq/M4UI9fVFgP2Yzp8xAR/8YOK8oLl4ku6
Laqws8nRF+jAUcx6UQuDMPnRbtxlUikeZMVOPA2zCvq/K1nY94rFJSk5CFWakg0zhBI86pv9PFLc
/oJiieHK8i1MQqOhY//Fr6+kTHliHQ+HKnOIkqtXswbuL1nlpNgtwwgGKbgCwH7A72CcZi0tTx/m
rVlLi2v8TgGZwNF2+zwP5ruC8Fjsyt0bs9HOAcUEHgiuP7tpxW3y0wkkKDMPXj/M/BOYl/Gj+c57
9Q6Uq/AJ1tk7qfcFV3NeAJ7Sj4KwazaBZnngqrVOJCR47khV2cVafg+wo1GbW/RLOmjrm7K0MtOW
dCvy3skZX8R1ZeMqDjeRpTBo0msosN17yLnOGSdQ6e86f2Zc/f3Yok2UOpI12HxiwClEgee+QEPu
3u4bBPkP9yTsOQ1P71mgCf/vo6dE6tUZqVhkK6/axLsPBM1BIvMkvqdsv+Z4KI3DObMVFNlbFcPA
MNCJXkOj5lUOoN1eGBjxDeAKYUQv0Y49s2aLpWWgrMPP7r+Ui11mkF0ALar/DdhFWUkSVne9x8vX
9VJ7/WwymDuExxMlgWfH4LRNinGD1clM6mvblkxOKLxlLGaWf0SOrRyCvakheJVC4Gz6JtwgbbPk
OGWM7i+V4tncLd0C5VX/ovE6at9H23KAs1I6jT2oyCr7F52GLnRrUoFdMkbbd52JvVRfDJhn8nYZ
lzbDP+VBuPysF8G6L37td/cjAnM380ZTj2oNDV39klbxxfYubrQIBAGokgOFhDL0yyBKjiFBP5/k
IlkDWckJHtWMHEg1wckgGkqfGcp9AV/zlVLLOD00V5r5w8uYc59me8bsmmum6LLOYlRoKmjtxcA/
KBtawwGOi7ILbpD7ePsh1L1LTnLH/6KLMEK82dnuA0v791OtLTHeIfrGSc1ClKVaSmfgWviBQAPw
0KazdwiYE0bbpgCwroJ+qHPzdm1hCimBSkuCUxR8cv0dSeiKfKFGFbsVgwy2ezAWU1rG2FHadxBh
PIWh0Tc62VAnvJSdtvhgmbHJ+DQ0d9qc3Tcr86VGT3BRMkgDqeR6v/inlDBVF0W5yG6TUrwRZ0ks
Ny107jva5t89VKfI5P961IPFs1ehxg0MvnFyIhvDFuZ+mO47zCt/nCv9N7TL6tYzPies9+p9nJSY
+ApNJ4U1xOhU3S1WWZ2/zDzthUDB7zagthaMVxEyyL5rQl5OqJLuzh5H1oAtm4AwKYPiQeWYFRDU
WMQORppxJOHNu1aAq0z3UsH3lfNK7ju8F/B5QcBEtIZErmOjCE7HqvAM+cc7HmTITJaiBT+siH0a
+EjfvQ6Zmc3WfIzv+YLDTtjK3SD9Tq9ksyiAkfq7t2kheNCS7HMPNtNASSYV18UYP30o9TZNzGwK
y8rTVV8oAyMKbxd+rgWDKxPgCYqqpqY6h92940owSSc2HzsbE+2MMBHZUzRUwQXS7Md3A6XZBHZ2
hLxT6eNipdx/G43FkA2w09RXjc7XAJG0FxKKaBAGtYKOyBgSDcotQuPTBwJTvW0/fekhIMQhI8Ns
Et74UB59z+wraaaOAs9uy4PZuoknacN71rw3yPFLZePX4lo58Xd3vEogPCGZh5hGEW8zKIXLlwif
QWS1p0vddQl/i6dn5N6I4lycPuydDrieab13KY9RTgpfV5ZNY7SbI59q8PqKZKeGL5eIVNPthNMy
bh8tZ7j8gmNxkLz+efPHPudD8mzVFy+dPVCvxzwsFSa5PL/WGj66fasASqZeOwCTmlocE8bQUR+c
XmO75tAt7jEdTOGemsZwMA9fwzA8SXQ99NihfvJtiQ3kIhbhQmxhGmP32CVPZpO7SeFptp4JRiJN
jDYvALTuGd8pT2gsh3cEWvrK4ZA3EcAD2Xh+7Cvofm/Pj/BTMiupeNusk7ZuypdBf42F935FvXFd
/iRzlTR+gvCH2QBUOt1Dl7UMehYgvSSBzpq38OKUZUfgmH01RswQFP+fZ+mKwG80rsk4P0oMHjFL
+nF2cVM31wEOLg96G5zy7ShYmKiPAN7JqA8CfXnAHdw+iVf76iumqYcfEVxY8QoMIjMiI8CskZ8G
mEI4guNs9BtVzW61ngmpuPtGEUwl+0XB4EpjzijdB/La3csungVK8b9bCexPDWW+4iZRbYXd7FVy
LPvuE/okK5el0uW3sRGMqi5bGuBSWynxtvt/hzOCaFSEkH1uKqH4rfcZAlRUqX+3l9lZk2V9TKFn
naJvBAykE1SucgZ6N+Woo2J5Cbhh81LkQcBrqjt6hecL5cjjy7584DlkzDvn8JXPHugNdQRSYrQB
gf7864O2aUAWNYdcD62OCzh6MSpaPzq6ZAyocHnq1GzAh4X1UB/kgb6eiUbZkR65xJveJrQi26NW
C26+Ukf1T8a5qfITP4lTVz99oRFHYLfijlJeG3B9iLRNmkIaHdni5DqzMbhEowfj42Q7zq7g52to
f1SR4aH7lYuhqXwYVXskOdN196Fc3RFMxhvaR0ssGZOVxi2/qDaCkyY3x8f0hxel2ody4iHjMDOt
s/4RhrKxd5E0pAyFk430Pazik+55DIX++gActQGN2kdHczrfyXGfbcQ50RoPMS2s/rpCOfkTH6Xl
MS5y1LDU80ZOAzlutRsJfX5RR+JCAfMPVkwSYNaSkQW8cr0cTtl8t2IBOUXbTsp9VrYS5S2O8HtR
9q5cKpmhrRSt+xnO8pHcMFEbrIRKm+lR4GLsih1pNiA/UPCjkfI9cMFMh4rsOj8AZRI0JNyMemj6
GhbzidYBkEyhhIrllLdKJyT1GfVKejuWmiYmHKdMoF2yV9Cj4cNf3TmdKDX3kwiTetoe3bIgh4KO
7sUeJY9mWdRrvwI1LFc7fDEcXYRcK5m+ee1py6DGNfnqIh6VKPWnrlHsL/SOwkNZn8M6+FtEE2hr
JzKcvKWX+hbgkAgSeedVZnz5QsKuoTKe4wTloB0Y435XpHMRSaZga5rioYIzhk5E1a/ehmhZEVvN
QlTUh+MTn8DGmhuUl9x6/dvtkV5FnQBHTGrer9+2mn7YbwJWrM3Wdh54XRXWg/LOhXo7ajho4NRK
mTJClA2yvF30liWDeA0xGqGfUS9xKzINxNgWAg0vH4vlLEgo0i/9gX6sCfsvoTu6KHBFB/JnrFgV
IOLlq1zfQnIqQvQ0zcIVsHDmsg8M8YLWv9/AVZGW5/wOA5OUcJOwRW4/p+Ox7mNYfTPzVNoT2Kko
XOQX+8WJvqyEc4dyynUtRPhUPbDt7M97IhiBYed91358P8nITl8Mk948OUjsUhuAG4MjBVENNTJH
X/cpw9bArN/3Ps4ZyCQ01EpMxIhssF6Ku+6f4+NLI2Ti+e0TmX5ShHCipJdz7ig23D5wgOzqjVSV
qAchJkimZsZZJAbJY14m9i0LoBiNKHifBsMhr1TI3HxIweyRyHBOzes/O1GuewVXONTyBPS5tH+m
s8sl4e5n2Rk2lM0JDvFAu13mh0sOu73nU0Db1hp3r0gBC9WrwikPHEdQsQkyWiN9qRevYt7qiVnW
BH1X61f7b6wOQ+EXfw7omC3cYC/rdHlKaB+KcYm8NsyVl1WnMGhfbWlTn/QsjXHYerigedCgDkSJ
zAoP1WVgZiPiQ2fwxox1az4QRUkopchd23h5ZQEVetimGh9IltlHQC4jI9P+ySD0H1JC+a8o9re2
1zROtv+ZKSLmbtr0UHtFwESEPggXwYCgL8Rm4s8EXva4ejddCNYTlUxYD1a79uIzUAtHJ+ugg+gk
e2IFWRsOmiTwgvCNLldDwf2qbimU2/24O88ZLIWsnvY90GWAOtHy/xtAyJu7u7bNumQ3Iagqn9OR
v3vCsxaPKPmZcXHs5istpvcnhnvYB78+IxAWMl04y3gJYsMipZ2YcqfRGtFYM1TLI9nv110wRVTd
YqtHFba01nUl/gKHOjEM5XbsyfHd9PGO6u0Z3YM85cfkpQTzUD7MKSs0b1MLNKQQhLbr3L44t7NQ
XLOgVimeQClZSBJKQKCMbN21p2D5akpCGyf5JUN7UEdlsmW3Ocw8HWhH6RW4TG+ZxiMyW1DejkbY
sd6XRc88PqyWyRp6bJj03iaGt8EzHMcJsGiv0XUohDBEYMwfuWLbmefXmafEp8rwaFSDNa0Yk37C
a+T3TJ4br3WUZKj0RKgwmWUFNol+lyYe2Qgk3DPqAMxMKYcAzpy72sI5WQQSZu5eVo3C+iSXas9N
pBbqe74u6+9jwDp6ElTBs6ux2ask/ZHiXvBaXdLTUKxg+lrCB1N28njX7MBzFd5WROmz6irzQ5rv
Wve9+VwH4dQuGJ7g+ihRKoFnJ+g8MxRp2xmqhpijuvNYIReYEoKTqGgkRCthxjnypSQ8jjeOoRWt
eqQg4PNtRvsVaQ4EpJqNSFEnKvdcVo9lMPkUSx9zzV/eAQSmO8XKstmbF+y3vkk7kskcgtONRRvL
BWSvXAHCeRxRprhCyZYXHL4gvKKA7IRZCbf8seSvHUXe0vSlSZ1omTcYmE2V7VIsMjHMCYcFz2ab
WYo2WMZF4mtzyFxGIWfbfiAEE+fYAP1komY4PRQxwnlpiRi1TbOQ6jtkRPlIy1XkqaFIsz1uk+8N
QLiLlhYQjQPKb+8143QnzK0mFVMSyqpl9V6+sPJxMNUDPkFstFHUw+ilpRpk4s/zHUNTtekMABsv
jkmA3gIazIuBcsjjXIGMQOhDE6EUS/HjMjr/HgP/0hEKtkQdaoIMtZMvn72W9V8NQ7o9jkwVcwS0
+NLYhzUDw4CPGseYc1++Xd6URTpH90ME3Bu5cE+jEtaQMy9DpGX9GddWx7wzSAfEOhBDymVxPEWD
l85fKQoOGt8YK0kIWMRt6VorcMzND+S1yE4cJmue3UoYUeeqK0Gq84/d82yPxwTbG54zhADfN3FR
4uQW82AkLBKXtgeUBH80BfgSfaxRT5eM/0CL5cc9+QlLnEd4Se0UO1XE2UOkAmIveKTG4UVWzbi0
Ehay7jl4NCnC+c80V53DaIMpZN9KnCafBuxi6RvRhaQMEjaOV5FRx5bZhN9IYGwnBkIEJm5acF06
CAEWcwf3OW1Zh3oT4DTQLbbcCg8CGiI8vj8q4FMGCIBVk9m0VWYVu1IdrBeJLMdcfQ7X1LMGQ/F9
/bBkbeeLC5qqgR+6oeQyTpKu0lCdKmJL4sZ5Tia2FSFVK7SOdX2RvCK9dpY6ShjIoW8o8v/efjMt
r5Oc5v9PJMnqwVwCx1qiVpq1E9F6KSZC3kiG/SOfHFVJ2n8LEkacBfpZBYX3KSLhjIg8KhXLVGpZ
z34wWDvyEVTOkRT1CznqgL7o51BbjGxZ3Vz2gAfzU7u8GiFrbOBWZve3eQD9Rwm2M57jKBAUEahQ
RKT/3zEfqNlN76Ei6ly4r7jBgZCveSpf8GX1qd1WiPyfgq1zyX9UDt3LqbHjRchMRGR6rnC4gp9i
z/F8m5H9qQkBKI1N6CVkbIJ+srRFF21RLkYXeB8QfiMw7hl7nvmN6sNgADeVPW/jFfjl4I6gQ+lA
jzDLh9ijlhV0M9tRfvSMeROr38TJ3Ej6LAt6QYP8kZiegl4uwmm3IjOsPRHy35yligJw0644WEEY
XIgih+UTBcCwsIkenjkMnNwzwZLbacXodvnPpVvwDSdX7bcudF+WmoRTqv2m6LiraFGVWpS9ikDf
eLr3Ge/tdUyrpfhrQTFmbcTlde/EK3bnM7667i+M80xVfetRaIKvhBYE02UXOm72ZKTekiFKoIpM
nXHpwWlDxYT/0143Ihku+jVyCbDdgTFEV0grkU2qHbTJ0fzuTv2ksNaU8MgIrd/hdHhsSG/1BKsl
TW+OsFjAzr/dJREWA1qL8/YZOo+L1PRZWJWPzMB7fhuDz8jMRaMAWDLfADpmG9ZMq2ZWj9h9aAYn
kACYlYH31Cgf1NRI+r8gsib0qhtnM7nXvGSiBkZ8wQ5fLlqmmHgY3YW/FEdrDK2j4rVn1LsFdHUo
TTVdFqo5x3LXSv9hxbSWwgAKUgMIMNJ+ty9fRKDV3M/umOppi3GkQXss2AAkfX8S2UJ72J0a18gp
BtJA9WUX4oSNpzUJlAZvp7h4yH+by9BsWCtiPbDjLgpGetrZ5ix1/OtAmBecjqGbIzLFvtNfH9/I
h0+wWp+ITA2UXiODB1DAUadOPAF1ltlJWeKx6MMjbiU3tJPqwGVJCMec7V9guOYi7GPatUvL+Xik
+kCrVlY3m9sWbD3PBaCfTyNh5k7KmQhWzsLCEhMg/JwYNFJKDqVLTueCkFNWvhCzlNiNiJch8XHv
fL5DnxjJjrWjt0krAZPc8WCQtinbL4b8XxFWDZN49vgDmseavfgLF63CbFcu32KltBbyHLT7JY/b
PklFGIfK/izy4cV6VkSUIkWu/BerNjRS5N4ljK/WpcRXuYfbXtbCL5q6XF3rgZQhAtKPQKobEB3w
bJ2mG3FbHN9MfdT+3NoxmgcWqWPlaCgCZRHVcHPV4KbRJQCqhSH89Agxy5qOhimmiK8Kc6rWFFM/
HOrYTrSTZxZ1wx0xgTplZBk9TYgZFvL6Iz+W1h71jAX7c/P1Rsj9R9OjX2Fv07toFnEaju9u7pWv
ePC0sXE8+opoi/NA/96yxtP2yZNkdtdUpKXK6kJB8nVn9VercC7obfGTd489u5Ymt7tENKZoYLnm
3XsHp0fJyu63D63XzD0/0H6MhXTNfufsnONWcvWAbUJAdX8irOY5R9w103GoeUTxmb0J0LVEqBNa
Mp74BB+SkPDg3SjVGSXiAmTEPksrul5x0TXJ0zRtwQf1IDkBcz3Mvt9mKv06x0SjgboAFYcJE5iB
OBs8Me7YzXZupCjXTp4eOwGd5RZvbBPD6QqElbm3eAAuKS56bkhzLLW9ywgvTdYX/gZoi9Ox4PUA
fFxIwhu2/dacVEIZSTNu/NlFRW+bG0VKC4Zxuycb2/7DlwBObw1jXdk/GwVZV/HNaFTyvLguqU7x
wbaVYuE/EdphGeiGqrM/X5Sm6DrvA2huYrB6EMtjnF/t6LFYZEPCQoeuQXc6VYm9yLeNlPb1/rZ3
6JoLG2Y8lBg1fyGUN8gqLnl0Vqyw6vmojBQrBPOEbBWK9ftfzREisvmhfAo45hKTnkp8CjPyAN5P
biiJqwyDVTImehQULp4Dw8adCqf+BOH40iW4Fw6cqZXvNZGAGOC4yoAtyRn9c5XM4u3OfluvCctE
oGXoiHalY1OEd0ho6e9/M1K9eXjX7O+lOEZ+fM0TX/opssoqYA9I2QX9RERpUz8m4kEeqc6C3kTn
boS3l4tyiQkxFEFY6vt/RiiDXcFwEgBK2FdygXAlPpetuZrzyH3JnU6XuipL6peP/Ja2ed/JhDIj
l1giT0BgX34PHnc9QyHm6soTRA2P+iUHvsverjKu6oEWmkqbDrSz30YExfGE+n1n44MVHa8tSs0l
TkkHwTSIEtgPNhQ50LUxsHbKIKCACFjuQlrkGKDTF7P62+vbOM+ewMB2wLsHFd0Q41yOsnFLBjou
8LVL6ciKeiQ3e5D5XaTGH88x615HuNlxtngyDP4HIyfxFgfeEzx7w4r2qArSL89isUqqdV8rYDVo
eKCFzmvSPC0XuplPK7Dl1zcc56KYpfF5/AyW/7nxasrM/3Kjk2CwNcNaaeC1gzW9cSnRHhOTUsRz
fSpn4tcSKg5Uddmd7HoDT22Q9jZCHHQryqbt5azCGZcJLuh8UYlIjv9TelDG5BbvEJ0YF53wQ1jh
FQ9Y1Jn2VKwBAPE/XuKcQ7Yhpmxq/28Xv1mwE6geOKqH1DuxjHKJEZCtINiIQ5dPFJx96PNHSRs3
bvpA31zxYuAtGGMxLzqXlY8gkiMI6H/q9cPYtg5Q1Xv1Zzc1+XBeSJZbF3pAMsjaEVw/gsHmBWla
rJ7YmqV2dXdckgs4Hz81ExL+W91xM7knfCK6FoFeFln9LzYMnDVHpHYAoxGz2aZxnFzUqZ3Gv1LE
W73/eQu8B1g18AZrMkAq3o8nAK3z4S1oNYPkB8Vnog7SZlvaCGsyghlDNv7Z79CebHDhi4ctoHRO
zSuagcxD3y/W9EdnOZSDBdZkrikKyEDeSS3Zj06UPDloEpczT/vRsRUHAh8ReEvRBVomcIk/1Ffi
6YSCCAtVKBREN/uROJIpyEYy73PkLxH3AlJRT988uI6/2d4/uLVg+4fJPSU8NHDvefGep/dYnu56
0e1/D6s5yUvmdPizUtojJNoMOlUTQX+6AUNJn8GWCnTCIK206gtOHTA9bcSVGu4/Z85Eo59pRMuB
VE5vts8IVX5oBdMMv8XqGEgExTAPuJjMPZc86cD+YnkMEbdf95dwBOQtzsnlcleLs9bZf+PtaBWY
mtZWJ4c1zbCxz13D2d/R5jo8Gjl4KXk0x8N6+PDTQ7QVCg4k3LhxGswppeuPhUJCMQEav7/BfHiQ
CI/3+06bTvz1X/XMzmusqTWHLB9UZlqdEWXBHv2ujHu5dLJu4R61p8rdgnpeZ9YqP0a0KrSuoEql
AMlR/OuqFpPimnsRLdPsku4W0zECMUmrigW9JSiX2cB4F6/2aknWxAdCGb/h/yZ7bRKHvaLoD6n5
m09p2jAFiceYvXkWnx9BJoH4UAwAdxg7oQIPuuGnZRUW/150IjOYkJjfwGn87krlZOkWGMzPch4J
P+TS5WBJeF9DGlkgnbDllZWuxqDPbtyd7rkuCc3X8505DJScsCpUQHkZw45XIoMXpAHghdPNPR7g
PPWrHfjEPAT5n0rDsyBu6OGXc1AOhrwzjxmrgmjUAz0S3Qf9fO9LgzV7h1nhPwFNQdu1xutYe0IR
rmcKzwGKOwUmfry3FdKG+NaB5rE73BZD9yq3M4GaXa9ZXB0p50V3cUqcDpYsr5Qx/XnKm6AwBDc4
pvWIL3PGLlMILoVy8uj5O9vhDQR/+c9Wm1Bnho4D5m8y7P3WL5Uxh16jsZ49r0Hb1S2wK78y4KXN
4J8hviBib5bo7ZahjLmRZ1fjBOM87JiLC3STGEqAsQOYSfXPj0KAuEEJZF8qmh8SS5s/EV2cAL6Y
eglgTNh2LJPi5a6Eln3i/UX7NZfTXheAsF/0nQe6PfP6GdpZDZjO1OvrPFt3f7giqj+Di/k2ccEq
LqJVQHhNwFDH1HFnK+BhwX6D9CZwGRPphxun4QQOjRfTT8j9XEZga8n7ArZ4LyoenH+OSsw/GIMF
q6aKNmxdFuTBiGXiqSJttbmrf2GybkoQr26viOi3d+F61q0csROGApeHASjj5t1W+GEmpBHReEIR
Tyi904bt/3svTf4jTg9KKK3/1j/itUb1NHidUtboL4rp8xZGcDaqjjtF4/sP7TcKsWPDQ97Kikw/
RiTz1GMbYqJptw9j8ByJInwSw6f8AvMYXithd7AbDFsKiKMCmZrPt0vzWpzZLr/WJlrtqUYYXY/j
3pQo2OQVOzLiLzEAgPmGGLX6gMHBETm/9Eh8+eUlC5YiA8sibOOnyfl5asjArZA2IFVeaJHO9cuq
/dMI6DprvwkrDOTq4RWrpwkdqac6BPKTyKbVW1sslyyMLyhdSJKW1uHSnBSHslcendpLMTMYm9wp
AlrW/3JEfW7dc16FvGu0GAKuIMkDLccIEfXKXdmORm9nXl/zLGqbGGBPmWdRtGL++pKjHGRUJc4A
dluvZkquINqOS5UsYm7/wx0wDJftUaoSAd2oxqDeqmJoueK1cHWzc9Xd8t2xJnIarR1hed1KZ9OH
wcpj4Zsf4u5svt7psjmKN+pH8bePis4Yp9l+FJxx00fL9+9mkZBOLQLYt2xB62kB8WUubw1PXwsC
isKUbgQD2gjuxvaNmA2ZCOMCg7PjJgiEUjeDLsEVdC3ptoprhpMR2E78JiqVoq3ysT4H3QRGd2HR
BUmgrdHhsMJQ14z1aVGbcPWybbUkvL4F3AGvTKcbTTA3osXXg1Z3MWUGh6OAJWICOlTmTC0oqhKE
LlkuNi8CYIaVscUFp6sFEiQKKbhnri00X9ORiQm0a4kcFmAbsAAzxIoUMxpvLVZvPt/7GGQWhdzd
vminDx1/zMrRQgGWTWSEz+jQN+u3aE53jkQiVjAaqx2BaJIuP2GR3A4Qxh+4erIRd3lO+Em0lgxc
yOOYJV7vqq1Lhy9/Mm5nlKeImVhQUvLEE0x1YDSbueLl9LnMpV9Dd+7uJ5bjA5fssV2aKVX5QZRw
qR4uQevmHu2SBu//EMEqWoR9bG5+poSMr6N7GCsx3R0v4o2/SjdYKktvLLxvyaxViJqeK8zpqXtv
6Wh3Ql7EqOEXy9V6ieH3On7rQ3dHrs2TTIlkrQUivDz1DB9MgOl9Qlkdj6uv1hu26kf7dKlkDIxo
C46nVIIi66TPCTKk64znZJMvJ0x/CJCj0nZrmXlZdwBUzb4o92xAiL012z7GmGA/eY/SHbHbMedF
IO9sgQQr/6B978MQE1MolTIOGJVDrOzRzC75nRriMZDMRNXjAQoajpdWgeVFbl2Ik7ve6jSH9WUh
LyNQVt3iCQRngNSwAecd8IjhMUDvJGwnTnJ0+tpFE1RJ7zL+1seO3UnIeihPs3c4ORKL0SSvbwiX
pyIAEA26SwOmBCrwjh0YkN+E3r8wvRonxBiYwjnntGuClOEcHnVFzQPs0U2eWYyr2y8FrxQksfLq
LBMBetdvnNKbD4IQORdZxIAhVEsmG1Q4U9+RQ9w8L9fUoKc3i+O+um+JNYMo0KCLRedsJa3+dm4G
F/nEOPwfmyivRReMeJWBT1JwRcL2DvVpK7wU5JGbzQDVRo5h8iFozJP7KRgPLu3mh/w6o5Uw5pZC
ObzXuvCVJBsM2FVLCnCHKr7qwplRiKmZWbjkSs0CIvaBJhk/XfoqrOrJl9wLOgqtLzDd2N5m3yPk
G3XMDTfZE9CbC9YnbayR9PnJMB7MhP3rAxZBeXli/Ng+asQQH9L9WSZjCPSJJfiECi/u1khyjRNF
2oFKEPW6waf3KcEI0W9MyMXR55RJyLYCtVapra1MXdvBdlw1w2cPPBb7GRCp6J1llxtGtkzdUvhi
HjMqHrTrFBHqGAbo4LI474lgo2BhgiXuVtDJlVO67WOMe3UsEHecgA6TNy0vclgFcrXQoQMnFrbL
NWfuFxQlkdHwbesgREHuOFQmlLIbW2t59FJ73bmEFhJ9DpzCRxyO2veNqg3ENgNtF4gi41xodrHV
0WrVbgdZffmIvEXZfDXd4UGkKVptFSq2U/i1WvbJ8qJu1WanZbIMMd7CtGs15xlJ7zJRDilOAAdL
6osfET/Nqgy/DNTt8eOW/i/D0/lmEkUmhT9bk1kBpCjbuTXxM3Lae3qs835lW1kI9X/jgxLRNw/g
3iaNLncc7VoHeP2hdiCLd+YHkuQc2FWSNgNY63tOgBcQflBS4rXqHh5Mk6dDsveDgttwk/6g3+1i
0xUTKae967O+ELqLraTTUjUMUe8NJLqUoSK+rQSTGIaEvo3jVB0JAF6NptQTUgyYeT/qrLU/qsQE
O/85kVr8FLblI4xGtvZVphKOhq/00M4DIQSSwN/dKj/BvRGGZuq234vBBFOXOLKQo4t19WmHfSa6
bnHvAk5yiyXVKy/p5VKbj/IIK0rQDffHOVEYApP1sk7GTxWCaVYleE2kdnr6D7NVXNh7V+LmDUCN
m2eTN68w3RV5ftRbNJy/jZoMeqGzwRaKjrjb2dVPlhTYeqRV9oaAJ5LF1dbf+aQUhwUmmASxdXxj
Pd09gE8HIWOOD83vmYVJszZUTDnXbQikxWlQpf9npWK+RkRPVHw5T8ixXL53C/8hMi3I81G+1X4w
QahJ0ILfpOc7r6QBFvUD8Xgq22j5xMWyuoN+qqnMVrL+MvRltNNgS70KntvI7SW+nPxcb9PlUYYE
EZBI4z08DcuCYHnBEygaK+ZCb79ipW3bbVWSX+JF74WybVZ4FT5aDafjTXQ4epfpQfB8TglK8VHn
H4knz+HRusSOb22KQ1+4Py6Qx4WmjmP4ltPKZrdo9rHmFRNz1r2Gd9QuW7MMkwlURg+lm+Gi2vfV
PqQAd5XaUve5/p7r+7jk1CSYDrTvUjGr51ZEY3i0HdnI509uRbtMYm9/Olh/U8oZFlA/lCqNRmBN
h3RnfvdVkzt9jKBoXzEsnqy6S1L4yx28j82qIAaVo5WYHg1LBOAiJdOSWAaxHsCtWbMJA+7o2LwX
CV/e9oepvcT20fbhL1P3AqkeDamyOQl9Z+qupzagiwaWY6wfa8Lv3vvJQq5Ht14ObqyG+gHzfe4z
+DighTWR5BzCLHhD6wnCpirwaQm+wscGzxfBaYxmzh9Y8ReCNxuK2HenSBpAQgP2jKp8+VFXjV+n
mh4KyaABDGXJ1Clj+AoLP0cYlPdS7JjtHnWnw2Wl15axRihicKD90Hxqca0uhqf2pjASowAUm+hr
mUmjiBO4VEr2BqOCiuErwUIlnMH+rhVCQJoYmfUmkEriiYepr+u4V1AuDwVCXeDnXg00w0/i0Yyv
rviUO7DVPPJ3adnmFLsj2ozB98vQuWkdBC/EVv2nDSZcZoTERoUR2lwvKmKgvXuFQe0su2Uem1kK
rn48P6ykfh34aGJyMTsymeA2TVthsf8GzU1owlmw0x8IG0MjuPGJYDVu7D2fu8LpryfUy8jgsC7a
SWouuJJdZPzTDBc7HjDBD0p0H/1mi2/vdrJ3V7gn0pBxagx2lMhKGJS8DsccUw5dq5sOoGB9zfYE
KheIdHRpzQ/EFstzUqPUaSdSC0tRu5QPr/xEGCsLH/JhlkT3hSvUGETSZp9Mo7fWPU09ZDpaQP22
M/F7NMBQAKI6egRjUjMy492aP2qxHOKkNSvQSTBRSGPZ5fbFaLFqzPhbCkQgTW3oAeD5U55vQOu3
IiwSaXJZ5yomcx7kx8hNjRuR653+hGUcpQuSzmQlTuYsyfYNDgs3vYxdUVk/ojRmy6E3Jp1PSwVJ
Y3jX6qBjaiaUm6pI92tbywL5alqkqY5DF/ofm4gStWh1xMFWC4vdZY/clrhtlZ+o8anQOMJ1Ql+o
LfzNK4ZID0mqx2WLj1m/fU5rCW6KxGywDz/0Lj9fVKQWZwGbmisREJDN/Uh2gqO9HZicsyIt11vi
2EmXVDYXrwale1z7udZ90yQrvluDlcGQq4pTSg9y7dpI7nxjGDnXMtDDYj9cjvPPJ2/0nS7hoDpn
XFG8xusrAhnjsyo4Uy1Kq69YuiWm8llHJ+bXVJqpUwPQk0YHQ75nx5ShhuXg6J+Bbo77qG4cHpDh
EZC+uzR7omE+3wbjxJQKmj0tjpXXrfJdlU2kCx1NHjCmOEiETObESEYgRh1Tx+dRp647PCokFXLa
2W2xBh0fy1Uw2t5CXCmC/u3lalRCqK8n6D67qlLMucZPEJ4pCEClWSIkvR1V1KXBykKp6wYFvU8G
W+HAhBefOd+0YTLTRG1ctndhhtsgExCcdv/M2bsoX8Nl0MdxS3/rXpMJUxb9txF7T6QcWf9fqCgk
qb74ABhGphfPeiGLGfJjtM8jckPQZk0wWKokIhVoxjHnn6kBbYhc9YJI8NNdMKkGZN8pGUmqMjMk
hy56zS7Gl0kp2n2HYvbQu51GCRd5WFcjFJeLfsmCd4cQb+0wMg6Qf8A8vCto5/+eDzdBjfZCL9a4
+e2GdJKXznTdin0xqWV4jhzCZCcirQaFqzbSAB1oFE8sEnZSp+aPJ2Z7AOtDldgZgbShHN8mpiJ8
MtfyDRW0yWArSEeb2+kTnrOZCT9uIrMwuEdM2D/ILGO/jOg0v9s5tdtnxMpcuCry+vc6qWeRwN0L
BZ15Epe5vHpfGWfYTAa0duOslnSdCmezZPlBK25id9omZea9fjQzcV2c98Hzrssz7aub2YfBJH+n
x9Vv5gW5ikmzXGcGbk9Lg1WtVfi3VhYy5QrnZTs9+A/jmk/12JZr3uPBUDCWt3tnRXKqIOsGj/U9
va8f8X3qKCiygvu3VLeWO5lVh90qeiA4FeyOkA1suYP++Wo94YUfMmdhRQqAywDDEaMEnds7z3gY
DHAiU4vJxrTUPT7kEoyRVH/ucSgwEFUp+9/48Vz4FuxHqu+Rxr0FOP7iPVAtjTTRCijfl8519jGU
Ae11E0pypjvHx4tiazbpoOytOUWBDrsflroFPUoTuP55SbW6AQdqJrlx9MZH3vub6zHETlnr508h
ObcQMHYOXcBPdKrCkVy/BiLaBSPk97b2rJmv8BjzDGuZIaphT4PVS+sTdwjaXt2VIdsLjC7C/Lbf
ExvK2DqLsGwNvpggRxyHiuznir0YZ6vZC/3BUrHtLU8/YmAjIFR8iv2pEtvb7SR53pxQ9qwU1jo+
x2EYyF9iR9Ub0rZpL9riaZHp5zJRCvSaAxIX7+7LPtmgJh+oqFYJ2YdK8Shw5/tvNfR15u31Wr+l
LwgEiSnEKqlr43fe9BB/tySbKjuGWk0oP/qIZ+VDHQaxSGbs+rIJS0uvgvvzVSqBU3fr5E0eU6Q2
l//feloiIjwMlEk8MVQZ6BaHt7mAyZIq4jJA0YymJrUuoReDlzRK/Njc25DPkTkRBzfm1J5yTddI
jBbAEWZi77V1u3McBCZFzKS2b9ATV8IK533hoVCWx0U3OI0Go0rJHUzy5auOo9ol+y8lEqqeh0jN
q7tbVlJD1IEyX7w3IlQIVHv6aK2IjNtl2Z5x8HXLTQoYv8YHYM6kfvPwFesGfLL0gbvvjNezlwwc
Ah0UIyBF/jLHeMs9TXYaZIQzC6BcLL04kzUXlUgfGEMir78JDnPivMghEWWxnKZLsJBm9UoVVyNF
DhkA4/P7y/lKkCzCB7We6ucyFTeMFq0Ud3uOL22PPv9+xRI18l3uVy8Y0DOriARhjdg5sFzwbbRF
938RSza3xVXX2imUC7R39D5wv6mRSdr07DPT2zO8BNb5zswu+ookh7o2l+fc1GynVJWwMVbzfq0R
iazHJyi6gdSV6YIdkRsTT/Fe/jMUBQ61HxfO6KziHuUvbHn6mEz1ZOaF6bgtJHFUHog6BkTQC0e8
yHECVSH8H1Zlalhe0aqmncG6V8klJdACcDLTcX4JxbMThWhMm7In3gzZ61Zwi/uk+uL+P4DAbQ4x
K67DZOpVhu2OJjxJieyvsZ+VZbc7+8QbooPACz31U99ZmtGdiHvT5BxOkML9Pl9P0kIGHRXTRR2P
GMExpNkrBS8B3xunw/YkuibLVxlefIn57mFfFlFIGba4jEC8ChU17fjtA+bP2Jdh9FYsCEU5fXb4
dHWQjNhh+85lt7/belpsumGQ2ouFc5zJYqCc465Uo/JU7acZBTXRYc877hDl6mYhE1A+KN9VtGST
012Et19bC5AhNO6A2O7eeuHK/svNePZX4XH30pjZKG9lsGc2YuKXxK0dlZa0nkga7WcFDsvcmuha
ZG1xuC4eIjmo8XDuyyBohbZGmEkpmb3jqxMZnT8Q95/s5OsQYhBkiQI1gwkUgHdf9bF0I4e5ZNLY
osSpXyyoiTPcARNPa7o5fYdOXlEC2HgT9pGphc+3cSZsVqZuD9nH4RTEVCKT311EUm1N8Nf9aOBG
jDWVMEQRFU6STPKQUm99ClXqNDdSogmejgyQcIVVQ9047CsOdwjkhxdrH0614mrtBFFrdxsLL9GY
1GVrM8lG7IBESwaPZJba+MrHPqwc7bsi7LbNZjiwZGdHKFtfkupLB6enMpAxW418zlJ0aDhRS6LJ
d9OE0zTDMyWNRmKJt2fu9L/ECoh7Y5bjMKRZ4fr5YQjh2DyH1ErXB8cmIMjkh+oSdSsZcsFR34H6
Rr6wlHgUHWTTRiU0QyHgOhK9p+Kin2qBZub5r0njKuFFbFI1r1p+n0GtvzQzCY3saQVL+UoHpMvv
Nn3TJDKvGtYQQyxnBwuwAOHiTACSQbxj9R54MIgfHpQIN1sJmDvzvJwIuWbAy5YGa668qtDIKjhe
vRTB+C+7rc9kFCmhqNmvlOWSt39LMIup4lfY9EydWFkgshGPHM9TKNa+N1OCxHGILloHl7yfX2lY
NLMhSb6tPbHlUKXiGAkEamt8JHa8FV4StBwzoS5O7/PCu5w28k//1+zV0xWr+6373+lnGp++oI1+
ZpYlS0b9zoLE5xbUVDjifpoBpIskbAgXOzYLiV+o36aB8NSqdaMyf8GyQ0SI7qjEamIglRpO4nkk
vxCkLmGIM2S+7JTtj+80hjmSg3Zcl578sze/tLtd4oCgAIMQOyn7LjNR873rCYMrE8DnqDKVob1h
HdbqRfC2gob3hykBsd12bimLiddsyjeeHkYC67qUHML1xYnxf6HKSOaowbPVFnQJk6XXqRreplpf
FTEzRB/FE0mhI5U+IzTxcs83wlpfLV51taSIYCf1htr2XBenHqLIa1GoLy1T7rBJSNaR0XacgBfd
17yOQSNHIG3PTEfGTTXov3/94CwMiMWX9lGqnLQgBfECon+RI1cNcldoNknZlM1e4vIAFh4M6BOA
WSXIFmdz8qIuOsEa53vRiHs96WbHo2tkxyiJTBikH+lb3+/Dz/ywkjtcYlvjHLQnNTWLeBBo3Wmj
vTY7gjgJVJ1xSjIpMTvJdFUygWCtRadaZGqCoZ0dDaumJs78CoxQx5hP5IgVWw8csne+nslxrAty
WiawW1cz4uKsMjdDBZjiWz6TvU78kKhqJ04heWBGNAf/NJFuXdMI4mgr2pDhrNktvh7gupUPgkRL
hZaQ1YBa0/HFmBcEdTZY7/9/DDHh2yGCnLldaAEvGWF3FJImQwSj4PJ1dSGJFwts3EBjRNmG5ysP
X7OT4v3eFi525bB+FcCIoGsI0Xr00uhFGrAxjenXhjrgA7F0oBSCBksWOwigp2jl+AjMG/tbwzH6
0+ZDX6qpxhqQsUMXTf2dsk++EIljwRd+ptjWKav5W1q4fnSW/SlsJ2LY2XEvO7exdueevoGJp9XE
34rCbPE85lDAO0vb8nEnfmYVTHxpGPkpfsKPrJ7ZZ9Lv6ZBqdxzkD9/ACOKTm6jlzLeGeSpgUfAp
nQ5aXIdUgBbVxKlU/+E4Y96Ato9mtcNaMNIDhA6eA5nQXYjpEwVhsDIzkJqxm9sYBF7VNta+/cEl
4NnctFzMW4EesbXmT7rRDrkSeRDuufh9ZqXGzvlfVValin7qG1cupoXvOWxDn+hqIlhFMmqc7//1
1xYqiGMMiPD1aGYYqQx7CnR1Rc+DdWcBtpJ06KKYS59AGPzl+hVHUAkSELZsZtct1guckBcB2KOz
S3WxtBSOZlzeFAWeN9/si6OQ3Q0niQgIOgvghxUTgDbJavTB8wyhl9GQjHLUsm+WYIo9rrKCaFGs
AVv3ySKZw9lqXMK3GVONVnfECdpO5Czle+HJoeBGOqFsSfSC1vBptib/CdB6vJ+D8KJQQBqMaFLv
g6i9ZTQMtPZkdXyWGSTQ/fTXq+hEmi1MvHPkd31YqjFOl1Uow5ok5LoPdGCJHfeYzqUfkoRZ3Arp
1e+ABqFl8p2IJ80cz0q4XTyGgwAAPc9bpvzUHcYuA7YOv6fvIU9+jnt2lresLc6fM+pcEX6HokQ6
PDXW0RGAHqQlOdOjrZHAQPibuL+tI0Wmgr475huVgK5R1K+PlN61dqc7Lni/wBojLhRVj5Sd9IQJ
vRngUMjGxdJMgOAxuCRAlWWKiJxwR/ICFuRPHwViJwJE7k4n52KIBEm5xZwovyCNgswbShACmSul
IrCkFzvLFH9WvtB1MSSE0JwGeKKmidkh6n22SIuYpnKPIzJkDfPxQ6HNqeV5zwOXEVzv02FcwnGZ
yCFdbEtkWOKJP+vWfAAvnyMiqgLJ3kFBGqe+to6hStANP/sBZ6pH/s7YwheCrAuh6ddac7bISUam
h5qQJMXOjtKVCqClNrVrbeGz5hE4Q7L5eGBwZbhfZXxzwWIP05P0Yd5MHix9ded3gNdWazC4Rpx7
7TfQ79eVjjOSMGO4MKdrhlQ8EtyIJ/4mtlUa1cN0yGWxIvuCBzz+mA27YI9qVBcsX8yeS0NHwSiV
4HqJ8WijM0wL13RxwKmgWJh+dNLAFB2qVtJghAqNqFh7XqrhVzAMvF8dPNCdBpmVdb8PazcEJ9Jn
PSVPc2UAsunyPP4yczZpU0abGN5BB3rz2jouSDxSPD69kmTHlRbin5A8NVmrKxrVZLmZ+EOZrPIa
TFUsjEprRBVtluDVwxr6IGnfgP9gUE7s8qlsu2cbkv5pGPSkIYF20w1Cn26pcPaipIFqyhFJdjZC
NUc8OLvNQWJvvZ2k4Em6CMj+htnIDoKAd0dxwdIC1/QuabZtbUZEADHRfyBWytEmenIm3jcjsEw1
+oNfHCPOZSZA+J39GICpAg+xD3Yc2plEA8Bcab2UYM80xYvMfGW2JAaabXmxI/o1Pa2/3Qu8K0QG
oa9QQf6fHq9cpZh2/wcdvSkYh2XSEp1O6bPfVteEwC/OkSL4jS+seQU84QMuh3bd9KjajN+kfhsU
QPFoV8lXtes1tbZ9DjwCHvToTwIW/79NH5BLt4ikeE5vD4ZV9LupXObVxaWLE7pJGG8QPLgskbbc
3VLvHsUVfnZz07kl8Pa88EXDkGCB5c6DbASneq87cmCtbxCiozWQ12Oi2JfbpuYREQ17bgXELvR/
I7fU5pDot4i3VYNthf0kkeaQou11TBrmKc2PN7oXGEModOdtf9vm+KN8fVZKQfN5jvZSnN15e2fs
uR9jeoNwqgiXzLylcFWY1RL0FZPBNJKbd7hwHImoT7vkdj3aT/JmBFc+FZFohB/BFRpgGQF8c+Z6
EilLXN5xPaLwUbN2isUISp71OBL9cRbL7yXPoRnMJGx2GGQvytEw7wgWWkqajQ7s/u78GBjbmTsx
8iLZoEevW1II+UqjnxPn4rtdu4P/nm4O3JL1QyphpkXHFfw/pfwlfpuAj0FHSs6B6+ZGc31R/di7
SIS//aMbjz0XLSnQ8bbXdaURjXwfEFEM3C/6kvcB4f0AH+Dg4PA237giGSXHF3+A6PhPUz7DYTDZ
MuJ54mZEKYO25mWutfpr5UbN63Y+kjTlHbLyHu1OWGR+CJF3CHBn4W5R7dZIwAiNrg3ni5rE5f5f
t6jC8l/P+d7k64N93vZEAjL80kjuwo6g/0zMPjFpYWwh0z72gdBT1zVlhYG/HgmDVrh2kQ45Zdh+
Uvxt/MiNgyiGkmP51Az0oI7CQ4WBRATqrsIbexw7ohqb07XfhNoIn09jNTK5Wst7IR7ZTMOotd/E
ROI3QKiBcpwpzuo9EfV26Qlaq1G9oy8C7CLC/XWW4+2FnC8v39KozisZAfdIWabYC3ZHoK5J2r+h
y470YCQwPf4Ye8YI422yljoejzg1zOPe7rGdhb0reA49bJDJwfLnoLoy/GVLdsImaHownwB8BT8N
uBW+pexdJrHoNm3w2fAS2BBChwDvI+QNWCGLmd6AbYJ0rAL25yFBXVj1nAjIbG+iEcGEh4euUoj6
OshGoSNju4DyXFSgQHACqUFoQFSeqXgK+c0hsiHA7DBIH4BwVjV4kAP+L65bTFWl+N8PHAzs4KSK
0ODjzD9SfTd2aNJv/Cyk+7eIeo1FmyzwZerj5INGhrVRs5oJy1zQux0mn/xg51Na1B7a+FmNCVd1
uFi2mqlo8um3KIIJHUTnXLgkoDxf/K5C5ewvlxGBJYBDjJNhZTOKnvBok0IQd6F44FoK6ZtCjMnl
UbN/SD2cTOzcwuhgG2+UeOd66B07ARb6Lhgo91+Hq7sWdHiwvLeEDavLUfxRjaI0LeZYJeE+SoTH
Lf/qUvW+oyA0OEHBtbaJ1fGHIGGNWZvdj3EbOv03zqFJ5q69y2YL8meMTmYkE5cWUKI80aa5OuCr
kpRSMwhRRmAPoPumZLibR2El2dY6rNyutOM/UMw20axmUqa1YnGJ1fSozpa0OK7kv+ynANRh1KRn
RXjEuM0OPnvl8xSa/eot4dOuwRf1NqjEhnOkO9puIVumGoFmssJvylOmcwVv/8IIzyseL2/atpce
g1f09OLTwbsStLR4qEi1Xb9XsARBothHlCWR4YG18O4YqL1qloOYc/7lMQU/fLDWKBGAmwXWGvoU
YZWhoPSncU5e7sKWtYzQycgXFs7L4MF8wVnxCxJlm/8qEx5l17ASB/d16BF1RLY85gWlnQsZ0P3G
SqjGNDKZvaMiOIp7LLjVezAqLmA+1Xfba+CuvR9fQ+TfdDjoxdGo0TYFJo6frGRfKOIeG8U0+gRq
9SrKH0F9was4Dv5y1luxyJcNXxqQZjVEwPJhF5IIUWFQsa69ZA9iGkmv3fgiYmjWmNrJHaJjXlGV
qV251SMSG1I/BC3u7j+U53gBhAiN6rwsH9cdYdzFBkUqa3HOBpdUsxTwilcY++wzbovB4WWZwooO
HVc3nBrulbtzJd83niixx9zzLJH2muwkliSoWDDrFH85NiI7mQh51kPCFoC0W/0mCSKSuV228bqe
wSX0Mmc4tRCBprsOL+xytqSGia/oLlRrMaHIjQXn1aXa2NPcgS6WbV2TLr7wjNZBePiOx+NXAmov
iVIzfW3Vjzm7IahNNY8CWZAzpOFH3CthqGVc1+xL4cfmZ4EjznCLT0N3C4U73N+g3X43KkbspYLT
X0IAMxU4aOEJ+0UkPOH9PiSAS7D3XQh5Hb/xgC8Nrz5DEExgFg/T7tmq1RHIgpBvOEjGGc3co/zI
T7Qb7/+XmWnY3Zrxu2bAfke9ieBH3VO8hBEYa+xiu3BuUFc2yTugzb1CBAfCdJj6TCdf8Pqiui4y
JyGCyN6ewHvntUh/ars5J57rtbuL8wS+cLXM+TH/DabUK5N8tm3DJzEZk7ZQ9AzV9BHTHDSlnwjy
PkXwk08Eo65iZML7inWs7YlZRMRS5k8KbilX70HGFhxz6dN16TtdMX0oin9Fum9G7Ff0QUN4qEkf
Rzivr9nwVg1rUfwRcEupImAOBX8v5GMTTsEkn0hxNjuUkMXRxZM+s17wPh4SMIEHtQ2Fyjd4YgrM
O9YjL8ycWOwu33jX3efDiNIB/Yll0PfxOkl4BRYF67SMxcFAFyrk75Z2KVaYJ8FscUTDA2Z/CiSM
MO4TOBVt4lO3F3pFvAlwgyXoxUncjofQ4JWQJcySIlo8vlwv4YWHXYk/qa5NUvpfMilmcvkq25cY
PXfonbIJjU5MWsUesPM9BrfBAkG3m/Qqmisq+TY/5QYREiheNPV+/6iLoDHkApnNtN8u+3AWJr0N
rCAnDsroILTCv+V/WVr9zGLTST0IQbU5X1uiQj8x3VpmA0wWPEN5CoSEx251stc2V4JkeQod0nIh
r/dIlOkYbspRKV+tcPCSBhT0hbI/+yB+YfEtnHJZOYMlv/Ndc1xQ3TYpVOFrhZhNYPRXvXg0zeYV
L7fcryTBpWak7pLtO1Cc/nzoFafG8PXc0b3kmBOgTYKkNO8FYbKmbetzqxIOt+m1+tADcm3btujI
ftuW7ANYfYvWcnVmXR4/hGPa2ayQWghQnG17KRbhDOb3lchjsbGiedrfXynmPafO1zyu4T4Ir67j
fSIRqtykEnhn9gAEQM7Sfw4vz8XJr1T+qNUjZOklXNZg4MIhn+Wf2gr7P1phj5MuYhMLpyKw4P1n
RsIKGVcWGG4IWi/D354QyOjO9U/5OorAvsaijg99T7HeI/8w7I565imrfxofkyIt8HkHXUlyOVrA
TPYwJ+QTWXYjZK/LrR9wUtPf7jY5addRK3YJkVeQmS+8TARUYNNKay2aP+FV4yp7c6HROtKUcYMj
PqIwRm3UL3/9S7uTdTGJSaNe07hksI2qFcfYn9AhTqX8IgLrmLd8D8PJPLzZqz+2WsIX/YN/rs3c
6jd3eryAHsV6Qd+zo8qwV28cmUfP/ykjb7Llxw/sv1SF4FNTB2Mm8L106EsNFdsNPPYWBOhThr2E
CcH4dqduAQhWAfoQ3MhrzHdCAQcvBZdxNvBd3SFkgBD2rDVuOAiKpaea0q744mHDOWJSlKLVrjya
Rcjv1aptbJ59HFBAPKAKTL1S/AAgnBesfNUl/gIZGW8TBnjBNUeA3tq3gm7QjpUeNyhvJPF3L89y
WwrCsKVbQPSGSb8AkMqEL/Kzxo0B0HGjtYSYX11i4Po7mQI37fi+HuF12e05C3UNZ38Ho7gMOF8p
/C8C2YuIiIzsquxvUyPEm8W95icvA+X1FWbvg5s7ekBZkePFhE9C00zzetMJvp/XbhGprGDUTMno
396Vd9zUXhCb9x4O+UQW7RNcWL3eriPghRdOz/97AKJeH/rrmeMmHRtShkqMWxl2JS139bdz6wn3
vwSRN0w9jUwrUfPnV78kwaRd+J/CuPU9clisadkbOICE41LE5+crn0GxIf+G7iZw53NAYerCu/4C
rikZIFsLDUYy48ZaZq5SSPl5OV/ZiyjrGX5UzT5eYU2ZfwJA0GcLKZLD+r7QfTWWSJhmcn9aj22M
o20yz7coZ4og9plH7l+mk6qzDavniwSSIdwiL+k0HWYwRmhTaJqYW3cODvTIiyPGWo9sF8o7RkZe
zRewWdxgZx1nuajTvOq7e6yuAgxiJaVCW0NfdlqPllN69BUcGdFdBRB4kCIlXdCvoysSfNGVI5Q0
HvCWI91JXIZVz4yuerZCiuUPMO4GhS02jYFSm3Zdg3v3WPH2bmJn4i9L5Xoqrn9Cl7Qunvf3jK3S
MBJQceTztTAiSc5PD1ThEgRHueLMLdY2WgV8kMbsttUTFy9+snDMUJS99+eWJRihmYZM8jb1dcZ2
GN9YsLOzIveA746jItd4ahaLyxAe0yscEEuyrLaFhBw+Thu1y10L8lhY3WeOW5AIonL5Kq28n2XU
JHnOcQUX756lbvogazzrMcOPZ5X00/GkFLnqGORM3kep7NifyvMPSZQyBJWJN1WuqOmHxEfKjyIc
NRJnUxg9wMytY/yDXXV/bW6fx59eeRS1vONqXwZ0aYhDQf1jNYkgld1RDkzBhZnD6+0fx5LiSUqg
EE5lRvYqvktms+vLCt0umUWCqcU3H2LRGfUuGgL85G7msFJc4XSpVz4nEGE0n6XYX6yzqGD/H8Un
3bTD3FDjuT3Nc/kIY1VyYZwTgOpAWAVUNiaziLxSYHHAmjXKZ6VFZH7q7mTYg3zXEhIj8eikGgDf
QblazxM9GJd30eKmXkymQgNnlOz+Puf3fcDKZaBgrFXThkm5MqJtDAiVfk1MJoQujkQNTjkkgvbt
glAa+arnmoh0M09Lc4Ubaeoev0sRb4CaU3de4hdE+26gLkEQGLWyeKqqM/IBBHi9pRHvLCesxJCF
v0h7CLn5hixBIL8QxUKyoyJiL3SsRE8wZlmJJhktlKREc2lpYjrJdBl01pvt3NS0gw3MmXTFsHbz
mGvfUtTYn2Q1fqvDfg4Egmgrt3szvNBumXcXwIr16AJMveGO36meLbdkKspEAuNOMMXpM2qd9eHL
5ITtATpiM7t93w2vs/ym9Fe1w0B5Lix98VRUM2/duZfel31qhViSGJk+fgXJmJslEHKeNKOulcqf
wHEhF1jqcuPk3bsBf7V7fwNBRxBj3KSphBoScrKHjnVoTgSByHKSNJsTqZ09p9+7oFS9hSbilJD6
v6erqZkKU1Rfzk2t19y9jg5hZUXoqbwqcQs2gXsKiyJuhMzm9az3RtRfySSbQ0gnNtllVyThO57D
9CZ9p/9FnZf3RjkXPAES+yhxO9XLcQDlAbEYc/H0080AtXVLR67BODWeDVgL2hxDD0CT3H2qfTuc
bmYNZj7zyXR9aqwLxa4r0DJJj6jAcPdqo7w9m37gDA/Sn+BlyrBx6wm4BkVDusq9Xa7M80tYDHrY
dnho5CIYEEVq7FtgYhxdKGbviiE6bLSG9CPKX2aekYUkNy/z1SOaathu7c8TAPfIZChnjtyGFX30
veDhy5xzMfBnIeBv9a7QOdDm9SANAIU185fPtRXqTu6fe1NnYXC6zqpPtAVtslLligNYRQJxEe3+
RZtasj4qpK6xt4JNG1iScR31AkuXcCb50egalfAITzoTDZsmOzOpzRmrcOoW/oR742TB0qZ0jeY2
6YEqzovUjGwvbqGb+4c67+DSfxNomPgKOJPtnhrFy/AiRoOJY8NzkCD+YX269elhWLoTkthhFDe0
nyDYuiq/2YMASSbe8FqL2LFJr7HGW0thW7hdHzGfhVT42XXylG8jzX8Si0DNvk3yEcs/IDRz1nG8
R5pKOaTkz9gjFvLIz72oBn0nYd7Z1Z6/n4RK/Pvyy7NlSJVagPbSHHc36VeQAmzMv/o78+ZDzmQg
MJaVuVEc9DQD9qZUHCMALWjCVU9DOBe7BV/lgWd1xgC2GmQ6kvQ68J4J8VAn71YqWjipAhtQRCRz
/OvwZGDcE+krwoW+HHtTXmMkXTAnddkFTLDHtPyZAY/J1qAkoFfVjOOrRhzoIphHY3ETnN2uT33n
KJgFviOPFKpWO2ScTlyo4iNaWIfevxDPnF+H44S7N4zozjVSvAi6wzovjhgM3LZzgCxWHXg0UxP/
fzCq52FVfWptvEFG0OvdnRnDwVql3fe2WUc/38cVkxaNJoqYqYYf2m0/g3LokzYRtzqB5Q/XIqJE
YjhupWAW0DNe8a2QHhgKGzwXWaBhFty5EfowSPRhJZM225EEHok9jhqPE7yiii2rVovGADfD7d+k
sFu/Qc7JW7gkqF/30PDPwEz9Z7MJ1b5vVFs38LlS7IWAZrQdcIaQCB67VNsaWuv4h/sY82IC2W+T
NcV08PTGZuy0pKuz7xm0A5Ty7Vf5GltxILch14+RMDL0lnA1l4R910Td+T1SUElz3RFm3hozADdp
8U4oAn3amqewyDELTXrL4QJzeADQBXEAxVTOZYDqsx6PmsXyAEF53hq4c/nuxgct9O3795v6pXaB
p8CiaaJT+/Q3g68PEDrr12JCVbv0SUFi8LZOxPLlZrumCWeGRUCunkFduLgjqCVidTFurMCCLtYZ
F4xrxW9ITXNRzOt3G6pTKt/JVxnBbHjQTCgdlV306W9L/m0ETyAAZ+5CdM+d8jnOLdVe8br+2zwk
xXZ7y+Pmo0Poycth1IR6dLbatQExOGBpCxZDRCNusDC0rMdgAb4gGZKUGqRiIaH0mFadmPiGx1Fk
Cus16rPlkqz9YnHO7/1ESXK2T1ZezCCcJLXaKgSmnDgtuucS7k9cdMBlYfTUWe/i3/wDrH+waV4L
7qR4oed/u9N0rugIfd8OaEuU5TmqO0DC7x3OhYeSpfRNa8sq6JP5vgeEgGzGe9f5LfhDpmwHblQK
taARo+0TTIGc1nVHT2wckuZI6eqgAJFr+7/UJFkE2i+11J9Uf1TZhHidDw9xUX4I+at42q4mUTcC
83/gSZrZ1CN141I1a4l30UjvCGdYFrxzwlNc60XQdu7iKifZRlCZSoNr9WfWqOa2MLPRtJ8B1EKO
l8Gs5J4r8FtvYmkwOzlj0N89fLT4V9CFG+DxRIV+UYCWytr6pABkjSddc/Wa8UqLUM2Ln8GdG+Aq
UEJtZUE30ys8mQlyi0SMEEJbUwvAzW4B6ysEWvlagZAYGdgFhSU2Z1PKVJ6tln6yU3P2mIj5ZnNk
kswO3keZheDNngmLc21ihu7PWmSPH+PlsrrUWJJLaxnNNOTpqUMNSRMJTqWiv1Of+BwlbGMgxEqN
IP+8QbyV7yE07T3HWzCYg8IUpffN4UgminteusxXRhIU7tg5DKRX8VKwbnrMMjPlMltwkJ88Qrf2
1EFc3y9DIrykLWY7nIjAXTS44wojFwu4+kLM31hGD7dTtabF8IDfQXovlI3d6pyWJytC6/9o94MQ
ASB5rqsrmQZS6fII8qUTVkAcefE4SNLNw66MCrb62V7nEQ1YzCOWZT4zRzzCJDQ5NZcxNg24Rhwo
gh7I2rFXPwesF7umQzxdaqH+gxgZiYlDsmV4t2tUm40E5kpyj1Xbmmy+xD9Ia8Et/LTcMjrjCpTu
U3LRWJ6tTIXZsbJm44U0F8RwfJXhL2fVsk5P6pUbH3o9PXOZl6tltJgD9/HqGLFkkB7D9wu5BAVU
QUGBJuHhFbix5ofgt1vvlnMT9/Hjp6dEx3JH/wHgPDHqzVXPS2Oqn0jC8FzGKcsxfemKFCPBQxhT
6hzsa3Ou4jP28upyxxEruXYtj6OUMPS45Xa+dXcL41SKFycZqJjQFcKUp9PiSq3tQXzRwoGhLHKE
DgGCYmxInqX5xwBkTQhBBrcuLFxXrVDbRVH8jwMm03RPjOccyhY2KjpPWegPdX0SsmCDRwA/2xEs
+njtzVgYbReUMvpHxIi8ygyr4f6a37pHmOvxK+Fb8djz9rW4xW05hd3PcnafpAxDl7RfHXtXzVaA
U3EGJMzLVohptZU6AvRYyTdsfBTEAa3kWNFWTlpjcCpqeXFPyH21/TVufKFHWzeA+jX3uZ1YxNt5
DvPxrbeltDYJIjKzhsMbXHRBi2q44GzVKP2/Se1CelUvO9HUW3smZNmfB3Dl7/TrzlyiFKua/CvO
Bm8lvqOAuxdfnq5B19Hp3h0lTT+ut+MIED0N1PGsDwqUEEFs1fSxDDEg/A5tyr6yRCZ7jLN3bHkA
m/s4Nafl+x+UHwWwoQ4ofrfJjlMMnI7R7G0YcfY5NzP/xe4BCnGFhzIJcE3fOXDS10sRmlmFlYlY
M3zpD8pxVY80D8nXPyw5qUsxghveoETBJ3KyeKvgjS/VWs1IXMUtG4IVlSqhL0FqivWGrb0w7Bxm
GO7Fas488bjpvBhJcNfUormXDT+c7Z737ajtbp2wGu1mTZkxYuesYFXtjzpQfnF0Mr9FjBzU/nE9
a62rW0VbaLtAQZTpQl362Gbnm7IAJ796bdhE/sgxl0uI3Rb50jGBXlQZtwhEiFJnt3JOpkKakBlw
UcfZgjV5A6Vnlb+WVJjl9dwa9MVz3FO2LMUOrzUirA28sPY7Z9QwPnAuZP8pFmnY7KOyChtOpCEg
pWxDbiBXnbg8nTtDOHRC6W+tJj/FOzacSR/t3X7341S/4YlZiLlkVNcmxt920c4QLcN4CaN874fl
yWKIalHd2qI6LT/Ob7G3h+m9VzWQMeO1RO75z81OKqC2U5Xbi4/Dd4YeR/mUXKba/skNF8HVWR4U
RW7ELRCdMffxGPyJDy8ZBchLFYVCMwdasp+7T+5ixmRL/rUXoZoBw/+5zaGRtZC/QIN2rwDuqH7Z
EUtTNfWpaorrzgyTnT/7sZz5VhUc5XDHRDuCtCkzAM9fV2vTZ8zKVK3hGGuLLu488416bqVhMp8M
lhBn9y0K77gEXbTz+GrCQ2eKIMJ90QPNoXA2DoU8SAyWPkUHHPJdvlZqUrCeoDgIVR3+XHLOac+L
ldhtx5UcE9qdlOKHTBjh8zvi2LLE8Xs6uHOAnxWMtFlSgn18zvE9RN9k+95Y4eoeUBoeZNyTywn8
FRhLiI02JdtWgSg5Y1P23BQ9JuF3Jaq2L7B5jXXPZSlNV5qyhi1gXq74MIpc8RUMPjo7/TjL3U5x
nxkDoFRKC99kOJ6068hvTmZZVRS+5UFZBQp00OC/YfV7SqtlUJaQzUGlzlcifzAvbpDORi2/Xlip
mQgjcUeOZk4BictoVAUo8TRhHTIqzcE2vTyl2fqs8b7kW0APf8vYBu62+Q2iJbHyQBhEsb7VpbR2
uSHoyyQ/ieadG/CFGKs/I5KS6J5U67TsmpozdaMwhVGJatTI1xP/vdWzSta6rH3JFGYrl9hwByty
vnw1r6uLs2mmoxHripTxGVj9IOSyz1Ed24aCui3tgsAHV3e2OLd/yBtR/fdfxOMRwj4MBEhI4KIO
8lToo4nbtiSij8/pf1UJFfgzBLlFqyNTqDc5dDtR9b5uDx8UX40vDBsQaZkn5oTVkkzN2E+wmdV5
A/PGuf9gjHARYaHMYwQYep0H6D+77MQfbSdw769mJx2Z/0US159etW+YmhJ9OQ6/zXkOuUL19ICG
ALbNwb6yLu5Hfn5kZIjjBoowB9g4NySEpZI0lP3EPjqCpL5sQ9M47fis3ZyqNvkmVfjzd68dtsfA
WDttoWizMnfGGCjF20Qw5vs0VXPnSa9QTFNpMY1W+8X4t+jeQFOipC34HahecEm9fkpYjfKMQW+f
ajHgcT3wRqy7ZmQ5rjC2Lp314/GyrcO04U7IObgAzDd+HPTRd2/KF0vF4Cu/BC9UjDxqt2UJ+h0w
I/bPtHJs6GuuttTLjRJwwdRJPLHKrBuJpppai6BIGcEYdK+DzDGiYyoaDvgfOO19m0ViQv+W9sgP
pMFx0tFMf+Yrd1VJ854y+JU1nP0w1qETGFrF6a/1E4/71rSA8+slJPuPnKZzjWm0RltpjHqTuhg0
o54L6dTacGcsXma9y3SQR9OZKdfsU6NS/Nkgdtxz0GNy41AyCRfJ6zWBZC8AhM+8Q9sBeiNkGrIt
mkq7GZseQRRJ7dL5FBvTcfGbDSbuyQEnHoAA2hfGB5JogxX9s7OPffbG0BjJhXpPwjryVPze9eEl
gw43RtV9/fQofQBSmHHZ8RcMbUKQHYTO51qHqxBOT+VfXr2a8KhNgc9+6rpuQLqI4OaKqa/mvqtk
ClpSdpHH509dcwYX7dBiCrkKND032vDgnLPiwmuiTr6uISNLq+9UOtof2RVGTJmF2ljtaWa6cBup
xqhrYgFCkaTCfB172pvUBjPrC7qsCeyyi9T43qW5q53ZNgK0Jk2e4BGtEm03Oaw/H+tNjigX/oQ2
/sPDOb/C+JYDnS1oIvZO6kiheaPjO/qPWvUC6v3Uecu1YgTT0iqJzy7qkGOgNkmlxxRf9eHF2SGl
KNesKE0RShB47zvHONMnnqB59XtiqzZCbj8lHhToWpRxLjHCgdG1gr+eRA76wLlWiJSQvCXIRJCu
3WrYilmh01IiolKtNmt8fn37ebUTIr9/r5sBQgn8P+xofFV6c6+PBi8ONsDzE0aOHnGNrJ4ohvq6
GxdBlUY33QgukRfXsgBBEIl2ywP9BDbUULCDe3PPhI/HqLSDKp2hdS1blIT97yTav7xvM3dqQvo2
Coe0PWnxoe2+YeNL6ddROTkEMP2QAzllM9m/zqmPO0LiuR6zfUh45G1zxlMFYv2IWofHfGMIlgWR
4VPXxjcbl3R3A5L4kkkOt7I201zdq6QQatJ7zSooHpBlEv/6D693n6eHtqPDzYuoAmohldVWg9qr
Z5d8vNow9+bAXGcKph0tR1z7JvJngYpJi0S74pxTC+in2vaBUGheKWtCN7n45Vwji7bG4JOSW9/X
qpd0RYPt1NoiUAjkFn7iwdH5w3FKzqs3un0/5xl2erQrGh99G5toaapM179SUri1PJUCPzLJ0Mk2
mfMS+VAsXH02zdt/l8HLn+TVLMogzThjH+FMAtEIq01SFqRGnMHvWtF4i2vXVud4iqPoUHNiIfjt
spaqZMqAvo3Bp630TtbbyriuM7rCzuenM3eAKY9BSrvcQsjlX6RN4pq670zz4smcWiRIGziXD9a4
xZD4Syxef38MtzxoKjbYvEYmokOVP3TUnFrTQ2GWS/PE4n1fECgq0BP90+z5igm7CQmo7yWYJ8Sj
r66ZSdO7EifO9WaPZPBDLcni6RWRWDhkX/jHz9XRrlwUqP3m2HGqaFTYJW1YWgm+qGGWujEJUi8e
ruOH2faIq1XMF8p7N61V5JT/BixRpG5UPFAa7c8P8LsDkz64AXW37Yrzrv0VVpafExcAaGjK05PG
3s22CaeJgKXh270haVJGBVpWwAMF44wmct7tkQc/FzqH5KDQyZ64lJoB4LWD0QoZoFcY1q+mbTgY
tTlvNE+xzr9fEQETwARa21gDlc9nPWJlfUSWmheO+we+VYdf4b6pxGJ2xkCzWmeIvIUbJA1MPjHa
cYmJQSoP/Q3DKi4a3uYwPUm9BFIKZaPSczsezZ/jP3IMFrRvVOt4pBXAEuiG20O4NrrtqhOXaYiQ
g1aRRZAJC0U53R1W3N1nlLYvtOaW+oFmiC4f4jhXoas0Ml526f0nnZRQLYx1jJFvvrKQpyoMNcVN
SwJ7OHAb/LS/bG1iFmaAqXy/bCjJh5xC8t9zQ28fmk9l1QdKEn8KY0v6u70LQjLHdgNbG3ZbU/9K
tNwOJWA/i5rKumiox1llSOqisiDEb2CFHdDjULerzhM93jkLFCEX9/Xk11vGdR6/seaxTZnvKDWK
8AWHDVbOi919pPjwFlvrbN8ik/vvCZa9MsXUHMLs0Xdji2C4zJZl7OzVibB/0+a8NW1NZzyrIz+D
k3wZsVnl5yij1TAyD5MDCwT9DHmsT5wS76NPIKCbxiKvh+WX+Sz3HXgq4efZuaDSHf8vlpFMAtgK
B/dRGwW2L6UtyNeSmYMCpiphEmoRov2bUGcoO9LlyM03seFfvvNkTeT/bLq6SacbAIQuPPpJMDPq
k8I+D0kxpY+uV1eFNxVAHJQaTUp2SxN7SY7fILdBGhuoZtc4rBL1FncPx72RMDIELJUIhBWPTvli
pJTFPYwDsNjF1yifgzk6xNcbo/icF8V6ItD5Ow3rUBWqgGL2xjnN3EvskAnOKww5pQs18sAY2Ekc
uU1KIbEZXzHaC6odJj8vOUSdyQNhBgTg7rDAswl4OckO8MO+B1IfDmlmzEAfj/D6nbAUh7Kvbi4R
Rolp2q378J8yO4r+RbnnYFNh6fiu/Wi9W7gJygaUuouZWG/7xhvuyNNGcCiXur+Zyy3R/WZnJzZM
mYUZt8b8NPLDKjw2vs7OpnydXHbW7Xk43st0tav9Dj6LVS5AgkJo1JSl8yqiaitcOnwI/gPJmbWd
p/2UCUdnkjN5Lm634g5cdf9fyzx3NqXKTQzvW8FMvB8NecZNlZ0wBTgUH1lHB9SXj0+nKodpq93y
RPkKJ6GPMcIs84pLg+V2qaRfynl0Icz/h0KHvBmMIpZYrGcoB2SW9pTKvYNiNW/6TzuEM8FbQdUh
OycUpqlfNDEea4+fL5qQ+qulamUjS5R3HNEaEQjnGyP9U1fjpuxHcP/+eZWmydmDtBfo7jsVK6TQ
lGDj41Hr0z0GFoTJxu7V46NML5SVeHwkD/rOEGTXmo1iAIRRkShWbtXxTJFZB/fog2dBJYma2Fbq
PoaEZtCAVhG06qJ5wDSjYeKee/mNKpFqaWhC3c4CZ4GEED94kzTWAusnvgSR2y0EeXxgt/p5nZDX
JGJ9lHyUkkfmg2mjj2STr3xUMh3IRjCfWOMm+g1T1uYdnHmQX5bn6X0+B5W2o9k8UEzswLXAoPLz
IOc2h0+4lovzWtKGCNpCGWL9i7VzM4uIhlvLbmAbeS80lHwRnaOr6FPZtU+NEaoe0UeO7L82Z1as
Dafu6P+9dC12hU0JUoxql3z44AGYFFpQsCTIb0ueRRTEKA43oPqt2KiHJYX7ZZPgTmLgzyR01bHn
MAH7mJXr6mp0jMenhgk56wTL2is8HsqYpM9F9l1j+3Wh2r0LoC66wryCwTBwyUYBs40hOUuW+XwD
Pr7fMy6PCIUMfg2tTTA58LK7pTssD5w1tCzSIXpR78i5Y+gyrmIz1946w1aWmLdFQNDI6hvxfEvq
ZnjVccZdyWFC3+3g/GP28ojftPHbxoI7fyHBpm1v5yXO1lclKNwJ83JFyGCljzr0bs2qmMkGMk5f
4srAdOsbHx0OslFAD7SUH1X7iW8rWp0PT6DJU85iDkgye2dWKVqOW7LhXVFxYQ5Vb7fmH85RfG1r
4NvbtFkdgdi9VqI6A2oz7EWpp65ZNx+TeVStvxB9COS5L0O8SsVsUgx4eHdn8molyz4mQtrV/wgr
XSFkQE8IeZdiAQzlTQe7nz1i9b5z6Q/ZAfLK8WbPc0OAcLUlFFp50m1SSzYjIty7d/sRxiuB5DRr
Bt/8eu9BwwqDOE3BJrKxL2XxzLgDIt0KEJ2QnwG7CdR24mdn99tvKLS0c6NdGlGlzF++rC3LVLr7
UdRLW4xS72BJpUFUnYADhBNzexHblYLaNlBJKWaTUNs6+Fndg74ESS37VLjKi4RZjwJvC/tjlaJx
GGzkHDaidm3B0FbEWKhV3LR/zPoZgoyAvcBaXZPWLW8SstmiyOYMNTA/ZFV7hNTlCVo4mim1yPZM
FWjgwW8u/1qQgg+GV59iSJaalipmnTXuu0nmNItanTz+40vW6XDHpL/V0yb9UpoCq8mk9tkCTv++
YVSiL2k9jCte16Cf4+lNgE5nlu/0erAooStHquUu3cFc0EtZ/A1k/k3N/+Qpm1R1AV6S3wW6PQ7e
xsDyaMDmKtTTOpjhXgHnOiai9y5lsQC4tjj+8vmIcgchgpuLso9NWf5J2TNeSt2f7jYl9pchgDff
8mMnNdW9gzPKqNX7CGsHTahqWN5j5gmnIWFwfqERF80Bar+C3I3J9CO8JISCKMa20sXb8BVI1FH0
On2rGuXMw138Pqk18h2TtmF/MWlPd8WyWKVXNpH6AGvBHv9ivkq4lZMm8QAKRGZLj9xp28mLCNST
Tnx1uhD31peLrvLj5TrHuEeLubUY5o5GklU333dxqM31JZ9wknXZQ4ldk0QaF50EJ/lOvr66jw7y
Gt/HD51Bl85oUNDH4P7wnmo0wnxQpqmv1Rz/4MJJmW5bKFSjtAVJCvUybjib61bKei7yCTqxOYuO
UBdRmQ9Fja1rAqtTMXkix5ci7vhde0JiX0EnDeyg9bJdpMQv+gtp2NuerrgFRY5Ft0ZMkGLQ9ReT
mQP/6bynAkOIM61GCCABKQqADe+h02PBeHsOxGmnkNYeAc/KRgU8P+wRRNBbR6SnF67HGGDJ/o0f
WxizLzRum0FKci13tkQCXNeGsa6Phyvz5PPKL6apxzp2IMaPji9qHBdVjrzplg1xKUzuG4WXkGmz
6gWxx2FSgNy7yqRp76qUte+cBOGBI4G7OevE6qj8XaOnDztZ32hg7i9SC29rRcrTdyG9COLnnd7M
b+O9j/qUiP00mMfc1RpdQ4rB0QV+VUidysGIQ0w1DxAoGUNYkbDxkpEL9y3lNmmlEh4cmWi5Fbbe
n/fciBg1if1i4RqmrLH0ED90G5gRb8mtsW9O8630ZCcnxz8Jk1y3vH7rrca65Rwdifu+GWQUgWKV
4vpqtEQ+y6vuIrFRJCLZjCYE73eQqL6zz2PvOiOPNDneSPOt1hHyLEmh52RZl63xteKAZU5mfX3c
nKS/S1y1STc1noUkw7r5zvWcIFoFBHUIvDGVpqqGysy3K9C7bun4SUSPCVuDtDDInftuA+9yZqCI
NR171c2eBd+SCV5PrnBGl9MbxicRN6W2GugrU8vIvya1qsxhjGoCyQkIWBIojFHiCq8ERIaCP3QE
dfF+FMnFp+PlAeVnxg43PlFtEr0z++dbA3htCqLIZK4hH9FmDnbul69nfSVxifpGNledC0aY1biI
0eAaNNgzfsTGYL7cGf8p77quSajJQ5f764UFNw8MmXgoT4drrEGbseoyF09N1sqFEU3mMNqeVrBl
n/d0I0/R9zoFUloautQp2W3sWsn7trjjgkiBTHWR1thXQnzJx8APed7h3QKnkH/Ld0K8JFWeeQtY
PPQzvttYf1hrU0woTRI+Zak/lRBOOuHbUZ0ADEc8IgHUdufv38cMWQeZSOAnLAC8fw8ue9lrfF6t
K1xH5rqp8MRUjVg8dGZJzKOStxp+99LbIsD4zIgTMkXHeWQ6f7YZzDAsXg7K+nZMBNNv/pqK286b
tGQibhyRNO94bQ8+lagvtW0mzpjM8e4u/uhygLdqyc+AJqww0O7sqgcEPVBPWWUf9M3mFEbYFjSI
h4SOQkzDLZfzcVoK/pqpRKa1XENvRYkWD30opbXukZG6u31NYWkfosANKkgUpiFyWrmGya8wVNkk
sTpiv+6LxmTcfNQ0VbpGAMzd/c9fHCo+tINjmpQSIDCJNaiaIwpD43pazVROFxtkSMIm90/QJc4w
v8sJ9cJvcWCFWnq6gxX+cilpbjR+ynoFzSBWaroLNGqs024upF+yJ0MxjOpKSJ7zYxdJtLY5bPdF
9/nS7k7mPyGcNu6Jsx8ce9fmNP2FNHMRDiLvaRZMqN7o2ikzqwdYvWj5Xr1PwYHFG7DQzRyoWVcj
zrwIFGJyhgNsSSoz92Ua8dkDCSLpFLCD1tpDOJuFSZo0dtriYpANM8Vl5rdfvdzTgt4dGZrcPcPo
kNARGXijqUt+R6i/yEV0zDCi8cciHrq1/givGyT2I/TQyuPO19zNAyn1Ee/TD+/PCfZp2dW6VhwP
b0gDqUFk3kKtUuCOUxqoOE34ZiLnOO1EvDMFWU3+EnNSOF4araUZJzYma86AQCZGuzqjdqAwdiiN
ImCDG/k5520hqCV2s4dyMzjAS0+x9hX1zy87pTljgtXZvmeZ+SLAS2PfjRYNR5ns6pTSs1E6MwRz
LV4MBKyEPP9E4rtIP9oHh1U1B86HJ0WMcmQw1CI8S2TSdtz0RV75dYJHjQo9PobzQI3b0lJMppGE
KKdHK8KUt/xF7X6H2aPMAeQYuDL3PEbbCnYUlhoH4UpIuFLLkrjX10tNvZXEcv8ZhSooACvl/Rnd
YaA5a+FxMfkt/MGSq/7bwZPoKLKbujB2L7QDBX698nBfPFdkfMo8ocs0BQI5hHtZpeeRyRNHHoM3
hC+q56Rz9IUUc02o6M4Xh7+jqKEDxObz4lObb5myjtHfsDvIttgz0KAZ9LzseZ7dNDTUqhlU8upd
N4DC8xJX/TST2jRZzWUkLDlhDkrmr8DmLgL+FK+95iofGpdXyg1yKWoUoISoNjOXCSr2oz1ZFuR+
vPziFfp6s8MP5DSO/SCmSMw01k+w9nFQS9uwUHkjFULdF6tS+9oIV0M0hKpIQhl9V/ijULz7sieo
nVVs8HVr2LUi6AY3gBBzZF4vjI205EyxoNqzevV+TRp0wgRfJXcltIq9KAbjCgs9en6cdjnc+iks
ShIqdpfVJAlyB6RWGhzugassbhaavTEo4fvt2KpBzDEualogo4/MT/g36zNNlTX5yRLCW/aqZ3o+
0mP/pi6c40Scfm9Yo9n9H50MFaxJhg29AY0HOZQBuxR3Pa/DRli9BUPHLaQAkeTDkTsW/Nj8lRPe
ELj9eSMTkrmoADU1rqaMnygj792wbS2b/xaOq+zmJ4/f/fBejXZACdX2tCcKzlzvrWhz9gN3ANL2
QgqIVpv3aRwxwZlqwHlrGeLgcu79Nyw80c+81/7ApqVw4YLdjnmFOIfATNra+R8RvbZBdyh2xvvf
Sy0tOe/lIP4w8bGLBZuInJ7iBIqf4jwVzJrNLBemVQHu33GaGSRnOqUch9MJTKxvL23p3V9ba5bb
CdcdKKnsIeH9/Th0rRHqcpcwctrz1K0iVFlurAVKKd1GA9jobL8InM2wIPesDueD4yPwZonY1Sdo
11ZImMMQ8pjDfHAHl9REdWcucUM1kfyH49oxO/QUzlBmAW16f5Zs7z6V0ZA58+mAF4mg9LQJoMCY
pJAZfwExArOlQsFQi73PkqkcX5Aq1Ai0pyKvSPFa0PuUq+UhVW5Dlq65gAmqjBa/ETaEZwe2d90D
Iupe3oUcMeOTSNc4WDsq+qtBE9r2o+vqXyiPy+seFj6NVVVuQ3LE9hbqTr8WuQG6QZ0GOKRiRlsO
3XUm+gNNGZyAX+QDx9OO3SLov9tVT8MCkT6vGftmU7iXdhMM6sVFcgE+4Q71fUGNlzxxn+rgasGj
LxLjqxg60hssvjqnkYTM1SaHG//NEppoa7FC7kppKHS3Jj63qv4Q3tfJTaugNwPkUgscT7XJtn35
IHvx/iLa7tYIMthbH79dfCh83YuL05qo2I18TElnLpTcIMBBygbpsXeKirA5KEx9kp8M/pdLuoQo
GK5h+yUhAy1j18DVXB+qOa7Z+gJkdrt6f9oFDj8mvJ31tAIsfyNedajPmZdfydyeSRYjyG3m1DRh
2kA7e4+f9LZckBJnpZCV8q0pni3t220pAICtb4/mC5n9ox0jujuVfGmqt3Ctw173Ndy2SDcMYfEk
Njo2RdbTuY74h3H7RBFSZPIF3/zspUdXwQQYa0kuvqhfPGJ9OQzRMfDKFSDyKBOHmXNecXjU9Sb+
xuKuaWfTCpWoLcfQkcF3pxIUpNGZ7Dr/bmWOgUp7vaRrYLN2q0BfJisrUcXDHHWZNzt/WZvmRVrq
qGTbp0UhCNWqOmVsT4dB0vmyA0tv3veRAaai8MbFRiRUHjEdoAgPn54RTilw4SAKl1RP7U3cFOH7
1Xrlof6EFhNnuW0ARSsCqNMHn0rEu3ko/4GvzrzTHal3oWkokQVPFLUWVVgTi/I9f3SZeeXeCbdw
6FrTx3ZLcadwKlW2QKNrJhqVfoGfRiEWhn/VrvoSMyIcq8GXNo1zoGLelC9HNesq4lBoO1CXPzAb
3SqH5wZLaNVVrwW7g/N354BWjqQeghtGMXTQMqfqrCDkQih8yVj/JeIm6YFHvJwFdpXW8BNxkbGC
uvoP4WMe93f/20/KfkCDafnpNt51eGTcPrIgu5YHqQ4OFJ8GZqlRDR68SRJ7rV0DW/NDL7XxAPhy
y/7arWdDjJpXjj0oVbsywFhNTl7AqbbIv9PHU3HtCVZ0rdb08p1Z2jT04RGzyjMy+LqRtFKB6HyX
LQ41p5ijfkms3cpKW9m77kAY8tTXAmFPAuUqc9mYXIaRWZrksrNsYJbaIoy/5KJCl/B4MimpmK8Y
eP9ZFiWC8nWTL4QklPlCUI85KFuFBmv7VXxZyGxQkDI8Z8/oJjGpuKr8wbpj+Gdzev0UOAnDR2k4
8aSoDeAXehEP2osrrZaUglW/MoXev+tN8fWoN0O8Zpz5q/cXGC/ASB/hfgKMEdF5p2yeVjKIHV6z
PmxVJQNz9indfL70KWC1EKhG2xmkshtvEy9WVR/V563QhxLc37szgFNzgV20wF37Txt9VeGgDsiI
5Mi72/SwyA+v6kNhZlxadcvX9ryCW3NSpN/MpPM2U2Kn7qxRgKGbDJUqWuVcMjbukqAoD0jvuoSE
YdJ1RrBy8avZ3gWltssYHZQi2H7AeQXUtddJPzqThxCEI7DhnUpr+v8FgPjO5yTxx1G4nWub1EhS
Wa4SSzKa3kG73MAqYrucu1XCEuLXuzVtpuEtc6FsJ+z4C/k+piwQn4XHPXhjRe1qhfzWjB2T2EQh
q+1/Y1aOLhU/4O/ot9v2diEo1AmpwBj34rKz8b0Uut8e1ARZ18v4pyrwlMSa/0POR91W9mhMST/R
X6hTrW1JFbbUx+MJ1/JMEmQA7KBL2KcpVw6ayfZje7PxE3VrKHpbUQHFvVzzoFp4/Zikv8dSClFo
EZ7KZKUOyt9ZZh9UYqiCaDJiWTuIxrUJg9KiESP1W1nPzbCFYjSkPol+Y3j0cveJjLDWicFjqy/4
UHf3geR9fYcNwzeTcsX1M7LukuI599kqHR/uxKGRM+perNWFJBDcwv9c1dvkghYpNLhtr0gPSw/X
flC37/6IQMP/nlmZV4Euw2bUyWI8qTghHjarEeCEEQrS3Bv9ihgVa6124MkW/vldWbnXUnqQ+RPZ
P3tIrGEFbeWEteTTgWBvEW0C0XzPgvcicd9jqA05dYyT2outpdW4b2XoaEWOc0Jtw2ndqqK1yOPw
bnEC/rlgPRvkQKTj1kZgJfVTWtMGuX3N5ZQjylvnInHMEw/psaM8RMufJ4CQr81cDtOkIxLaQ9VG
PLNyGYfkVme7AhCKTMd3mkt2BuSKEwSIOLYo8Y/fCDr49PbqX8NGPGuG1iHObefnXxvxIwaRBYNC
p6xA9f32BZav32quuWnwB014nyeY4dleAR2hmFSyYJgsOwhOQSrNfx0YsuxDrvyQOkijTp7O8+Vx
f1FlLKmCXbz9GTUDvbVPtdi4xnYLqPkIOzxaeuPXT4cphhIc/3vJWkWwQ4/qDgu1/g/WHrH9gNqZ
DrgXTVRvq4XCxuYaAJKjk9grA42w3+/TUwR6RVMIsBlU9N9LdDJtfV4DsroTgvKHq4Tbnky3BVek
82mvwKQIKnbOzbTY0tRU8suk6Z5zZqpweVtB9pCmn5pEbYbs9qHs4X1IrgKWaDVPflOJsUE28Nqp
t1EpmbHPwZRwwdm8aoxgDFFzoqX0W6hskPSWfzOskGA4NMuiC5OGLtVRyJAy7q936XR+e9dyPRPQ
Cl81+4kAUtVVzNpNXGtRGwXow9U4JP2cxArX/ihs4kGPgcBGm8X/wpxk9QkQjYvW6WmW7Xjd+Ohh
tLHaFdKo74nYC2pw8oBPL94e+RHULJpxr46gAoQFTaS0KvZ/Clbo69vIRHEy0sVfRGLHnyoNhILB
ORMpfEBbuHxpdJuXbIyjx1r32reKZphSBXy/sFQ3wPiAj+H4YRfMc/e/WUZ2CYKiExADXyTYFdS9
CcoJowitgO/eYYKgEPGOTVoDKRVfLwNehlZehYrtnM7m6jGSYQETksRpWCo9kjnpZ0xa7sgoSifi
0kpFoslOhwYVwkqormO+CZdf6M8ONFFb9vrnrWVztJAncUzIBr/w/YRvzn44upx5nBKdgDeiuWlh
Ff3uZ4eJuv9Ybu0h/mhHlYpv5LsfSAdko8VIaVtNhJFP/ZPcfaEtKNLqfJsLIb2zie/uUKangQni
l/4vd5Z9Y4DoItKhr8k5gpBdB1c/5GXJKMfparJ9SHo5jRlPHtWlQcnXJQ7ScnbT7dic04pGicK9
5vx94orKXmibBooPyjz0ieFiD8RFHsuiBZ08iN/mi726mq7d8+NgeZUvOvC/yG/wr9Y586RtyMqn
nza/pTEYxtK3uqadErpzEhSfxspqeS6YrlZ8vcc8cxFw2t1JTmLmm+0bodQsXaO1cDsFv6JVa/K8
vwxsr6acTJD92zTpFhnX1Zbayq+GTuz/ozVj7RaaIt3a62AZOYfo8Gcx2Uj0Qc4wu1GRUX6je39Z
mEjjm7Ln+JNdzustchb8px9DVDm1JY6GZdZ2aQrj5t9u924VIRZ32ezUUIXQ3VN09q9/mzbRQ5Dg
2k5UOR3vOFNpO+moa6roF8E+u0b6F4Ei7XZGYZOqDvoPp0/O2uk/B201oConnlHnWVWu5V+Ogzel
mEM+OrO2Byha2j8qTbP4wslGX2zcCQArWyVtUJ6AvEKpE8r50Lb888tsLMkFaBKdFUujeseMkFBC
yOfAhKNOamO7WKnqUT16EAUdUyEg2xhyJ1xOg+h3uQ2CJZGIfS4eVKiAq4REtTLkyYhOSML/NSC6
ron1bG78bfcpjkV7q4ZYiEo9wvmEmozJSe2xuEHZ/U+HvbAqJ3nnF25fZz0Kyy9EvaQgdv4VbKQC
WYaDI35fr3cN0rsyFzVOSWwYfs/JQnov0/SXMzPGhuWH5TjiokOiL65zOd4twXp3Co2bQdqk7xIc
ucpa47V0i+aja3333vgVBMvRymCM+qZZAWEOIdfn9WGp3glVZ5EbRHLZAVxmFY5Jqd1eACx+1n8t
+XXoYS5Cr16MirS6KxsjCfiW22h9u4FNCehgO+lQVAQjFXxTlZbxhZqIrjBWvIFYD9tQqJ7sNMxN
drKKlmrl68/9eSt5Yalwyk/18BKXxn5TJqnrfotos+ejtsni22i804HZGTQrGdMxVcHEl71DI14u
xicHWwFN5krovN9jnTMeu2DU/HF5ozstYCFMu+DWhXnFeZgqXs9KrY7daMzBevRCc0PybQb1/WJt
VVRxqqmX+VP7shVSn5nQQArqfFlEz7CMK/zoDcGTa94TbCGE4AMKmGQDSL+u0ZJRECdZNq0mnAYL
943HT9slRhh0rgV5VnsqEpX5qSj0uZnRfvg0Pla7YEDcC3BwsrijeDCU6WCKcl5QzKMMm+mcVXCN
/i2UohEehnCnhPJNKPqvVRhj2GB2+UnvEIShv2JNX47wxFHslQixNrnUOhNHC27Y95Y3YntbCRP/
3fiG4ygDCyl0c6Z4D2cf9co3Oj2y7KNdfLyHtIPZI0x8KRVO/nwwkD/EgaWpZvlYJeYpO1QbeOt3
RT56vUVpP7XXG+6kPXYHoB6fb9FTPq4yj5ALjjf5qG+vSifFxORyh+obT5EnatYAGJohmIqkRGar
Lq2SPsktLyoRwYjNva9/7/VqgwiTvBdExvuBu3V4UwF+1Fa9BKa33IHEQDHJe8by4Z1ww9wE0hFP
D1YIlIIvY3wuTPEpMPdAhUH/KVtafttJLcnlUzyfERrzMkKP3PL8Wg5SQqjr51xJ8vjLGsSG6HTH
weKMs/hy8mmzVKDppFgdmi94lp5RKoqR+NYeacaGz/CdKpY1Y/jZn12y6FMN1BwhjNZcLupQqGyr
2SHAUOB78r2ycbCXHd/Lx3/+eqm3FA0Eyr0sRwgJ81POiTHTXb/ybeDvYlHlF7dGLSRKyhjR9jcM
JLUPb4U7FcosYAiCSVXJRaMxyGevLQ2qdAdosW3376gVYvgj0mQSz2cBKCs+iyYg920j3/rVuIjW
8V3Lax45zYzLrTuKhfYptHXebbnSjWcc4kHenlfQ6NqRv8fO9aQtXFilfjDVWLiD6k1luITnBvTP
W33Czwgy4c1R2OJ35kEEip+0gzWhToSbYdgYfdTrC1U215ucOCKbWH0H2VnN1Dqx1Cfm3vOnfKSo
d+dR2cXgeJ4CBIn9c9mld80LAqAIAC35DXqGlvSFLitCuWrL1MNeA2YChAm96WbDN4KZfDcaHSFK
aZpBUvornYAncObuz9ZysO8CcZX0SkZa9VrwBmEw0m/V8+GRnD2n0PJdS6F2McKv8rSkVbe/4rHF
/iwxJmUTscYlD88VYG/BgFMGtP4Mu9q8VrOfNiK7YWVvEni1ULqCdfbS859yhel9Svxu3sxlzhH6
f4or/bnfYLzHmfcqgIj6mx0tlRprdi6F42v+PCVUq+gNwGxPqs7QxGDOGaoQfMMjFipHgCauo4vY
AWb0KDMX7kLj47v7If87S0as7BWi/n/IBwkjAZdbNW9RUKNPjfjK4U5uoSAy2gPvDNpziTqGzKYQ
bj/F6FY2Dz8IJTft++aHITHnB6BKM0xcmbjWdf7lwtR9YV8vQjCoyv3kM0MbkqfeDlnaLkGRn1ZY
MA8c3INOBEVQ+gcJJa1p3V4MsJOXfMwGx7MABIZN4ialu2sXENvKA9oObqdJlaUKa+r6x+BIDntY
gaS0YOON772VNgrRTnX5WVumkUZWI6uPcetxZlH/Pai1pgFKVU6fKvwo4wt2tKGgVbmw8fao6h2j
TlEIFJmbbpeMOfG+gb8ktwZ5Pgy0ZHLjTR1Mx5hrWoo9RrVncp5Ts9tIUNPvv9X9ETHvk6Rd7KOj
8WfobdnvYco2tCIHB4vW0rS34KSwzWkooDj52XHPSEzuNy/2YzlZFQMOj3Aa0d3u/plOkq+JE4Ng
722zmY/ex3q+iajYScHCH5moOoZdTC90JssQwls2GBVjd2lY5k6Z5Ffj50Xap/ruOAW4L+pRbmSF
xQTnY9RPoZFh/i5LoaPwf4EKlU/nYQuYI0OZ84sJNcpk9d26hz5jEIhrw6nuhayEk4d75rD6ULx9
6w2+cmuhZb4qfgASZ08ju8vrT7a8O1NWdUxg/eAfrdq1nBYWYK6CzD6iAAmerpSlNcNOyTulaWuX
DKC10wId1ORUd1oDsbuK4UGp4WJuqD92zmEqLFFCGyj6ApQS2oqupvf1ozH5uZDHlGQINohFcbfj
i2uCaFWIw39cXAtHjNvQQ//XVJgmFlm7iopCywPvDOQf/c/DkUr/5tz2kJKKhrfEBErdz/O8+lmp
5Q4aMqHZq3PqGPUW/QYr632I5I2//s8TjKmJ22B0mjbeGLEOqN2OW2wK9bXcoaSDextZgqBWiEEi
Ql7ourEMuXupnIDZEwiUjYdndXm5b4UwCNTiv7hS+i79RDRTVsF9Vdbe4LI5P2d7NPckCQKMO/LA
XR5vSiIqEbIZARcEbK/7RToM9dBloLiR4VHJzdJBBSbCuh/5hSDwYB/yFky+qQ8CpNv2RrEWNeyw
V+7gvuTUmwnr5jxA19ZC3wYusd00hRWoJvqjaU78If6fmJmOhZktSh5ViCng0I5HX5GYOUcYOC2U
O+JaBwpgbhequKLivWKyIDG+hbqLGswDIsFpNptRatzXbEdpkjJtizMCPTntvo4vrsB4jJualpf7
teUCMUWzmRqRfm5R7EngkDUBZWVLTEKHJS7HOtFpR6CQ+UDCoQ0yDw4QK4K+jr53ml1Q2cm69H33
guBDsUvsDT2ivitEK26EOkhAR79SnEBkX4Sdx0y5D1VuArgCpenGWnGXaeWaV0vWF0yt5Dji7R+3
6RMwtmuGFr9YC6cLW0z1zrzFYf0bDSuo0+RCODldBipYF2PLlyEIEAoMVNGrO+L4i5czaavoiPoT
cs5jtPbhGrRA7Di5eTDV+nAGNlKCbHTnCHvbWy8FebbUUv/P1/1ahde8PPlKXZvU+NcnYV3eMqDz
uz7olRuYXJdfSYiaT3H5g+4JeqRJZhXs9PV7jo18wvCdrEGDKUFd6wE5LFinCwpcKAQ3eKAF9nW5
LuJRyY4FGomnMP0nFnPgYj0VRexiDu+QWhnX+6uvcK47+/roKaka50SgPzXGXGF/Ut4S8XLvfJQO
UwhZsGDRzAJvCPcRcrIVtFWdALbidLNEhmmQev/k2j8kUEkS0tilvhB4gtCXG5HOwCjR7j88Hbgy
A3NMlj/WXSoCmxW863XVjvKsR55zv0FujY3zecc5iIVfDdNMjSmiFER1/qhcy20FwTUOw/nA5zur
XazFbtVduA7G0EUya3ovYkD5cmW0T+AItSKDK6otmzsjFdEswTTLk92DhhLVDd7MPCIeRAxrpDVP
wEoz5utxrZAuKSYr6jzTsY6DXlZ499UFNpLXrRz8C+1iVqXO5DB8IgpkYbRVyBpLpVW4C+gG2UQA
RNSRyY4vtyNJ5MzQADsa/MPwo4yWpwYzrznP73i1UCUoGygco8FH9mMDdHp9cpB9Ej4/nq/Ph6iZ
fhcOfqx0iKsA0zxNy45jvXDkV7KTjfqkzSrgqL9l56mZEY44H9y9rr0oMZKiiFw6o9tLQtPFkGOg
oK8sF2ttBoNbw3fvnTJWzy27k6eelYq5SUnGaogHrJyHwpoVKUOlNhr5u8YgmNB+f6nlwg0w2wkt
zOXJrMjv9ouMz/InJ9dbGkIXvfxbLeXMw5nZrT7eGF1VUkh4dJtjksbHTc+VbNFDEP2ZPzSuRI/m
cy6drjIm8nEeILHeyTP5hpW3D/KjG5Y9j8lhytp2nOGK0JOL89nIe1kUmY08XqFOi98fL0bRvDtC
gC/4bTDGWB4WmFZtvwF3yV5mo4ql3IDgLw4q8iq60FQX7OIvdD2+sqEBFMfPVO3KGf2gO5xGLqxL
0TqUWcgts6Z16N4qI8QEJ8UeKcjo6R/abEY3HAiyB2HOinZnzyzuNdDtFF4+mqEHciXTcoLdEhGl
3MLLH2P+hUhTVkjxI7G5GGn7xaQHbknlvRgBnqrjEsOk2zQm7Oz3IwTRcqUmE/cBprTvBP2sJ2s/
ek25YHa4j2GdcXhSDLicFtVm5nEEAh6mZjdJ1VRxUbm4Na1E7OWbucTr00BSK1eg0sl2UL9lZrMO
vXtpq3RPBXh7qJyXWoXlfb3Dc+pJL/I/21F1HVygWHcZ1ioq6n+9WH7WjkyIwHdfvfm/QENtA5Th
FV3FUIptZ5YTVksWnlI2yt8ojnXVyVfLKFVXsOv5Po7Q4066xp0RiRZt+leZkBCkXK+YHZdwi6yv
Bor3e/d6AFa+1tSiB283oMEYR/jtA2ssN+RtwDdY6yIT0Y4F8TTu8vz2NG0xPI7/0MRPa+vSdyd2
wk19co1O3bpLd3Y5jcI2vjF8vcm6f9GiTQtD0egtre8NC0S8x1/8Qrq9MijKlVw1fy2h2vYkcNtA
vqpaxHflyMJU+oPovBUv4jju04lk3eAg1vo1sTAWXOHdWU7aVw+gCsCHbXhzNzNDVGCYuednYosw
RT9n5c5B0lExehFW6+IRo1+rQTv23A0+WL/y1c+rL1hXHSqnoGI3b8OSethTOHYYlPbgNnuS4sq3
+YxlQGmZ2sDeXNRRyZ9IVyk5SsGgEk2kZOXJH8CIh8WQOdezFNt+OUPVop8r5uTBBIZ7lTMTVDgF
M4waYNmvYjSCJgzQacDCazHUpi66PcnWWBmEtrSO9eYDJynIiYdB7J2blXE8PXSjhvH2fNgZK6zQ
fUIZWvqVY/pq4OzpZF48ha5MZZ2Fsfto7wmQPBxxiZ6wmc9mR9vK9KOif4E0xnevPL9m69ecN9xl
78eDn4q+0+AUG+Lkah9A1RUqiZBC8++P288NiD/qB9IITi+/NBml01ygV5l6ZgEuUdyp64ZcT3AX
SjFHmh8T1cV1VTAswvR8Mr+9g/56KfVL7KHgZAGWyMUw0xjqSuqH/tBTIqjuyIpBxV1Dw5up2nNX
mqGVHOiD/Bb+xpk0CHOcuFrXdTs9898QiQO06iK92A3nbrNTHmPZ9RYCJ2XPqIs6HJqxFg0foh5W
l/+bH1N1EultyBiLIqK97v/DGSXYzHBBv5oGrKTO/GoI0vH9rbxZD3FMy3poBwQnkbNusnfa9x0a
KLmdg5mgqg7R1H36jPd4lQHPW01Q2AnqzxOUN26EWavWKM+VidLZutb9Jt555OJJwL8r7kwFaV+Y
1/M0NLbPSmRLsF41s86vey8/DXH/7wu4/Qp+OOSo422r6UamiHsiSmIamVIs2eUZEyPE9LM9n0yf
Nq0K5tl+u9503qvgm0SSDpsfivoTdyqdoNLKxAsP8DmX2gO6Dw6ZWtbDjWn083Vl5c2faYMwk0Rk
h40UF3EuSxnQ6gnaFAHYSQ6T1jhrwb6oAo+jUkJnJow+KfLrZtB62mN8hMTkLtwdcmJ1yG50x5Pu
K8VBdIj2S2BmdRwoG+rhc7uqF5dfurd0oh44pWDN4Qabo07HbDa8JpIgwlwrXa2L+fnNPCht4jHW
zEH031R7ABAqdxycRVmy5k1WWDxOSVd1AzweHu3qTWNToVVI3oG+qC8truhEIsP16EjXPMWjiY8t
ZqFpoVtZ/tiYPtZcX3IGF2YUWcBCRjVWV3ZkYlyF5UFrRjZXMcCVllU06Pij1Bi8EaCNJAc3plJ1
A5RainNpCCa5X+uKA+qwR9V1AZC7NCC2DxEEeJizplZvUZe1sUriVJv3Ijh1PpnltYpOr2Gp+lzz
u9XlyjrwIH79w/7rl8YSxko49a3/sMwinSjjuQjGa7bxzQKv0N34DkmLimYf7hZO86jGEh2ss2HR
bKSKqjhUsu3Ec6ERzMKaPg1FMZ3dBLWxq9mAGCwQtyGcgpDw7RDEU3uaTLC9L/h/8R3NcGb9PCgE
UaaBzYA7pjOJhs5u85+ZPJyzSw5Zv5zfD32Aw7G45sjYv8p5JJn+hDFfM1jEKa+gONVaZOUJXFjG
7OPfawrbvdlBhLtJZv/8jZK49Q4nuR1fVhQByulQnHn5LVVOsWT/IzQh8xPEP9Yot8iCGO9Ojdyo
PH7ZkWPow2Y6K2aWaJAB9rksLtR6N2JoePymmsMXedNZV9Cpjlz7RiaWzAub619b6boAq3VZwnZA
UpUJWKtz1nbG7NGfVN/W+KZ6BjxdWaGhdAovtHT9a3KRkc0rfTL4jsw/joI0yQ5p8MlZUl8mUiPw
DTvjijFao0w1qLvjQ7jVOT2ExHflWZElUaJ93zM/+7ylcLuEMatrJQx5LVypE7nC0oGTrdSpnTPM
DbtJLJAOeEjBpU6LegFaVIu4OkqhHC0kktNU+t87zo02sBhde1EqcGwla1DbIlD+tGSVE/WmDacW
QfTZ/1p3U7YHc4AsrNGmpv5Au1VlY3MccYWVDxAMpI7ngyazJ4mSaJVSrwnQirNb34QZB0PHIKdn
3cMIjj0FYRzn7ToiKhEoiyI4K9R6AP6oWkDgDgtsVHzwocjcdyQUgGwNrLBAl0NFzoo57muhPeF3
dCZXqopX48J8RzA5RkKO0BYR0qBZ04G0XhFAv6gn4luZYreoqVRLG1e3rocE/A/pZA6jfE1so/nz
+P2PGAKWwVYgZPdDsw4qXkyZ/P+rORHXIRoiERahw7FZt7f8Ow0T5RwwrSfv/f1R+04XDzZkjJXl
F7s+gRWMW3LsLWl4AViQQS37a/T5CB4OwaxlfoO7vITm+aEuHT0VeslqSjQWFPFxhjtC7T9yCa8C
5aOsiOPh1+WOXcPC/xNzIzraXelZ+whd01YN+iH7o5ijY4/Y3Y0xVrfEle1HeO/syzLPG7dRfyVv
MpNUHarOxT+lNsA2do+EqgIbUmR8yGp4+hVmVIqaqI2WG/60S5Fp1d4zDIgjjILA4NCTcznJEomV
vum9gx+eacP4hHMet5LUztHZdaHppYZRTf8h20Azeex8u5SqLCT7x322+H/BM4x5mVPG0OeD3A8U
1DVDW0zWyHu9Zm2eGL4r73wC8+87IQneFVqsoUtVnxLkR5b/GU1Mwcy5YLXtFDxF0dazdLZz10e8
P7E2WL2e6Eg68Gi3vRIUCX8PAmfmBF5ysr+SXJmQBL/QOXa1GD+edNxqlKailFW51BB7s/mMeHbH
GEIQVBXlySBKMv2bwrrRZpy5kVHJUGUi7CWM9GC3nHz+xG9EchOXaNFK4mkYeVHOw1ZXO6YDJX9M
s6BBOiUNTbOBwzMjIzh3dSenJl6jxYAb8OHSrRsGf5yAYcuAFXdWOaxJHSM79sr1ua8SfhWfi0SU
mlbGRmRNxBN+7Kl9sThy5ClNs6KxAif+hSbyM0shwcRhC9YZoyUu6MwAijyIKaSa9ZZxzUNdczGZ
R+cZ19KsfM78VaIGjamw11ENb7K2s3CQnHa0TlezamITx0sAdsyC3k5EFYt0SA4/PlmZAoyQ8oij
HnTE9hKdvg9wMSss5B08hluyMo0kycPfeEDL3uQI7EmVfN3/v3OCauj3ViZnsuI1BaR2ncvAccOA
YiCTca+J8CikZbLve1r0sINHxZIeh4O2h423F7RgLXD6BjsSWzp65gnm5UMINfEDPF4nRdzVFLbJ
16viFGln9IgHFN1+9AEykY0TeRFEXHez1y20L3gwfmw0SfngiVeyX6KOI1npLABOc9kNvUSusEMj
XqpKgyFcHCXzv3iVBsT2upoWEGw6KdLyy3m9FkpPafzNGPn5e2CeNjLTy4+zW+44jT0Nm+l+Xl8K
9p1cSpyViRhJxnaR5dHvd8ojFozJ8yDXySTx/OXyiwt5Ns8fVulX/dGqGwAkzxfuhOrR2cn/BvR3
u+RcmbiJncEDGc71nz7B4wI6ySFzLzNHmtL85BjG98T6LcPg+TxOB2NuBAS1rxJkIG0nvt5ptV5l
hw0ZekaoRGheDNryaa9NZ3JmpxuD2s7sTzT00CuV+/PL93jFLQOvW4yYf63qyn1nB1pwiV1nt35B
4OBVPplz7km0Yvwc2Z89SgYWdKdwbX/nFAjGNz5vL8TKS7iM/JgzokBA271dvskYrrXRXxVzH5iP
q/ymHrBMLDr8/zy/UNv4q5z1xHEJk9dDe/0YnvpMc/72bgnMlGp5opXP7dlOiaN0vYe/90jK6IF6
JU67Ar3v7l5XTazjUgyRhkC8ObyJcg7L3E6V1IRgYMgkxt6HDF3gsbsJDEAb8OwQ0h5zPicvLa5W
gDeRnYC/SzzEKpoW7D1+K5ahy9udRaMw4C2ZZsXClvq3zllwutmj/QQqkVPj4DvyBPhfqdJI7dZA
wPMX1c5o1pMzFnHGFe0wDcXRyPEJrZIVieDNo7W5wfE75sQ4uJCyp/DEwvZBHQlDWCe9/lr1y4B/
LH6NEpIj+OrUAhsReKiD+DrOIwGAJgnAfbc8XpKrpbEWm5ppokvjX69Xkwbi0/SeAXfXxG5ovV6A
2DeKlyOmlZAUrM9aWZrEPRtzaZX2Umrtnb8iY1Vu/eZGtEr1UsPPomccf4ASmuNz7qj3fLBcGJ5N
ia6AWDTvVTSI4yyDCOeJRvs/sa9WqpZURs8WemPPqJHTEtoZUVsKHTgu5qOgb3v7t6otraNaSpkO
Bh9wDG+5u55vHW/Ox7B+xYYbqZ02FLWJgs4I91vX8bcZGm1gonD69c1PCGYjx1FyF29eI/6f84ms
AaI3QPFruPTbtRL0b0FhiGqE5JD75O47wVVOHZTzVND3Awn2n+GsGfRRGXvtgghG0W16FnDRhe1k
UjRHSnTSGv6HxKz7CAh6/nZeui8YOB1rt5E1s6soADTiLuvq7+E887K0ZLpuvfZ1T1Hr/NZWRH3W
DsXZvlPvlyYJsvJdCmPBLAjKTDzsYNLl4gg+i17vuAtym0q3suZ1n1yh89cyM1+T1bX7JTBAc4TL
JiBs6+XJ5fpoaLqNpUhH18ohiUGqyrIeWH8Up4pwztjfU1R7LtY0nQR+4V2YMBUxZN/etWTRBzQO
OdZuOFjRZovT0FUPA7XobOBrXtGBrnNgP1BroqhUg7R3KyGM+ojMCLjphnlmXbKZgEzMoTiohMQ4
bgeYgAJJp2FsSGZiK2qK+xgYljvbHfx56DElPVZ+qumNZy+xwjnaiD5LqKzD55nrvIBVIrcFKS8v
H5bBIngE4P6NHrSLUWhM2KhxczbrRHb/JTz5OvmqyGXJ8W/fPtEsgsq8pszH9knQummgBlQ+WBuX
zjhA563oZeXkSk8GsllH4j5IDgtXMh16pDKK6EYIVb8IDTw7hqIqYU4Vtc/ZpYwYlpAQfBsRjaQO
BJWBLOlpFjTwsEdweEOpmY9wf6iWEjLUCIkXt9O0GVRB6yYvO88PRSR8o2aK+dhYsgRAbWbEDqGj
dNBWrdRZs2gG8t+ejvM1l55/VS2f3x3JUoCA2tWWdiIPecWDIvtkhqfzTAww20dAILRTY13dBnL3
nkSl1Su/amy+FbTsFKRz0zewyKGo9VZqOGhfKD6X3JV2HeZKeyxoqhGpZlmKdb1MMOf7o7HmM9ah
zMKAwUtRxreRqn0IxjLBMqRQaFRkmKJlYrSce6ka8vXn+kukFvub0Cx1OdgAKJes4lPwHkQYppiv
/Ffmfaa+y1FRUAi1P+5BdvRgw/Lq8GAamnv5lwZPC3AcBxrcs70F2g5rnatDT0BgvRz0YNVewanN
zfYU8KvtVOSe7Ekr2w4KdWyAWA/LEubWYG8MNkx/NMTj1oTAFk3LfmYUXX9CjgJK9snezvawaWAt
Xt6CFI3jLnKBmo48SBfKhK0Rsy7XU0YYwzrxS6NyXXm96Jz8Ydq3hqnWRoSdjtq9Jiaourq/b/IX
d76kKfF5r9zlHy58DDSS91YieJ9z5MRY+rlEaWyFwrz7Dm5mKqsOhmCJlwk/c8o35kwrpju65nSP
HDlLGFaou72rwC43sY7JlxFCTU3xww3p2RHqouSjtctGsrTdpFBXTr4MYV97nJy2x/5D7IQljsuF
eEY6DifwQq+GrfJbgUP9sW93EZRDbLyYds3w7e2Emx1T2UefdGOGnj8aBpjqbkLoPsJfFnLxcAZq
U8k1heAdhf8ODXBSamraRnBfqft6nYTn734+hGO3jpP08nWjk+oFE4AZC0duQALCcGF4tu/OSR4O
7G0PdeRCDmUHuV7FKA+9hLJ7CMw0kFmDjOghMv028iRAfqq+6Q4/4cxK58tl9UO1vXk3yuTehNjT
A+h2JYHm4GO4R5KWzc3Yt4r6IQsWgCJomPb+aJLpHLyPp0g0+hX1h0NTLIRSE4eE/FGxyJGK1EFD
epFmQKrMcgzTnXKv7KZKdoEL0EcfLfEQs89QHEAl1+7H46mGPPphaembW+aL0Hmn8njGiADrwFS7
ChESmt26VbXVIpVYmDeed7C1y/PRYGUcmVopQ2zXnPGA1+pvln5sb9vbKzVwfT/N4/fwjXbqRINm
S6uB7KgTsuhU7v18L6Sr6ezW/NNrN4s+lATqhPu+y9SIzM18ZkDusJmZdDK39cvHK2dso21T2P4x
c5LKJYcfilOj5K+gs6CGc5ZckhdSrBq235pW4WlVIyIAWMfc2ORCUae025psDUeJ8WTBWj7p24pf
Ks8heihtNWxb9fZ+VPMy1IrRGDcrKqgfmigqpR9D/dC8sUBdVWZcMa0NpTDvqoz9BHitxcEYuKjl
vleU3nunUo2CJGsMluJcSFDjAb4kyXIq6Hv/1bRQf1njceja8ZvB9ZJXVIvOSU6AC4fFCyK7VNy1
dsqIYWWDtqtaQ2GB4PggJn4Yt3FvMt2cUWtCTxZ6/yjKJFuwbOH+4UmZ0gy5pWA4Afr+sIaEHBk2
XjMCIodYzySyEQ0x+U9UWP6uZFRK/k9RCAfJjttIqVQysS+85kL6Yt+SqETWK6xou7M76jMEQdQK
v1bokfAtm6az8pwoxwJye8PMHFxSHOFKSdkGb77OuO57egLnuacIY2XIxP/Sm821fuDnQfwjBHvA
h4U/0tr09hQYhTxk/8974utQe7m+Ymez7Gbt5Ng/spwmpg17qlY5MpbI9zfawxtb2n0s7JMF09y2
bq8ZOw7w/HqNpivKfmK09bu6eN2HOn1cP05Yoibzxc9K3XySoihatNtsb/TNj+4nBkeYspRS/KfT
jz9nsjpJK3t5b/xeNNPIG5GVLbNxoj/f24GHKdrCLLa9vJaNW66HVNKRFHMp7EbX+E1MoX8M+Z9J
qpJ/rbfXEpoBZQv/7kd3PFexGAm/i+QhXcAccnymUd53VqAcsL6wPKzjW0vtv/iCO0mpqD2rqi/V
bODhxtRhIirrfGz/ANfEtfc7x7PLhOFfJAgi+B7tUXjzJY9TImhg9eNaAfhpq0VM43s4fASIKgRv
2lvNOUyRo1IIieJlnXVUKm+HJdwR4hHSgiKmRu3fKMm2klllMYqCVPndJHJ8Lh+bCImkZue4JpCb
XE+AU6VYVCIkWop0ZNflbOEMV/trnIF7IA2lUETm0+m5et1NCcPICAKb26pkKSUqbGUgmP6gCEAQ
5lc/pAl1njMGRjmInu9428yLoQoLZYdXmlMNxM1ryMEna3MJ6JwxQhEiQrUzRfnp5VnioJJLSHFz
ZcZcV5ok+AAh8rhzvLIkCvIxC2/QrIDzUXIH/9XKoFhnmBu0DgkreoKEhGNdqU7y3qdqmVT8Wxnh
QrEdLYeQ4etmij0qs7QO05mCjXhIH10tDVJIRCbDlScIqfGXVL7w3Oqbz5fZZi7bnqEYXe4Skg95
x4KMRdMT9QcsEkQ9R/WzBYGbVEy3jP6kfpxtJSaUZWKQ+03ic+lcyAd45qOluyuHQPFK5E/xaNVz
+xN48vgdO8168ge23rVqtq9eZ27hrCl7MqAMQBri+GGuGxZpfrSEAWVKXH0QHRWdxv/hzelEekuq
ELPsS2PYsctt3ZbXofBfq7x6rbnp8s6mHil1ykiSUd4kQbybsTrjeICzY5zft9ulPdrDixTyCVJ6
DtAzIdUksBB5oY8Q+TuK0QbWepdshVh9BJlVfzCZU0LKhiefLx2a2/5m4763/xDcE+K4IkgIXusU
T6gZ3qoEBeTb/HdZg3pAdVpTAFssF5Wja4/0faapURKbGRf+1NV6Z5bACWNVEVSvHxzEY0F5ql3w
CHxEZpyyiroXaebtQMV0OoLKgWtBwp22nMVfbkKzpXLhwgQDgsGRBreC8bmHCVgqvHUwkRTVMGyH
VgLmfW4lMIJlIEj9CVzF49lKuLCcTuhR2RCmxXSoPLF+hrFkSug6FDqWClItt2TwDtsLpjsyh2eR
JQ8oUr9EeEhBEQHMmxYQ+x/vzYD6+1fN4rImOki7DE7LIip2GlZw9GJ6X5BBWPMcxFkcVV6c3VGR
aJk1RwoVjur3FJPmwS7qr1kvp6kp0veS959E8SOpfBDR40tIbROXMMdEtSlfY+Vzwhh0h0TCAJ52
oJ8dihSrLwgiylrX6oCAy/EZJ57mJWTS10jbeRA4T9sP1/G5yovVRaUdzg3bAX2Q7PRktp5DheF8
4lgYOOkDNS4zV024O4iyZjid0YaAeT4TKJ/cHjtP0Dm2DoUiGONEKf+dnMKIUc1wHWQKEyUmWg5q
w8I6MC6DMUKP8gTtEbZkAdFuWYbW3QpYzZUpDs5wmRkM1GrZ3m3BEpl8cL5QtLl5lQGm/oAFqJ0i
dr8oHpjQb/pZd+diMz5DC3xtTJBL0WrI1qrbtgIz026g/svNAX+pjRmPQ7XizuM5H2ZZmUXxXqCY
GTKa4m+B4WmaevXZqev084yfwoer5Gv7yH41bb8AV3yBW0u2/0fRWDAGBjlO8fkWzprWCYNDgie8
ETHOhArr1Q7RCthvWxIHQ0WcywbJ7cjutLX2xh1pQv/d2gxf1pjFI8ED4xFnbav9BbVYltYKCWh4
P/pfM7Ry3xQeUa2bftw6XV9WNFexCF7iTCVbro6mzWe9PbpCNtoob9xkCvfXHg2IgFaFay6PCgd0
ylajVc5yOzUKy2Cg0Itj1uVqRSNIS62klw+f8whUB7U7Gy9MPxxQBMcsj+f2K4lfCljlQJSGY0qv
mmQlrGS0mPotQBNnDd6ro9NNrvgdFFthBi7v9Q+hO/AP9eE+vZAJbFTS6ofKHH4JZEfRp236X248
A8SQB8yBpCaDxUfpvVS6BrksEg2K1a4553l6Keo2KsLlRKIXiLjiN8bAdoDzVHwo3TOHvcR+xQQW
r3p7nIcSigcvboiIG3ZiZyUrXwmra35ZqXHzAWhjL3HZT1ceK6biMaYZQUj3aEJeDsXaQOGOrw6E
h2Skf4dVlcszFwCTYbdD/eMMdLDkThI6ErZ6U2KOTCVXQPnzoMdaEIW1QeEhhUGkiOWCqj111s6n
Jxts+92Pc5IofokdMZufFiL/4V4TjliZSPpR+ckOg57SgrZw8jS66/HwN0O+5rIZPKxn5iwHBqZN
KrCSctObObtkxZvqo87cQbttnyk20yKpnQT5a6OsAfcn0B0GANyJRe+sLGjuS7ewgEXpgj6YHj5W
dAEoGWRuaDYeqyZ8+8esujYAbjeLPUyGgsQTvfWktoJhGpqpRZeeH1Wks7w126gKVQUnk//QOPwQ
yPQspMeDKgCEVnH/RzGAxsnEeH5KOwFzpip8Ox1qpn3+BcvUWQWoKrhTV0gDEzzGJFeHSeed4q4W
ShLe+F7AZRF4kAYXTebCpTs1jcadpBJqUrsMbK9zfwgM7k+UdndFJTfbg3Z6d3VhfYPYdJHHepPr
Sx8wjCaC6NXSlYrpoNZj6hzibdTKk7au7NuWDT8sOBKB4Ay16CTH8Q3G2/ermEt5JXUGY0UxFTqJ
5Fekc3YYXFjk8cY7BOLWWEXjyHdvPzPR001OqZLbjlZnTHQY6TNM4234oCT0TTVjTf6dT2dmEeuZ
sMNBOK1usBlFO/CCMSVfyVTjb695Srr7q2jk4qQaLp9fBoFMJhfJwbdLcjR6ozr08gUx4RJfkcLp
j3/rTmtiGYyOGj1bLGwrvJ4KiSeBV36R9yi4Cez4qX2wvuesXABt9gne9Df2ovpCX/jntq3Vj1r6
L2QSI3yy2qhOJRPya1WvaSl53rMGsd7h+TL2aeub5B+M1ukZQqyotBWRjMXOTJRb/ME1iwqwMgjy
bQqQNMGPYnGzn8uA6vFIKsyGRxeh0HV5yhbkYua++yiJhuO/+azLHnH2PhbhNsaliaVdEvJvlwAN
IV/BJqGF2FBm33w2V+6u6aaE7dYe9IIQALR2aG0bAdxWCTBTfiHhFpYd5NX2t4oslKmlV5vlhkdG
HgC68Hv+1mWPbDjUgboJIbl5nRNT5roN7vaWJXg+dOSgD3l2WxSPITJByfBn8MtjDPZOucwqi9C5
B9Bq4/7Fo97opKW81knH+9cw7/XPcn6C7BxcPcwiRuHE514zJyEdEvuIxF3FgVMn9/YL3rffgSEd
elb75qizBmEiW2kRQu3/theNKX0fRV6hnd9fBPnHGIwApwtnREM16vMBRd0ktyfSoZUfCStZL8Jm
XCOhkdUtpZxfasM2uqW2YAVNLENZXtj+CMaMh3c83Oznh/05tami/demw14y/hZ9Bnpy57j12VUP
PIYBJdB9jfz5slkgxcJmY7fQ2trA2D8iUk1XEdsXYtDYotRmbV3fotEWbpR91ygpupiDkYk2Lav5
UP8gntIiyHswIiWxYS13SrB60oRfbFYaop+ZZfWmSBZA2nIYlbolBlEQLUa0Gnuyr5W+/jLq7TYg
c78EQf9ytcrgvnxCrZ1hg8mwHUXNuFbU3J6n4PenCfdqBw1bn3VdLhnNPTSGK+7L6fbIn3u6FuwZ
VRByuoiq7fuJ5UCJfwhCN0TP6EF5U/REzauEu19lwoI4gDfZw4gnKCvORm6DWoyK920B9rhsCpLQ
4bnDSYu7abqsKRd98lVwymSlKNlvPqVzYyWcSIpRvzMb4QePbvk60fEhu1Ifr2qfc8fhzXOlFoNm
KcWKxN9tNW2xQCxVi2gHbdqhCzFrBkSAciUhhv2n2ePTF4l23xv0a4aKihCc6U6aZprgYq0EiyWg
WRRsXXM1LLFdYoaX8aMdz37pIkC2MR/Pc/hDqk98RAtsy3tLXEieri7YMxebC5+fddfn9mT+8Kwa
dHfPrP9mRXlWnczvMvBH27RrzugnWc8d4tVQDLyT81PiM2ydnYNigLYO2GGuC78ZRXBmGJkaTaqw
nJQpPDa4faD/p4n7Xpk4M0460b7w8fknaIBWs0TYANoHe1At1nANSQyZT/lEbk+H49Sd1e3kvBzo
IC9PytoZtszXjQ8X8bsPVPHytxjzPTPFSuQ8ZP+fxReY7vF7URb4TDv9OxMjcwfM5azarettOFZg
tkou9VoMosmEvfmC1QPzbRIXvSL/V6A3VrnaAQV/Nsu6HTq997rC/V6d9+lwQsRgAG9stYlRp5Jg
RcOoYNPZtQMyDBrnwQteUaekNQxcKAuhK1J5k+V/vDaj7lVRJCn6I7PTz9We/lvQNPqnXhnSdMCF
tO4zQv3X04Zy8/iQ3ut6YjhyqaQxXybNr3FtfbjI5fmnsiw1qYiMF01DyKhkfj90e+V+ssVlVgc3
Wu4ECRupC+C9W+UzmKq4UxPKWZLmVqxIfrJsk4+J5oOq983huJMgY6RpGswJQUiZyC5TZZaOuBDQ
3sK4HLZU31W7P4dmtUPzmcPxmUmKVF9NQBjNJuRBECwVaD1g45cFmSQixhGoy17HgoJm8kaG7w+8
94qN3mfMTPSoLgScvZKGc2jT9whdPntmBCjrpGodQAb/PZo90KR2FtYzkZB10b0W/iCecJ/zZ9JM
1ojyEqAzelX51XkWsauOuwLmQZhh806L7WvLZWeOikqyrImc2zfT6END+iuBVq/XtiSkJ7s9Dlxf
zZTPjpZmPi+jfgsFMLfYYLva2sNzWQ27Am+gSLuvdMXnNaRdC9C6rTFB1KGaSBEhB4Vkmopm1Hpr
ZaRFDmirujOMOeZG0u++ERtd6T+uo8NyXWqU03y0vPIzcXsF9nLI4n1xBv+bqnT9PtzF2ZL6ezni
Y0VZA89dHoQBUpoyY55e1iqdz9yRBCLnR+Y0hepvnImHhTQ+hrVM84/Z2JRTwZA10lIeyz26iDdN
Bbd2RDAwGLlKCRuTiOBG30nY4MqvgfPoJsStF70+EGpV/uXbT6CPdnHyU3/CW2toTLVk/aSO2Nxc
bTPsnjgnjyGHUMZh2UluAyMAAL0BVV8RVzDF01yuHYeAEKWk2JlcMVXXGoEE/lNkbT4rPwrtAgAs
nCxUC8xaL73macgf+6ppZbaJIyHexTPnKxpRRcYtdcVNK+A5djz4udE8/+GR8FCgKmvr2KHSZUvS
s7NCza/VQKaVOIVDFCavvMAX99MRD2hL0cGFI2a/cKP9f/HLa69QllHtCNn0/Tx8fiGsFFLbz+2Z
q3VmyQ+DpNzIGdC9dW2+eDesgNGWqGyNBVMhHWWeLtF3Tw2B6IVSO3iXkv+B1Pof0ah+Hod1nqWA
ChLcGnsS0Qe1qVl59FFQPW3ZuRKaz33KWzJxXS1R058yc8LCcNKFxG8Sq2rRqRSSGCcH3Je0vKpT
RiZbybw2HsGHwH++qb/YNWB4Q2AZAg0Wt/L11NIiqQj/TMVRnBrJU8x7zaqwzuiH9eo8xWY10lPp
3eLYdlzmn1lr5pzk21oAEio6fcMBRXqYC7gD4NnTmO39oSlB2l/QRxL2FouxS+hkjLK7Hpiesfzu
3FrBHJ89Tgf+BiiCN/5UUVuFJeZX87gohIAghJoRpSO4cPkGGsepn2cLZTmsDywSdfYpdTAAasmL
5D8NF7gO+s5DBDYNUzs/OZfruSOYKKXdt5JDPH/xrbQTAuHgoYKjVFMljLk5ndCiiMBwZqlLWvg+
FjNF58O690fcbvz0x876eVOyDkuMafgkFlp0Ps0EElfODliLpFc0O5AOzFXF0IXksA+6Wg+NrQxv
l/Rodi+XuVu8cRVrku5u1fY49xtHqZ+EdaEURBNon+STmXGbXdyRjs0SVoGOvLPVRkxABMHTF1Sf
sQwbxbeI02ye0HMvHAQGbhkLAfZTNC7/Vsj86VLS1d9BuSdG/grn/E4dVaCHxGfURJ9hdHfF1rFE
BJS4VhAMcmPqoAOq8kFH+dk09jtc6snlMAQ/6rUUS3RmVpxm4q1OsBqWlyq47mCtEJ/QpL3d7Jrr
auYbIDXtlA7w93QvQvQEMJmRYQFnX39qiJRB366EubUYux/gkl04JuNU4exCxyDriELYsCv86XZ8
WSIWb9tz2NsPku3QGK0ZTw5DS/EozxaNd6EMBM44dul+URwmW/ff+NZe73QK4hvDbC4jTd9py9i2
fQqGNeKe80WHbXLUaSaz8tKFpcP62CICuMZFiUTIux31DiiWZvZJQikusAcffm+81RE5W/4Yfrs5
QGveSZZAw1TfVFWCOfnMHMNFpkkUO00APE2TKZx5M+8KRu5g8ZtFlZ+YY7FDXEpt8DEhZzErUgGS
uI8DnceLlpP1dT+mysdW9dvpEvcEPVv2RiwjdA+9oeufdiQJqH02nPFo7bMdsvk9YFYONDxeKSuc
18vOyuIT6DSBuYErZWZio9aRI0vzeIe7e/ypaDRnPLV3H4Y5bzVqixpv1Gq1UUxYFj1zKpoAkRGY
CL04xEF7gOHGdAQAG7foH7Xr9daSi3QVz7w/uWkK7qzh01dtjnBHO5mmrCigYntGvCWZA702bF0O
gUQsoAjv5i7uJaDmTFGRKLoTc3c2NeE32vXCOrwv2Vl0ranAueaxtoRTAxo9HNDRkRO7Tk9U+Z8Z
7tTrDYGmSK0VFkyLDlz3UcCO/PyOeIqdEk+L2JdsflXgrCsWh22xJ8Td6PuECRVi1m8qyD2USNr+
0LQKCx+a3F/qqS8VVgwFLUjPWXdGy95DQ4hmtOJxGchi3AMF3QfQDZCO154rh444fBJCXs5PcmOu
38zGJh/OdSVRoEPY5LK0yzch0D5Xz3d4udm9zTDXbRWbWdUtswGfmZOJA7FE063Nk5KHCoBPvKg4
Z5uzJwWWcFpYHxntwjsL0OUXHQcFQo706jypAkBQD7cSgy7yalbA9KXoCQYPL3QP5UKbdBLcVSlC
rYomWoivJucU3Oh8xEm/rAnWjBzoeojXe02HdmgBgYznqIuwQsGyHXKaFujOYNy6uoSM+mIX9ilZ
D7aQFQgA+AEHcvGwajYSDV38QA+hhX6uEMZrFuQWToNtkMTxbaZXf661W4fM9dQRHve33SWx1fMi
e1Y+7mqy5gc8uHAswIPPYCSIzW/YKY9E42Z7EDTIdBDxKMECNfAwR5zbRqcK1nAnhBq7RFy3SMng
iwc+JPUXqZ3R7VAtDpuavk5KqCSLhgXPef7IsQQPotJ2H+nVRlmWhl0LgUAIZ/CWLGXrMiY5wqL2
Nfo0F4g/RfedORz4NvL2q71Dx7CSChQoRsohbleNB506HcSKHjDowqaO6Ya2gZDjj4OI1WC/U1yT
dP09U4/5lQWwcR6RKx3mD5ed92wodPl8z0QF7Sdizx2qQGofPvaMUoEKzVxJMI4olxwYOfoOzdzJ
74pa0I2H61+quChfGqmWUrAU9kjwZaZjtOd59qyeobXOErJzwvU9FNf7WNe7Vujc5O9GVUn4OMAP
M8kcCmQFqTwc4f3SrvXf9Ou9R7ls3+yw/Z03VvM+DXM1iqYZS3RMDf7bDAs6ppgfKJaX+jsSP4qb
KibJthhsojEM0cMM9UvEOz/RVng5izLxYzyVCsYzfyAFA7JbWXFBMYkkKBynnIt2StOnPsuL112c
uyZ190qfhFa+anv6Gmpw2iQxUVjdMBHEeO8VaATei+P9F29HnL8akK5HDbGYlhlQzc3sgFVJMRgj
yQ700rkWN52vRCP/Zww6pFN/9hWue8nEdUU4ux0CQvYEx7m58h15Hb5jIrGvaabfvwhEVJzk5zYM
JQ4ZftGzlXliq+lP6osxD949XczIHM4uGBmKoHP1NsventZ7DVqxJIJnCFhYXQBPyNUEJecwAPrl
AAh+EaHiz6zDV5AdppKmz/qyR/22eEDBkz+lE33jWWSg1999j+XFZVFSO6PAZkMPCmqvMDjuIlvC
VrRfKQQ5XyCu4vv3AGHgt4ssjBtti7jXUgphZy6LVI4UB/ZmNOz9flrozjhOXMBDAJh9VAflA1IH
1siNG0ECukc6gFnlQG/gZAXAsJsvDL1wrHnBK5vh5+o3lhMpj4/FDy3p30OrPBd1Ynr83cX7taP1
3y50Es3IqNVTQr1hfMMzxf44H4oMFLqNyf/4D6U+8nGmobAmw3N+C6qcjUNphWeWhWou+YluMNYu
9KsD1jK4xSyyUPy5VzRhKdH4HqwcK7XmP2Nt+vLtn4n2nNpZ4uxO0kUrSPINGojzPWxVpWHR4/8L
8citcDyN5RjaOhDUNwZwFAXV2ROH6Sae9h488SJyLzLLWGgUKX6SgOQXBNFVQlGKwkrJyVWI4ONi
J2pynGjdRHM9Kztzr3Bc4jXo4h0kI6cPVkQVXwK65cS5bAVJwlQpjcdOvVGhVPFrtEFTBnAZ8cL8
MqQfZWsBEYlC+nUglFSQ2pesRRZgo+fxS76k515FAO2cCUNUAQGw3MEhdEl8cn9TEjOCVBN6BXHg
TlYsRnhnFf/TRaaOUySsHtLf1LgDBVbkIHCq49fSOVmKVsJG4xAAW/KZBg0yY+nCI/ZisD/xSVpE
Fs2XXAPRJTkhwCt3lq/1z6B25yuyJP5hK+cXMWQfsgE6adja+2BA7SwEI695aO1cdmYEoNgq15P7
+3WWrYyQqW2//iRRlOZfRK4a8G7HRhkdB0H1ztq/Uyn9aWU4zPFM2V2tHGXFyAaJAQMM/F7KPjml
NSxwu05tUY5s+8zNpUqeUYo1QjIUw8apnQFHjtCJ3C/0KljVDlMYkqwOe2B8HExl5ZmMT6/salne
Y4+fqKWsYYx0Ka3hS8dGh6EU8ZbiONJoi7sUFTJnei1fgei5osNGYw/DZvSqNuCtm+WuGdEVFCCj
tUhJJ2B4XO10spewo9v4HrBip9pEzT2iyqpcXM3T5jXTxyG/gukfL29dYz+JKEkSPAE3n+omkvaB
HDcWZJvAsxhUUeEI9LD/wUuBF65oCb/nfqz0JfPOCw/eN57Di1CqgrKKqqKQqCTXJB68TQozBoGc
3oXLdZsLYSnkW2JYRjR4vUoMltULOlUu7gsxKW4DAmrKoQh66hZH/pWUZpVbmL8q+eJ5iL5IEhuH
f/DPW9Q7jIPlGtQbkI1Y0IwuI/94CqbTtbegtTYE91XynOWL0bldLMl3hg0vDd4VYhSJyt1RYFLZ
GM8lGZ/Hd/5tYSTmMNsuGCXfv52KmEspk2LjDtAwt0C7fa4RdJjOXSfPNaZ+C31Iep5tf7wsvahp
Z7vQ6KAIGQL/OAkHIyRNzS0oy7+eKccCsrtlAmrJ5E0uywM3UYWEK0H2ClsgrhfRVztQIzmLXBF7
f2RH4mWa9+hqQYl5YqVcgvZZCjU1IzjMX+jU8qtpMWw/A0srAjQvfcF2ui1rPx86SLDLv7MZlxxb
yf8RhZKWpxiu6lBguUxrY/06MMFplwDZNcPmUpVhVJKqhvn8Cx9BBMOJjFSCwJUQHn4MYXkEuDFD
2WrUKosBRNusYZI1f5IGnLPc4EFn12jaXdcrjUCtkMCuF6xzu3hLR+ZZuyBvEdYaseuszwyjcETL
kybpW6TMnFBTScQrFwSzp10XjjEIKl0k5xQwKUs9PyPQMQMRAElfxyftIaJigVHm7y/e5J7kfpcz
dWNYp1rk8doDxTBZ2QVWKAXbQBdTCIInGEVmOY1MnQh2oY/IhqMZd35Ds1xTOo/9NTXEdlZefety
vs1kgL4oX0zXMP8mJmMnnzfadx7uc+O1yKP8TkyLXjhSP7+W0hcjzC845d9BNc30ah3eP1y+MNby
FxyskiIZ7WLdu51DGNoh4yfZaoNcA6tWJyTUZmg6AKtna/5WZ7Al9NdtXutVOadt9FBW+WGD3FCt
yUwyeBWGmAY3dkqqneVJTwViqnd0IZ3j0r1HHFr2GsR7P2wFwqt3kv4kgCQqNGraeoRciFhO5UY7
eSMhOtVu1Hj8JhSP78GfF+dRxVo7UGjYgKH4z0/in6Fsw4VKwpUpj0ro8QHHohdx6itEqBqoPvIc
kgwWFuG4kkrEl+lI74qrq1eMcMY2307/sYGmYgQ/QGxoV1rJCtLuSe0YRTwXux5YQ/aqE7DDIztX
aNbgTyNZYzP0CBZViQxEHwNdfWWCYmAxQe7oiosBiwOb5+ZypdcpCKp+OAqXBYJAJwIuQkU7ClJR
OA4O0MjnfiruM8apvAq3XmojjvF2kgRdH9gyhncHmYjHIosfLbjPXIdlZRrV8q/RxJFh+JuGDvBL
vUEqHMnlnq7EUInxNWpr/aHnqcCRjCCnu2LkO8Xr/fxrrczaHI0YAkRujYOKlGZwrJe4nT+XePWO
TTphzNG204nS2IGoNKGHSTWW5a/wbQ2+AcdPBM6yBT4xf3FMGZaVAH3+ZQn32w2IjOgsD6INPrcZ
9THFEmRsTpRaRfa8UvBEyYdWbCOmASKiA3GVqxnn62vt6P/N1oSD+zu0/3HYllXgnRae0QqSQSaB
pSR+e46qq7oFTkMMulBOXLLmJAroNZA1kr/8VD0WONfg7GEQOD+W4aS4Zg+0dgYqlWxW0EzE5IK0
0Jqce5omRZN0IyTZIGe5cSsvuE5ffqu9gAGrYinPWLXGSI8x6z7Y40jovDNGdnEyZ4jq3ouPXpAQ
tRxz24E0UFcSi6h7QRbSLmaWVruzaFSqw+Mq92YoJv3+AWpUnle+cN7pzSbKl53Xj/6cpkVZfer8
ZErmMEGmAGbXaNmzljA8uiQKph3UgLBQjTzFJSH6AQeEuYisB7W/GUGZhvZSyf2BJ545Xt06CnFT
zgol9WIbfix9X3ZA8LLO18+NHp4RIQNj8ItuLoJCR6eHWseHdDlkTW2p0Kkqa40DMWVaYO6CQk7U
YtSsidhxKGul5+k/TovIWjCX74xkeFMdRSR35mOOF8cw4McMI71flv3151kyBAUs8AVvub8o5dJN
e9Zz6/qBaN3aBJZh8e2G26rL3h/4SXhvTFcw2Afo2L0ADV0I+9j49UUuXBqPeW2Mj82jeFCc6Png
GkW38Uc7s1H6IReaXus0HqA0sQSkoqXq6w4I+lnQI4rc4LK9/5o/6oIeDUpRQsd/+3/nV2NP6wDH
GjKS1qQIganFys9IiMkclhBU6Et0jGcU9TGABn/gG4GJWYByHXUr5n47bTvd9eQXavSLWqwunwkG
QoTumGeb8Gb7dc1II+kzrN85Y/yTMcKYEoVNomLnjlFA2o3Gak810mKKMWqrXNDWu/vNg0nNJuCj
zEJ/Cgpm9nJ8EPGPV37ITp0NXYfHOQT+87I7f8OupgUBl164TAWoHaQ0Dr2ZfMBHGgC84WDkGRFR
60lrkpvKx5+PxvborsNEJFh/wNeOxaG/LxJL9O71ztnndJ4WdzNi6nPk5El7xud/PSttzI1BdVSd
Ru1ITJ5A6LFCPXBYtFgdH2GLirqfzYY9poIvae5055ow4VKpXMe9Ds2MxyKe197uKFQQqifeBkD2
kN2nTomgnU8BJQQ4rPv9lxSQOsgbU7XZnhuQ0tBMs4SYukZ/uOYgx3v+e8GynK1SSc5LkEQvC6Xm
OSSltlpvwzhj8dRC7AbCMrlULiuqV+a+Nwr7xxxW6hU/9PEpzU/xigP6h7hsK6CZcNwq3q/1Fl9A
xagtaO2HZS5EfP29Im82cvQcSdRZmtHcY85FvoIjIdkyr1jl75+eB/X2rxETf1UGP7qLUVN4hl9S
XBsOr4vJCT+hiZOe5osJ7FNzu7p2zECTvguW6z1yl9YASZo686vkPLr+VMgM/DB2djkfy6Qt/zUI
FbfFuhYEhiMgYYzhcaJ67I5++DMPa9JzS8hfm6kTlTjfe1gB2YCC6TJlYB4oE+ieakqId+Lpp9XC
7KrtitsolvzOmRl4ycuPNJ/eTJ39HPq8XVv1WjtCELk1m0vkrA6hvBHXskrIBC7tD7tMGqkzmBWG
ekXQPjSbDSV4jPFwNV18ys71CmqHya++C70cz4Y5xhA8Nh/dJzZgPzhAVbuhHvHKZEkaOKz3QBAK
kFlkYJ8sa1xDZQTTo3yo2k4xRwAD5MfPdV3lcURT3tJe2qJrspEddAHA9nnr0TN0uBMEPgIe8S80
UTBp6P7Q1omhjIMGSDw/QABzLc86M6knYV5fojDUqqyjOimyxwKgYbp8sMmayYqNVfZ0lF17IPA7
asNVK09vL5WybHFVIVmpENxQwBRBi0/tob8oI/qo+RQ15uHD9jQY0uoQU44OB7CorEasq68Cq4YJ
mASk6XB5kMoZJzuJS3smtj2xbKETE/+bjRmvnTVUfGLYOq0GCcAaIY3pmbfNzf2sJ5uPVoh54f2+
sFMHVJbZ6N2IPwQo+4TT6tOjynhULekajvut2rlwzGYQYwS1cs2Sqb//ttWoRb3vajLt63RHotXk
sG4TqyR5aXQjvrcfIlm/+kcQc5SJdcnxsRFGnVOUvDwoxlGuJ/8NL3a/3PNLZnxXJeSm8Qnulr5C
yZoalisRQ4WVxyiLd5k2RFMBf8AP0LqwIgCziXnlLTFJz5rXSQzRkoslTYDRrUgka0SGIa8o9CzX
XWZmpu0T5+ihKl1dGjt4IQ4nvuglRX3zuX2yasCA8JnLkIpvbtDChoI9aUlKzRIZFFsOwbSYTKDC
fWNKxFCtEdI2iztnbaF9FY/U2WCVra9roZul/hf1gX4l2nL0REwZH6CvUzM9LSvJNux/zl1w5Hpj
vI/aegPL5YF93gTFTJsnX+qdvIFiHe0+RDnPShRRRoxig1grjNurJUAJeF0k9Te+xYI3jXQmgCwX
xG+S5DWAdgdzoh/yZUE4EogRe3+hLt3PNP24zFgZeCW4uaOhmuSpUfp0xSQ8Mxr3bSr6vdtnNQrJ
MJLKKVQRr/lRhTh1W9Q7LtrroctGhOTcitPhLpdM0U5+yLVFVmHup94uzgCz8ZtyWgkIJfiXMBDg
q9ctO1cuwq803EJjEPYr5SkZvXs/+MltVXsvfofXKVE0ZZFxQeUde4AVe0CpVlWZ5QwWaUWicBTa
eDa3jSEQC/igRYM9ZtkM5oaNHVDyofZ2tcQ6V+E99vHKFvV6wZoBUThUf8TjUyk2m4O4kGB3txDp
gacn5KfH5SK9gh9rRrjcBxgcQId5/03gauEq7jp4yI9j57K18Zc/wpsO8t8UgZ+be+8tHF1gulRl
w/QxUqMmM/DYPVIVIwv9qw6/AongEMt/svDpHvUPG7zG/1bn0e46MrGaAPMlUbUIavcSZpWv1j3M
ac95KpCTBfaQr/BkdCT45Hc8C/SQsZciR07EcyA2MqbqGw3Y0rz6tdAnf+QmiprSW8XR94TUH18I
6QMoBaOVJzDgTIr1TToyTM7oKKts+BNlRi6igelt20PKpwqdyzeKzY1pPA31Z1HfjjPio52ai2pp
NBb63pxniUcSj0nOp7UxP722PELg2VZLhEUqiuUzUtDYSB5IWRgYExESIRojafY5xdBuCpZ4014m
W8yk4zmVQXzTunXW5IrS741KFJm6pIO3Q2uUKZr6nAeqcaRhAlIyimupiGFN8KCHMAP0EU9nFvVU
EjHRZeaKNCyCf8Ur22UvS+N5Bt0Zi8ZoIc2lKkXzmoIXmC6uDxOq2Ol2HWQsR/LiwLr3SDpLQH/i
0DGJRtZy5MJ+QHOuFW8Txc2dOE6XxFOq9WeedI2A2PHoiih2FG0mdUaaiGJCq6/DAH9vbB/ctyOS
AntLDfwi8I6l+TP7rTFLbCfffu+GnaX6kzEB+g8ISVp86m3dNjrIKXEodlPN6jjMERps6roaRtZD
F4Tn/2yMhvAfb1O3Wa26ceB8hERPGlozN5IoE2H7q4icYMc5NubvHMxSEGP0h1ukF8ZgA2QfS83N
Z+spr4OGm3k1izT4UovOIoQrWww8hX41uaZPvoAodh4SNxhONbKLjRVA4ydpJaM7aygyR8q2GKNG
iWRiBbj/16nRZecXajRZl3c5qywmhYqb3R4RNS8ocIcHUzWRL7HmBPiKBmLLPoFyUIaOKsIhd3v8
tIM9erH8Xc4Lflfbq3OsvUU1DvsqVVUj1dKer+d+ZBwNHrKa9Uvk2KYSPJKEY1V8fbRzv7LYkY+V
VyJGwcuFNzg8yf7z5cl6Ve/+UpHcNeK0Ii+VFgnVJeC4CivjSgisdMsTl+OTm40Fieb1EbcihRDk
3/hu87ih2TACk+K4mxmt3I1LAaNP88iAzda6k70MOiUGo+3yc7uo6VZ2ISlCStwqKLXlBgbTXGKa
cbWWVrc7qrDW4aJzMgqu6/88+lwzJahPfOjorp2vnefXQMr4/vf1qh+ssnLina0npsq46iJ2jwtj
u0beWBMUAdW1GRfo4xagoU+I8c1vfZzDC7AMeIDBKpbWgmwuvgoXW8pswRQAGfz+VEPM5kdA/4Zq
BhnZus+3NwklUjIBRBro0iM9ti1emwYUqeAtZm7KDWJAG2Hy4nYu0/CkTZs48xSWVXSltdWwx0Nx
d/bSNUegyrMO9Ifzk5y0394oSaRs5x17vOsVj4f+rbB9mG05dOHre5JWWpOyvewTOfxxzzXZJ3TU
NJTR3+Sn2Hzjz9GCTn9fksiSFhRt/8E6Yn+fb/0YY3+rg6Qt/0hjHc07SgeabiGO79ks24ff+Eif
2HtDzuqTVfjFHiFtW1twrPvvJPs9MyY0LlxJqZkjCuMBso9ff73fMggKhqO9Lnd5zBGNzLj6z25o
mshupF+xfPa85CnAs1ZdWP3fjVtk1k4Lj3cMJjfJ7QDMEa3dxe7j1EgHHyrJtPTk53OkKSWv+m1M
InrNwcJMiQ6NGAZr0anQf1zR3r6v1QMEhKU8AZ+1U6rhDUHrKkUHaradSiltM2lWUbVrA+4JPxTQ
Ix/uWPprVFQWsEti2JOEJa38UuB4VeYRJsFTcGSsxG0UIaVpmYIXQFJMwGskewV4LU/JbF3KGWNS
7vosUfH1jqT6XPZwRYbbd23iIQlDfCVIYc4GrsQGTcRhnGxFjGwMYS+AS42pM9EoQ/Of6fOVVarz
moUZXLirnn6FR5/A+fBZ9cT3jAecKKldcCKg8jVB/473efg/4kR8zCd9kQRkZabVdYbnBVyg4cXX
oAJzNVyAD3y6CZxvVpSr5NUGT00iAOoA1W4N9/wc8yGVv98lRZ2fNhh6HICjx87xSWxJqAACZpQo
slvhnQZb4V1aqQEm7diVhl/c+O5t0W4ru4Rp2IcSIXWtDuZpBy9+3FiDrqoEJ+V2MEt4HsJ7Cpkx
zAVmf9g5NQsGSsvO199i0xQVdjE7+qL3p5onZUOm0JoVnTWCsWvot5HPAvADGkUaSmMaOY8ztK5o
I7TWdJkQNRJV1HgzMdnluX+ie4gdfAOpLkuFsjt7m04mV1snHSjSvf96e/ntjJPp4Z/uXoU7zcrA
O7CFrVpJFx2gdWaKjHInm+bTX2OZUAx417jS8HevsXKZpFrYXcKph6S3GdYGnOGtduIyaNd4lako
eDm4LSvyUFjKauyUSkYU/b+kjTHvma4uzRh2cV/dkotlItnGOPwX/FdkB1V+ky8UUnUuLGVB5tp/
PfWuq7rsKPCOsz5vHn8kfXoZPb7LCvSgl7CU+X0kTC0R20LOwuI2vE5erqIcKZgX1gX6++S5foCh
11STli8Q4QKcoPKwvOCWTRBAddtUKrGz7CRiLIVbniPvqab+LlwD1zU6MnSmCQhJLKqEgVetQOtB
En+fSMXR0oZ7Nq+JtRmGoH+RuNx1UvQHrVGIGSUX7zOg4yxa+D8MdJEtUx4mhjYQTtPSQBhyOHBk
uztEKfdRnLXljEOvLjNx581TfyoKvZdbXK4QD57TGCLi5zL2dSqkEEJ27fhiWOyQummGtofVKSlS
/XjUifMJJFlYpEGrD+HQ8vsPod69nu0oaimm2klpiRA+eNY0KLKtxNv0fID0ygjD8jJBfdzFtejH
W/GMk+sFRsWInLVzyKqjSjDF4Eaj+Lx/AbnoGdkkzkk4t9voSXGbEN+T9qqZ4KIX4Krj7Hg1qyJY
wH1LvmVj/NYYTsgFaUwt+sU8f2aL6tfJSasrMlkCQaBNl/iU92o3dQtSuTzmVdZ7ft/eAu/G+U1V
QrUsg9u+l1zpxCAfZ3/NSXP4hmk75XnSZzt95av6E/3L9Y2nHcKFCHPWwXgI2cZgWAKcuBfodfJm
kGbUORm3XW8j1QqVhxrunMBpmgtnrVPjuSTh/Pxb1WdAU9sFcXSkXtdMpgolVDBuABK2vVKov1vx
m90+4fa2BWT1fj63V0DXclT4V73NIdgjDdqdl9fkpRxk7bqypjFmo2yVwN6fRBTxkGcZcn9gW70L
rml6JoJHCQYJaNfc0MsDrJO39eF5SrtUvhJ0pvKg8UMuzVMyNW7BHK8r022ork63xrWOJNw1abQF
l6cCkJ0ScQD0o2PUJSBKpC75ZflXO/VCpfCHCJrLHtJVnDvKvJOVk96pmcYQrMbxGEKz0DVC/LRv
roETn2LpWm6iUA3LimCWGnRL2XdDwIOc3no0xHzQ/6Rmk3AXczP0yOqUuZjWVywyH4bsPSHwuBVr
BaLY5Hi7kmTFa+rqN4UIJxyK0y32W4urVUfLgGXgMP3VO9GkWwrEMVYpgGXUIEx04uCZSs772Sxj
FcY7Xv35nt4wBWIMWbDXSIyXEedczjXHnrqP3FWf0tLryHS3vUDA+i4ITIA3rC7CUsHEtfxsWGCn
SJcHRo6S5NCOyvUMD7rrnqnax729xOm7G5gaKKHWnV4+Ixjys+o6o6ogGqoMnflhOZ6z1rrVC6Xq
kfo3UE15pxe1tWrwzGr9qAxPCV2NnIYEXVIXo19rjgPQ54khwRuSj2x804HcNZoTHfVPt2U7FrYF
6H9dSFzj2WdwCFd7BfCGO/2/udUnNHH/WYtDTjBj1LtCGDuf9yCbr6+zobrV0Ot5ChnalmkJ/mO4
qVHcZVtzrP0xerUyyo27MzyqG0+FFT1j0HkoUVSZDN52WD4Sh4JdN93a78KX1FbJwtjKBspklwlX
hOGYnzfkkuNDgoS0FZUL/pmvX98lFzXFgondCBABaZPUH7AzaM5HFCoBERIGOYbDdSvvzJM8xpqu
EVL90TNEtIZhi/K4k0J1oXE39ghVn6mDhkB06Sf2sETZaLsIT20/1Z1WZcpEn8SjhmVn1PsyDext
c6cI4BWr0pgUgNnrCovtPZhxsPqvCM6M6oqC3tFx8aWonNaUrdaMLYJYe6EnOz4gKq6nYuIM7dL2
kErvJ1x9kRD957rHDPRSyaPYQG6tln5CNR7A0TrS3YfuzbXlPRkipbEJcM7o9Tj32m9EGcVimSki
kT6Q6xyHrvvjCZ8biuL5MUtohqKV4zSLsP2F78zHtMOsmhMhacRhuQQ2NL7IPqUKUSO9YRlpl+3h
9n5dcVHUFusj+Z3pNeTqAKD2NR0xnitzfTy46nG4s7z3Q/GAzVvkVwrX/paHWOg2DZ+Ggim3xrn9
02wgIlUVizPPxnFzlGLVn67LhyU9p87ByZtrsZuMgIGYD8r84Fcb+Yre9dz2u6IxnEyVYzh7JtzI
etMfmwQIeY3JjBzC43ceaNAd4hS95fRhaLV5kJ9B+k+WSDSByeitimCZaIl/CflyE7YjRuTc8H4T
DE11dr+xcOUAMmsD7Iw0w/rgXHAfaQM3fXot8Kh1juyrzR/wer7Wf748qkQW0EvcG20qCG7LROIw
o7F45KmheVHq0nvlTqfrHetoBhmFwux75/d4DcaQO7E4f1nXYzAegvYhpF5qZfTD5+0fwTK6nb++
ULgNp8igH/pKO+JGM8hku/CE31xeS6FOTGUqnAVB/36Gbb/wmym5HE4ryiTr/g5e6h2RWQG1fQoL
OSCO/thWicI6rrkXin4n4jWyjQxsFCRy/ZOCLSohY/AXR3mu+S0JAY4HPHDB8UNB6qJyJU/VUaCw
v3VcdBnFCe/cNXR4pDS6kEp3b6/5YEeHkGHsin74ZgRPLkaGsQoQj5uixsk30Ja3s76i03IR3k3q
wGDv/CfemZKetINz2MZqFqypSeVwFkPd8X4Ja9iL+8P7YLWaP3ETDQ+HQB9udDaE4Q36Xg+qmvgu
An2L4XAzkUa+5WxHGxMzyYovwI4MDB9zLZuLKldhMs9aXAJlQdMLeHCNfXA48tKQRmiTJrbqSWLU
C2LEX4rigb54t10sz8+OlpQTaUAe/ILorNAMVo/E8WGGlsJblZF+yHVfIDDZ5DDpY8eo8GKEpO0f
CTuCurnXatQcmigMqB90yF4EEb0uM7XtVBjlW2CHIE0ejsXJfkJ6qKNJuA/o1OQ2V36JNlxE0d/g
IVpjcSs3/LUUt+8/LrHZo/+JCkq1WlxzHW3vg9LZN30uuwPG46aJDrPjGcRMJhWTFK37TsqBg11/
vLCtsR8+2vn80HZSpHRFSx6o6UotGF/59+LWImL3tqgtp4mYpNxrwbb/mXg2MLQ4JKsuXWwIDrEf
46imkFRcD7XCJvhYALzgxJaL0BdGp0zbdMbZeX8ob+6BXmq9Kj0pRqv5PF0BRawApsDjc4iKu5Rn
qWtgcgo3Cunkcjh8f+1kQMSBT4VcvZuBjhkilZWjYW1jc+2I9avBE/aVcemKro6rhTHxl/6D9I+y
oGHdGCf7KAB7EWfJxRU/zL4Ik6kLWI87tO4QkC4jpa1R6tolzdBnn8o3uivhXygAyJmZGwTa5jgH
FDxLVvJBiJ6LrshQURf/Chgd4s/gUK/qEshHyi2q68Ry/fWciAEBYRx64C9QAUcC2INuJ3BXBvyb
29IhRW3c9N5z2w1H75zKkWl//I7eQrx4JjMlursuHb2JblJoNMLAkUrKyE7gYm+U9x5+marhzXII
rdY7FGtp1yloWxPjSwn2vDhHlwfClTNjqiuRjwFSiKgG/xrEYv4qG0qxZx4wXJ8QpAjNSIHmSg3F
O46uQDa4MxnSI1PlXdeCGkmREHGc7Oi816zy3cocM15ziLM3Vyas9Qd4RZESX3AoP7CbzQEaER3l
zuWbQT1xcwDcT+h3je11fnMppsONAktnc4scRmNl5hbEZ6dZ/orOcDllELWoWtRc7HdeAg7npHzd
MmEvgb6ZTG8TC8sE23Uxpk1bpQ4YBDXv9IqyTgJQSWzMtwRw/cNHQSJ3SqT8MMQS6tmNbcC6CYEI
Mi3nPUA9jIbHwVcwPteS6PaYwqid5pmxSxDrC2taedmuF0DIdGMpsh7NIInXJYEHGjBu0hyG0Lw0
1uLu9j1mD70YAqfeEJmYlgtadchjGvekpz1RnVaqs36GB+PYuqdK+eQlzKk8+BNoeHHCzF7er4Yf
t6gqJwEzBYhnZgv/6LwQmPTD42QYNc9cqgLhQdt/qI6epp8Liz1zpPWsafyrk11hToqb2gLqu1bX
4A1u9N+eA8VWobfSUh8VGujhu1a0Q2BmDzJRBEEXseeejo9RUNKMdlrthrfiR889/RIvt5SUAQ1x
1wHUDaViaA62+51xgJ02Jx3ukhCNVAuiMEjevMDpLUXPtFNnDg81hHNzKIyajAISvQq0ry6n+ax0
v6DBvjZDcyUAmuFL3d5FNkvxhboq7Iu/Zvw9w5e+VUw1Yw7K4WaEnUwUJEDt8N3aakX0K79hbAGW
oE8fcu1U00DR47UkNLwtWC+gwb1Rm5aLQs04Qu7qiarNlsou+Xfbu1+82vuwxhxjRh5Slm4WHkmm
xidOgLLRafgsBM0Y13mnn7ncKAdcq6pm/8xsld40GMSRkG2IZMGHWqyLMBNifsqO7cmIEZMvonDN
FtVgjpB9EqJnNOx2pslfH+QYufz9uyxd34HCFwgBuM98NNyXwnTnlncMxUzqWXbRQzhVSZjOIKn0
LtJVB8f5XJKi9cOqYgFuRnatOe1o9tPpCQeQf0hYJi6OLmmNPLtq90Is1T8aYcUmHfuZRDeQz5Fy
JGbPrmirqhnbx2aedN2YPh7i5FtPU5QXptJ0d6AfsyMoDPS6/vTmEyjyVsObC4k7taaPfmubtPe8
94whOcCpvFz+VzXYjR+JVsMwhGGrRylcmpEzgTQ5Ys/6JrFukQPEzCF3JBZ/O2/5scFdJCfd3VRX
gJOspi8VfxUzocxPnJCk9J36okhm8UifZllitGxCXr4vMCe3UuGgiJAh4QBvpVgWOrEjkXrMX6Qj
4oCXevFQ0VJVtoVX/54978BlrN0CZheHMa18EZkBR6CynWHgP+z0FSUfF3U0yNjL6Qq6gaUHYUNe
GxtkI+14COtmAs6cdWv+4NFfz15yTPIA45814cwrFgEc3aSPehQaCF+gXbNTXgGAxNS11NlVYcas
kzsYP9GSreddITEBQ2xFIJdiMChIz/jQHSi+J2qkfi0KB+1HQM/VimvM4Y4kVhpaOB2wiijUX3aq
UkImUUliRDtScLIfOZofQ8xuUMrgihIaa3D2lNdSM8iSWsRxPusFuopBBzdvhp41wMN/DhKR4rGc
2TzEVR+D+i/N/QMVcrBG0QFM5xahSSsURcplMZ+482afxrFEbiXF6F51EaftnrW509bp1jlIGT1n
HwhgUldpChfctCICPnL9jDFELwBrQN88sBQSHnZQ+7UE6WrmPOCuRYA3HBCzjmWVVZbQTB7zjvEb
rQJrWoSPerM/GgHH/nWvDtxXuBgA3N6ip3MP/kvH3f+p6/UbIjz+n4wWlqQ5/hQ2nOEyvLdbWBsR
nfgX4BT5UPq9OZFLI/qNCN56aoOejgzrpnL4+VVdAS7eQ+GPWugKQFRKlVxvdgsl+SDj1PxcuU2t
yvphShvjGlT9HMnT8L6CFc1M4WBlKPNwF4+PD3PL1nujnbP4AhjASJpQvYgAUImvO6z5dgSnEE6T
s92V9cDs7IhV2a5ausnzHWwRjLQWkoHqk+p5rnNB8ZpDYEwfiXelpH8WUoOD4E9uuaff7YB8MxRQ
BCNk5qB/LoL11rJYabwQ+mk/Bokq8o6d8S+Zpj/6zu1vEfssGcuW2T8vt25wmmWOWoimgj7owwmD
M0uYxaFbXBacKiIgdzfmsA852VFPmTofkn8OCsAqxk9T397sZgqXys8xpdK99oPn2JXH3vxp4jfG
yVFh05YJcAFzg0EirqcloqzRjUn1xbsekJIntPMu6ea0PepJgCTxtBKqJAoxcdREpxQhtz/p/YHE
fPzVM1ztaVJylz5/faY86TqEaFmIrzbAX79kgPPdw2Bs3GahPzPrriz/yoorFgVl0eiCE1CmN4yA
4RLY3k3GDtOJg4mB/+gWAtOPsua9bGfQqJ6Yz4b0xePvaEiM8ZSJtlnLPaWZmASAsnmLVTgi/uhL
0o7NFUOqAL4W2Nr6Tnjj09VbDMTnw+pON8ewyaJ6f9r4Pu+ZpiDrEo82tmhqSL359f1UIzG41PUk
IRMoLdiZIkGFw706sIswuhOw+yuF6rdw/6dwbC1GhKKbbFV9IusAqvDyr1ViL8kmuEbFctlAgVY6
9lysywBrl1TPQrxuBSAu3HTTnu60hIl/Wl6TlgNeRvg2TRM8wFtSykuBMguYeRrg6NzjwIsPYvuq
Be3+B2yPssNgslzoyZ57pRzwK/ZhMRUOFPOBueZBm/UocSXBH9NENyM5uNP3WyHf5SH4TmSDiFK8
PrHoIEODAao1kNRL8ens0jdjy4vy/5ZaV0i+VN/0Muy+rVF+qs2KltUs0hNXCKkG0Gk+nEZfaaIz
hU1AODbWbfrZBan52vpGTNoQIDy3PMkPApcuiEAp8xp/1dopBcxtCsUZQEqfFTYAeLn8f5E1n+WX
Zbn1SZsUGR+DAIxAYn+l/5U/VIMV9jdVkpEt8inHxmNls6OfTwDknlUgvOPgN6+/+Adbu7nLx2CV
N3lcN1c79ps1ArVqZxVmfY6R4ebFIPzm4aQEAYOpJQ9v1/hTmdqKfXahtKksvEcoaf5i9WPqzYMr
LREc6WsRHnXn5rMlGGyRRgOI2V6Hqhj8hJ0X4ueaerGXh/g0o1j7wlW+KiZbFYgOmFLyFDt0ik+p
cGUAtawi8b4TmwivreJVUIVuW6w1lbDply9GnOyb7ygVYitcJYjTLbcaa+U64nkXM4L7KZP4OmVj
aTbN0cRgdtj7FQaCBGGYg14lAWAfwZ2o86rL/rcph3F1RHTLuSpbf1GbMjzUMRQtV+yXebwDRckZ
keX2NQhXV1DGagYugPlH4bjLxYFsa2Gy98kkm+m2KBN2vLrTGEH+ZfJ4oLqlZb2kVUbRhIkK0A79
c1+E+KzRGd7c5jHWF4+hzYPQaBvHO/z+7zSVkXCdthr9s7ByWUPWtq2SLKvt0Q+3HhKzhzL1jSb3
pdDS0BZoD/yQrf46xfCbx/ziG0yULDsw2ndKqMnD1Y4Hf+iWyFY0iG6luceWXY/1muTEEaYN1+Fo
Rz7LFzAD3GDPwH0CCQWjM/cQQjIWu4b4if2ZB88oicCw0fnWEQQyDPjaosBTB83b7EkI2scZc4GQ
8bcFP/tLb5rgOIPRoRK4bezojwgtYec10ZystxfBq5El7Gt9WryrdmgfeznovNr+hNIpmIiTV6tu
EjgRmW2XPPExYCvsxQB1L3Uw78/0IbgosRiVYy74mH7Msmeg4I2nfJiY5rE5b+01mOASXTbD1Hw8
DoJu/8J4z6sLD0+xtPPMlK4zwjQrTOReyjjyxxyKe9trDutMi1KpiaNIujpBd9cI/OOcQiXVEgjr
h+iguKJpVhcPRVeOJasQ2TIBunVw4xJi1ri0DTdXWqqvHSiyL1U5nhNRo4X/efT6QNQTULB5m4A0
dY8hLqnCnln7y29DNJgyct1Qs13A5bfEp+0hzZ5vkUH0ojUD9tzDaMQ4p+or+6/mSDO68qhKnrN/
8gqtNUEyhG7TULBmejrx36mbEcpx4avRpH+YZeUewK26ek9zp5G3elUfW8HvH1/RX89x7LTMZ5N/
JdWsZLAXH/LbjCYaEO8zf0wzS/gsp8WbWNP2ckWoi1VA3T5b69qRiTNjudPwnU8PgrS2xmj8zDCx
0N7AAewTZI09XBkkvlxOo1T2kf0lMfJVuZ6RbW36skRI3lheVZNqMjgucC68Z7RGBo+v/xoG7fBl
4Qi7YkX0BrJ5aQCgTCzr4sWLmEev5AgikxygrvpsauA0AbKgN73I4ZIsK5G4vR8yK0aYpXasl1nU
kFdV74S6r+L+AZARSRdafDebRM7xhn0gukWa8JKtfeqvZovljpujo7NWScPmgGR+Ynaco2QCRrJR
ty9qWlioDXoXlBDfgmUgYWbVKI58UYYOhkxzyJsKI6DmDcsjI978ZTb5kKbEPEli0HuIsg2Ea1AY
shFhk9c4IJeWf1LZ+X1anbgMPALBKhXnZyydjhFimVCE2o2fs6Ek/WBHowx219VCeBCgZG8zGr8t
iBkMYVU8LO5gxWJBCxEhfJOBzbxgZThxmmvYkVgLjDizKOsMKVlZHXmH0OxfNqcLgNgSuo7lJcgM
YhOKA3wlDtTmU7pRZCrIm9T9kNKvp1MFlbvfM7xOoVHFsxtOSGJzbvwkuINloNnLCOEvQETXItzL
yCisn7oe4faHeGAFXi22fb9IQ8TjBCSZGU9yi2eyGysYdcowOJ/ad7c7YU1w0TAEh0AYz5BxBZ7I
Fr4IFPDp6pNCaCuod6H5nKFqPQJBG5BncvTF8oEumDzU04VbNCeanO5oqc6AVOjYrftwt7TKDJPY
W8owvgmDoy4T8KducJJ5igy1SeF5bhOOJdi3jbWbT0Nokq84TBVRJvlv2KXOUV9kcqCnzWP5bkRN
ir0bDk4Cwwr+d/YFYLFnj/yAdUerB/37IZDoDi5nMVN3rZfii4ezsg43FnB18KFbzONS6D+rogpH
VCcJh14szOgaPmcPh2DU7TUsSdHwgGPImXUJ/g2T+fGs9+/Kq9USMFpVgbOU0zsYGXKcWJ8jXcf3
nKnlRQU/bMdapO6dTolM3aC4HNBI0E0u189jwGAFpb9dkcIwa8HQybh+RQ9MugSynk66SzIHrLxW
wo+77d69FO8nK/xHyTIQlZy4Xnaj+Pkk6oHIhQcy0g52MFtJ3aJT1aPP7PtLT7eS92jUHuTXQpey
mnd/xbxxPohxF63RaT06/+iXBQMEPp+uS98gblmKXNcTKnGkC3EBHwcUukgwkWi0EN2GFnEOvb3y
+pBcRPMfkKuroAXUDvA+eGjPFWNZn/K666kIp02D9AO4wttequTBoo6rdZavCUOYR1Q76nvUkzlT
OnSdnsHymCwlW2n5ygEyY9b1uXslToTUrIEkXz9haOUHF/iuZQjaM3KYiY2PxJk8+UyvZKSyIFx8
GKoATNRvSWIMmsRjJsAhvjwXTB3pgq7qVgCSh96URiYjtQnv5HnNOpHMNl26lnofSsAF9uq5ea1z
gmd40WIPNOkt+OQ99Mpco6Jb0in7rObDh8ECqV30Y+HnGBLA7ZKAzWa+248/TjBOjrQRc7n03DDZ
jymK3dYINB2DrlXsQKrSeVxDti1mbRPwtWaUERXA4r3XOkNLT7O+8gTs871h7f7miZc9JMEuN7S7
g6/5qXvj6pJqReCPH5MtyHko8JpAFNooSRugxLspQjMqpzgg3ecK+UhH2GWXx1AGLXCLf5gUXqb+
lguYh/3kCmnH3QtXQF7anbnzrZLLL4XEn9u6DD1VIE6qLoisC1dTvrw8X5WcO1wi0PniOvNcqoko
YeVIZmuOhsQaOfw80qxZsr5rcCEycvDTecIEfWUCvEh7oGm843MvfQdjKGedkCs2Q0UGV9oM1iyO
eyYuS/Q9KpvVxYKyI5FDp1xqHLseZegm08LY3RnoRdQf6yhXn7aOpE+qV5FCpU00fFFYLf1WI8zv
s1l8pH4SzMQ2otKLRJKy+bEtBfN5XMVLDmq0uRN6fLU9BwjlzUqEbY/TLriUvGS49HH/bZm18STN
K5Gob0znkoqzpoNH5rmp03tCQEnz7TWyqONT5RNdxZfonpBYmAX6PuxUX4BJs9VMwK6U2fo4y9Us
/hjcWcPKE3KPhYVTdTruGJ6jpsdBOvFZNE6xJj2JqPFJ4xjapsPsdqAdjBvFloat3m+gSQxh2OqP
lrA0V2vO6iEtqKSw5jUWHkcavoNETA68M5EFo8be8XIq4D+aBAaj3oKxh+OCTQdNdUgqqbDWKYAP
l7cC8bzy58TP6J2VJem6w9bakbet2FwIXAgBNlRU6TOEyuh0AS+kMrpDKQVb0sSRqilVKr5Vqk3k
f4BDbfPUY40uPWNsM26w3UVhhEFgH6SycdM9mrboPevFhGYi2wep0FpTr+FhSo5r4bD2XH2h/Syl
ew7vNOaFaeipvkE17IPM4jt2mulZlOPsz89LSz6uzDT6g7F8k0p39FQkJUXNSrWjD1LUZfsOIlaZ
Am3iNKuH4qQRQiGyJRMoq35ca73QqVvX4mnV8V9T3kkOQ8yKT3EgrQawgMVHLFHhV03d1mCP4U36
0Pqq6eL3iLT09DJf47lGPfRLUgfcnSAjA81invkvPLTTFENUdLW0wSzYih3a6P3rPCrLqcSyB4BZ
k1s8sYPWp0OFFaNCy94cRX39Ru5HhvrI6raubK9vt901qfpmziOtAezx3yAGKr39aO0LhWZ0y3qb
LXEIHmqMNbcJL19HSOSC12xgleLIw8LiLbtjSAtRdb7EOp3UXVyBSObaRWhs5zMwPWsh2lyw5fY3
qhhp0CPfv5bPEVFRUpiQyK/PXWvPb0VTi0NgeU/CzdUrr5yAe7JKDQjmzaUmtsehgp9UkQ8cjylF
IvqktNpfFeZYZOx3NXNwrt3q0CSl+Ji54UPEgyDQTHtBFmmyYbl7WOZ0ToZTG7DdtcvlhJjZeswd
FOsDPRzHMwBpVU/5eeirendXaw8oT0NS0k3xQ8sXSFDrIDT4dM1h6Y3b4+2mEKbsOQDWVHwDKJ0x
oBxO2cO2RXcRHUzSATpcoaopFJPjUSZ6c/CbOszf7jfhnpcKWaAzm07Li3ykj3Aqno4L6b0hx7l9
qKgqALmuYCRuSoemKV4klCpTsi9HDAg6JU+mdhGDz5qFhUt3wSDXbiuWzNivOjzjOsFYM9wMMmwC
cBYNURn8ptDNdo7mF8ZF/jKFUiSzMWUxq6FQiZd2nSy0g7c/wPfLA4K/TtmsYip0Ek6P5S37yOo5
tzbQaTjjbMTiqJNSj/uZNXDMvapHc4FXcb1A0PVa2s4gb5lUkUsbNlmYGmOURKwOD5hhNiPvDq3Y
jrQ1yM/X2uk7gylVe0hu2IhQj173hXvDcbeS2JCZUBKRlD45Pq6fHTVB5QPUX2+qqvUED9xGWaBL
dJjf6mS7AhC4Go8bnbdbVhoC9pRVHAxFFaOq1EOvKK9VaDhIu4BTPJdb5AwpEVJ+oGhzzPLUJuJx
WXYn4rL8S2gvUG3y7K/PCRa7whRNzBBCgSKCpLL7uARIBIM/z0kYLuidk3wodz/b5suf/zUqBeuV
ql9I6jYDs8ooPCMUOVVOGqnZfLJL1xCFWX44f64GRMnhoQtUi6jfyph5uPjJTSI5c7O/nrnXayJ2
9WplKxYnfOfg98b59J2WoBO6wIXlcNxa8jn0a994x+cq4NARHiRIilpNnWV1bx2h1khstAQ5tVw3
y1Pk2YYfwzDz/mmh2VI6k8VmcBfFwztW8KsIA/HC02ogHVAYZnbh8/7zQDtWEdK5OHGLzeBcA3Dg
4pQ7VAiDtoIolf32M1BLY2JA0vowW0q91dN5NhCIJDF0pQ3lVHqxprnftMFphIMwcS3ONDDG3QpI
W8c1dExevd0agQVVIRpL4CSOSI43JD95QjF3Ycgy+t6Sr9Q9lN4nO97zOA36PnCQm5hcKgHDUwrG
UYzvXfB/mh18n+KreQBZY+e2zGqibHRnOWexcAJA1TXPJBH2NpP76IJKfdPQDu9TuLuoeOsim7m2
UwRU91KyL5mSywbNjyqkdjo81rJBN0vA3MYqMJ/gJCi2sUFHHzeoKbHcw/9zbtzeOUXe1lQOIEmh
l7c0jBeS/y29Aqufztq/PXpKiWrexP/tEN9Ne1qqzFyYyVGWpZNXo6EIDUpFu4Oz3aQnDVF8gZMW
zBLoF/MTA2WKwENmGZaiG+Ah9FX1wficgWNnRVsoH5b1uviga0v9PA5Lm3+BqjAYbTp+i+chJyOw
FFamLPANCImxIr0IeomRMKHbxxk5wjlvURNBKwibyPyow1rPkxuYW+LsQG5CUzhkAtCI8Bo/8MP9
epRa+IrGoLXGqju1cNl9dyD1SNvzoaWFfZ9y6WbkOt8ma+l/egVCEhSu6hNPSR8zEcG9VAUGAMoV
G2/LVHwlTdK1OwIlR237h2zeoXAMawBalV5vBqIIYiKND4XqLOvnuBXc/C6f6T9bTFTuOMHD9n8K
y0+E9y2hs2Hl0r1jMq8ja0z9MfgHP7wgFSF5KszgLu4c9gn44pfyJOm2eopvYpC4jRPds1famHa6
jiyiqcYEpccnNa8MaS6XtotpBLSP5iL8mKan36S21f3tiyLmETnqcMzbC+xrNmINJ2ACxSq7zWve
iecKkae6lDSkFArGtRNadTTud9k4XIpYDA8vQ3dFqxB/+7x+WxLUjrhUB3VETcoKcRbMjw4MThAx
lb8hBSXTh5PRQ1TYq9LMwFd42FlLUIShYZxRYdb/1Daiill8CQATehQUJkOvubkxHNqxxX3hbxiO
/LaA26/coSLKo8z6RVqSDm8aA+iwI7YY12iyYoXO5ADvYNwrsfkHwYeLTDR0S4uKMdNqJgJ0yHgQ
DbRfZHCSK9MKB6KHq/3YEjNOXWQBvq/fp6Ctk0KCu4X2V1UXeY2gLIqQivmDJbnjYkQSPH39BamM
RWrdACnW/PUu7wUxNX8y+QEciafeyKtnIGyweDCWkNtAXfqu8yjq02lSbsMnyzZa4gyNgvtgrNcj
ourqCO1INa++tV9dkjz8GB466p1UEFc37HT1CVHUzMo1fnflKxb+F4Z/zpBDQ9JVe2ArdPPatDSK
jzBIr5vud+//5p83uqMgoweJHMeqCBw3eZQppEgvgHU+uk3K/bZxARPcRrmY86qTxcZWuUwoC5zB
AEXTGTAWDCG8WFeANJsY3OXR7CQMldY5cwahaB+YF4aUBX2yvPO2VRSmqBstzu6/zSfkDbgaXq4d
8OqYqb1fod3uqLiYQLrpgFNz7x6vufvA9WktDakEXZ+PcOj6b4/SpIfrChXuskIeBPIrjsDlaHds
ruc04NBQNbD7D14CaxHmLk1ktgU5xs4H3YWqRdIOYjY2jQvwLQ7z9kgcdemMzdy1oCiwPPrDDsUZ
xPqWcDFw3Hqpzuw6P2+H8zF0VFMzRtul6y3/CP9ldtnLoyI2nxlZvdzGkTTMADpWSt1UvvOdrbtX
hsW2ydZO9VkBBn/vC/JrDTeyRRzZwaBFm+z2QRcGpfsNcQfB49CuypZXFwOylTWzph3vG3dw0J43
qIhSFlGFPa/YI4TR0tivEMqrGpfs1eXica49reh32eBYKVP8cQnqOfu7K96pe5g3qGrRmsYtMIV1
GdIpSn9MMZO6dN+nCtVu8mWSLyT0vdVdkLKmpS5QRumaoP6G8j+E86k2WOZCMp7FNKUHXVINlTwn
rg9E3l+iozhb7LlyQOFpvll+AwYymScvalU5PkF3njuIvRGBGrBNi9sUlBrUiTvv1HWxUnhfhLCg
m7559XvmRy4gKv+BYM0DoAsACtxefjOPoNTJOyy0R10XvicIOVDnpcd00qm15CCc7R8528zNuyDF
Jet2ejpIoJDBP+Tnc3FMQ0tRyC7nUVRNVAnhcKs3ZAg4UuwPTJnU0rer3p6iBce1OVMey94nItI4
FFGRlR+4PNdz+r96rRYK23rXZbFXxQCO1EBNzh1pljL9vI1TVp2Wo9X0V/wWRxG07baW4qYIFCaH
6qYPVAcXxklBT/GfGxVD9UfFzMeHIjSiOKY0g8gBoSYqxBTN4GHUYuraO6Hjo5iD+AEZJxatHfUU
fR1e3D2RxlVad6po69h9/nwgriHFHDPw1EaCernQIH3QlkexjDQwZZyo720SgeLP+2iX5fqqaY6t
9GEe6lyoe8pWTkpkxsWc7T1La3V4YqcvUBO5QveEQO3SMNnnsyZX2kryEhJz5251dTHrruaLzWn8
ZLSuaGFkfIPgzmMtXiAKJTqKltim51Lw1zqRLNu2g+zlVi6Rqm9DmJEGS5iAAJoX39nktFBmEZA5
yw/+d0t6yyKA7rug3Hm7ZfKUMOcOijVPbM/yKEIDPPqooiA36bPy+0DfFeH8qDSid+/rOy+l3xtb
0dsLX28O3Ap0YIWjB6ByOu37wv98YUMecC/aYyl29XOGTgNMGaK3cYKNiL/g79k9nO7DAKaYS1iL
jDQJNSM8Qnuo93/z1DsqA7p1zN0iIZj2FxOjaq9dMXOSZRLy96/7JEEcTWZSC4Uwadhfk1ttdOeL
hBYfjjyR1UKGV22xadLU1C+JFccWuWBa3KZY/+/9sIg+Q82Ojc5EK61ReTPjh07pZ4hSroWWOpoW
71euvakAErbatHJFaoUcinoQlvCXPoydqRUAq7XtxNk3Slh4bgVKznOFZXencd8Q/ot3ZvV+EEKL
tHozZft1HzcIEQLqNmpptamn3I7HdVsnIMmE64IqGMNH79N4av1BFSflC1Xcbu6+XQ9gp4iXJbVU
MQJ80ENO90KAb/jHaaWbiBYtWGBomXO+8JklZU3Bqfo1Fr5XlBng/B5au7US8WKhkvRT3o1X0OGF
qbP8/tea4SVDOthslDFdmnksGdMJEoZSQBbGJmwnUQg/fjZyDkgQmJeKTjh4T0k1om2aZHtZOW0o
uH2dFNWrlQenFNVETT9HF0Psjsc023O29GPHjaL3k9dA/qn/oQ2WO3ylts9h00REyEY4vywXVGO/
M2y/WLlXnxmEIpwTQxRB73sKDImik2WLB48sD78xxTclSakCWTf7ABAG+kfVtNNnu7dUgsjoR8LT
xbn+l4PoEUs1LoU2t0b/mlgA8mlt/k7rcIcHtvGqnLBU42IAh5Gmw6UojT2WAdnnFJnxOXBGk271
dfjP8a+xWpqJZc7FjVocs6X2Gki+gUsdREgoxjWQU+ZeGpu1DePr7bn09ZnaidKVhkmoTbU5TqmM
VeQusVh6LdskfCXAUmPRPbPfzSzEzyvQyGTfMTj990oylf4JHrpNCssfxMaLyGZ6zONGr/cex0FZ
Y8Yw89kzfA3BfjzOIy3bFTO9dRF/oJuPPvupYdyNfiqLr9k/r1WFryMFhVoFomPn3mVKn9FL7uiX
FVPUR4pynWNPjrLOxDqwu9DfxtIU6JgIKwwqmDe/cXFf3n+zJb0+wYyedk+kvV+4W4mISOhaaP59
S/NAYKSjzUX6sRDGsfMal2TXUYtBXxD2UEA+JEMmgUBcIhz4Bps0g8ruLwHuxf3qE19DX4BgqP2x
/essIACMS85L4G3qKcSNnjE2SH06IOhEzgWLMd9rbffeQ5fE0Jb5RWVdiGKyyVXw/40uaZFE+RCH
2e3r3Ll5wNbP8hlBKZVAgcEodqi4/a8JDFKRUXPeEg/OxbIqBjBvREwauAbpWC38sHlVBVQ4oxit
HI5OVc8t+p3deQKcjxFC6n3UU9Q70QtRuGXC0GMyVe3AfK1Eo8XD1J8OfWC2EXaHrbNHLazpHRKV
sWmsx+GnXQyyPlxNHt9rlchcCNOnhzwZx+pDicLM3uvp3N9Z34znAYGSoJbTVudzTiFysqQ87mRh
4g7c6IOcDSfAVlWZO1Lra2mG5BEU3pPZAiegcZ0IVHyE05CRqhlRjZvbD66czJvSK/24v6Bo00Ra
lRRPDdUt3BAtEFhAhgaIsQE7qXX7K6XdVa4cXcbaY0d6h/DSNqe1eNdrTDEjiWw5CG6SJJ1s0FTE
rQAiuUSzsbGg7SFibHk8GmdwXyyO6MMSz6pUhjhZ9+4JQLKXgPBvxMJHNTl+x6lPbw+3WCqBgikE
vhYkCUY2ZsvnEG9Az9BdN4XMaBddxQWJGd6Pi6oedGgwJz8CTQjvuvsMjG2Kzpsm8GiwPwDbMhdd
J2+MdlgYBKyAMHiRQmT9eNpR6LjCz06G0MthKHSUS4i8YsyymCarxegLSnEfcdPeOrHF9sHHfoAY
NlIKgvTZ93o5znWuA3w8u7UBRJQsCjTOTRUCgZvRJ+AyebMJj3NBhRCcQY0jSEzIppG03ctGoXkL
tAC1uj052Xl6rOF/lCUly7Pu7MRsxs66/Tdkz3X4kOUyfFaHS8h5ffkQGyr2ZzeHIzJ1uW8hujnY
POBqaTioPfq125iobwN7cWXBaJPCx2/PIQCz6u7F02eMc/R+1vmfnyZWtR+G/2jEfoSvca3ImiOQ
OoL9pZCxkQ1A035iP3j+hqX+zK8VDyfhdxc+cPW26ldrtqGexVLNY0LXV7PMScak61/iZQEbQtCF
ZkhOxKO4nV+nZ5l4oPjf6KvcqcsK/nVeLcqSW0RgIhb9RjXRvdBrMoKBfYNw88ZhghOKAoe/jQYb
pe9KYwwNagMT0NCaG254s9lVpQzkQMgACYDpfR0G8pVrr3k/FJBpjY7AGeHD8FDqbhMOZ7j5Y7u9
VEERtDJqQ0km/egxVe5NDr8D3Y1L7pUblgy7d+bYXgMT/hPb90p0En5cy4JjsPQP3X1S6qE5lUNz
LMWyn8fT1z+vCP9WthqIgN7oR2ATzsRyNZcMIPYb72jt9uIhZz+Hy0J/MJ9KJkopVVsJBHUgYCYK
K/w54D16nNrMJznt78Kzs4XxdUOOgzJ8CdTUmdU+tX5RxFBVPFjmT0LEYGGFw+fRasKnjEoPict+
qX5HXOTjfZ5XplzDFknHc/kDyLAMdPVmfffRMNfP5kUDXI1CE/Kq+szSrbNrr2G7aPvpKSY3ncI2
LDOqMrBbG9vt2jpKc30ctGroWVDSmPmAAVBBhEEeoFBe6SNIdJBA6lZmm3bg+IUhUtETt8l/0twd
C6dUYiwbBucqn1r6CghPgJ2wkBk8RBUxeCT0IBEYgW1MI+9xkA4Ty9ZGCfm3IfYAZ+Cjq3uirjN1
7N8/tArn+7F14myX7I6ogKFIjcVBn8+jR+wwUC4tHyHa8ImH4bB4foFp7lIDPZyvMjfgYBRP491T
ioLbJBdd8mBvQ4HDFndIMO61uTl3LzF2ARFNZjQKv+bKxDKxSfI8Bl4BsdhBnb2PtAd9c88dJwDB
rlZm0aSxa9XDycpg6lP48BrEgvQA8UOA9sWHZopMHmr7T2rLseFcbQp1NVld4sKMAk92hYzBY8/S
SC66RkSWPrmDGMrdqvFpR76wUvQUUXfl5g0ltRQ9AcP7ePQBfmUc27E5pfLGRodEghsOiwWuJXw5
J0Hd677JBV+p8iDl+Yyv+M8a1OEUyXP46kCjjWeFv/bpQPnwxLOHUhMPK4JgtU4aRFMH4Cspl5jX
aUpGhA3CEWjRaTTMnWu19dt+ASilD3+AmV2iAhUTD6Cy0akZZP8k1wkSwJQSAnd1iqNH9HRTKQ2Y
U8P6D92JFAKROAgMKbwNxUc1sFFB2veWw8NBRgduBfRy1r185xZ+Ekhaj1h62xp/Mh5UHC8C1pfk
QpLqwbA02TrCcKnyxi8yYyjfbc+YnFCqCsSxScHI6D3tpN5aQErA/58LoNzkzRtnQiyWr2m8Rvp/
vX4u99sURcQ2b6d4A5p9xsTIlXwTkeSN9T2w15Wj9ojJnyeZPQb3FOcncAjhC0VD9ITkZOBHjlsr
lmbe9qmYPl9EhxefuAqbaBDx3tJGaf2U8EgV2QfYdsPg0E+H+2bV2fIyGIcI81QR/xtXtlxFpRUp
+ukV6n4aYTwqNm4CTY9V0LrKARZ3rfGEyJYEdIdrqb/ysNEn3xcKFB3XeSWePUZJE4gxRjXOnMw+
T53IR128HVXSFhfVDOeLAh9adPLj/xYcIH9lMfkz8NmUOKV+eSjxehiGqc7H6FcW66wiXdLwDx8x
scpXOExcrQK3xB9rwDyWiOXNlWQH/kYcji2pe/NBbzzhEdERued89j3vNFVPTuFuQt7b1iezifnF
iUKq9qKPP74ScAt4IbaPx6pvQHaT1MxAh1ly+MpiwsT+QKKaxUkUtvzA5gdO1OSdr58582UvwIsY
ZOLq6tPFFNXikF/ovSr/8i4lAgu1FuSzAUm+tLk/2PHiOMED/tHALV4RDe6wLv18DtPUK+/XFfgx
gWTCPuG+MyNVon0FOy+Kp5zKo7wPidIm1zJ0DDPrkDXBlbauz7F6p3DFhr4YXyog4LGAqrJomuIB
pkwYnjJSY/saMNQkbQl64b0QTvQJV10wfCMyPBktfQNIbYCNGTuYTyvT5jbsTZKl3a/UpMsqB9U5
GAUyJm3Bn6Tzwi3IH/ZHAdWRS66cgF7WvXnBE27jM+Ra0jxtbWMxdYL+rkfWp4ABj05FxLhhLPBc
TfxMnp/d4QIevHPoKKDje7qr1r5Ftgv+qQWmeNq0DxLfziR8nbl+07PAq/PJIVuNEkhGLm8p93GG
0igvN2OmH01xelovp9EvCR32auXEJPpIkxDMksPyjaxYJY6Wkr3lCKQu2kpaq8Wet5+OyNxIwkuf
eauO9LbXlWRrhazosV+vW3EAbAS/k15N4aA5RJKNL/ddfl8gbOBdVAq2Z9gqIGbhESwe2HcBPhEM
rRN03sKRXeWFldd8YmbBvBGrKaXmplAUMZ+UIX0Yn5LvWK5n0uDvy1amLCHMCe2YDKApsrLVcsxP
0ynWGN3NbYUy7U8YLuYXlJriKUSREFQ3lMGk+28w2xX0ZCpY/xcenGqI00c+RNHFBvSgehUakDmt
TzLiEAGV9QPvmTJEMO7tTLwUzmQGqweUuNxeaQOljbfQzCAVTC5CBzsDr5Yhev4HSKFfxxeL0CdP
p67Dq7pcIegEQ5OUSuEidIr0Tms6YpYyYM6mVj6pMbRVeAHzpnNA+jIytm0B0936qyH5hbVFWwjn
nYSU8kbTxRdBk4tYJ0dewNvaHBQA5BdB1RFCkVVtaaCrQ4URmaUTWXrnugZ9tmM3Tpn/TtPGcVQc
wmpgujzEtqA//ttVtnebw6jlfQ6VX9xNv9bL129T1YogMq/N/N9iSZGEmesyBVB6txF28GJJXGEt
T4hsYJUzpQ/A4NXffa3L/tivLqSxdpszkHOCIOh6C6DADV9gIhVWseUXHqACRqsYtPkM9HwasFWi
S9+BCGnkAzoe66cfFhWE3b6uqkhj4giPnAYCwRPqm4jTFpSUgmZZNzwV76mEQh/FRMoK3TEsfa5x
XTPCNe+HqgE4m6YxxFWMr/aMRqmgTxyctiGxb6kLh2X6gNTiwK0yJEa+bPe0J5iNY5gLdZIa+vhp
Jt5x1a48rnQJkgPtmcNy+ktp8rQBzCl051ifeCQlX7ZVk0InMtOxvHN0i+UbZo1RHjGgkjz0BdIc
Iv17BlF/vimhOi3XEfvJL21ZmIfNl4XDLxzxZY920JGkrQPOl6BkXU3y31tYcXdNGivTDALcVsza
kRArprSP2HveEo6tZnSt4482g+hNHZLgXjtNkc2MT2wQ6eQVLNT4RmwZa7wjwiL+41VohnRMCpdY
Z8uKkItqqtn7YiSL3J298i3Ba1RxiQTDOzVIkbxVJs1nqltSFV85AVLqfHpSyzqHSVOXrz85YcHf
davhT/rEqrJQ13bef9zYKJaFA8Cy9XgCzxf1rqomzbIfDCEnTZeDhS/2xYoV1gO7ULzWfjtGpvFp
OX5H70LemqBaQ7+xveDj6fcTYpHIu22ZKIaci/Z/oHoFOAqAFM03DPL1qZcj2TMjVdpIR/vS16XE
fLrYM/rJNHL9BD7RSz1yT8iPN4ixnRJQpWiWburmUWghTBS176D5H6mCenjRVWI8MlNw1MFWEQyt
5UwCiZhzzXJIY2YcCKL1QSHW6EZcp7xNJb/yk72Xi5KWCb++zp7amo8rBT5pthRguRMZezExukBe
fsoAi7gvVw4wSGH0iophzu2Hu3dROI6h4LJzmApv947ajFK4s0mOaVyhXm+f9rKBTsZ3qivwwW4G
OzAlReudd6EbzPhog5OhlXmkLg62XHaYJG+fEGfZpA3FdSgbfaYHM89iTkHIHOZy+PIoyh9KhtoF
PrQhaCXxct88SKSuIO3OOnU8ACljMrx4rtBqA2LaSfk0+zav0QY8Aeq51yz7R+XOoqH3rL/vtfvs
EL3TbwrYMVyZyZX6cUidScDdEGkdNxHktJeYNJgzV+KWXq9h+QZJaALrSp+bLrzUvuCExtRle6MQ
KouO58QAJCtIMzivaO3g7hsqEAlbkpmjbaxf6/hc8dRrtelzMdVwG3SUIQIaULdaWb9uaZlXla7u
rHcDzQw9EHkgZQDzdVDGFzbDEWv+ZsrKT2ecBO2Xj34Sp8t7X3k12zWwqZeeq6o06S0mtCd9jdpd
i6sfPgVWPe+7ed0XT/f9qLYdf//GR+ksXFhmZb92e5YtwZoR7RTYEFwvQ333uqhx9BBBvslAA3ae
LW0U/Pl7lBkqlQt4jiWYPUV1WADff/yY3f8X1ZPaDRiMEWqfqY1nUHv3h3psPd45JQvuQm6kU+vA
qo6pqrwaiHaCM8x+AXdTk4aWtMdShJjaV3BJUS6dkCwUoFTMqL4sbm07AsXwGmlJDRPChLOBv40v
4lxpGXi89uGnDBx/Fxrq6jxOuuKXb7ujCJc/q9fwYpqFOVreCdzUStsQNdjCM0QoGNHEOfPorKX7
Tyg53ih25lU5PqKDkqSf30chBEdhLPHVQkquphNTDFUhh04NgvR4AFBW+mHz8/TobfZ/cfec2y72
wuu7eU+eysWa8IFzIwHgxgoJKFH0EzfUKFjEcy4rzPVnNmVvkSXi8llMXeIkDglsRV6abBcjYH2v
mm9GoNgeuxW6PLTcOHmO3eiBUbES6bvUCf72hT3u2gak0DnglhZOdU4Z0J/4bZafTuQoAMHKnC7l
9ywrCSJucTGq3RWjbD0MPAES9SG4nMAuoGQ+8zIekSqoRT3I+evyCKDpbuZiw6N73Rf4JkzX7qqi
JGnhcaRtcUqNwOcPnc3/XjLprt3XoQ/3RhnM3mPdivVIlj9Xg6wr1C5lZQauvTMtAvFsqOgK73G/
MoKmUWx3e5tjs5Iqd/r65LhzzjuK4Pj2Dq47x4NWs6RdUPHIL97JixuCWoaaDnkEfWSr0qVGT1mG
5/n3fhDaOM/pPcGN10WKVA6pbIic7HNh9eec5bSaahy2j0jfGO9DHK4GdklD4qzSg6nFnkfdDaQK
Fs6H6JMVJOOCjWTQYaYxSOd0mGJaGQ+zW00e7EtbUk1ID+ydjxwuVBHM3cZ+nbm/EfLeEu5YbLUN
NzRte4ptq1ctkBrJZRPGGQc1xAQ7PEYJs5HV1PNBkLz/QLBu8LEZePilpEFI37zIP07dHGY6jn+J
/5JloX8Zb6Gl3dca0YEcG9baQikiJlVn0kuIFx8NgOJEilcyAJAaejBSbUOr2xql9d5HLNE6FfB/
5IXCPKfFmja6vZM+2yHpu/32Cvb2QqVGAbhi6rwuiN58HbOXKAdIWCcb1kzzJqR2eRx5cwMAIT6u
OoElElA+2GYCNn1HsuJ3wTX+Wj2TkStEjtPz4t0W3lFiXnohAdm8+KXmtvlVrkOdR9KmuatsjhFc
ws1BGNGN/i+jPGG2BPalhNyuuhKM6RjYIowmiK2XCLA+da+Geta3T7ckgcliEV4pIjf7U/ZXSJND
urILyARSwXydVfYaaNHgTTPaFfp3xTyRIj1/vpMmXgVroxMFoPH65LEPyFQ52FZ7xvZQGy2ToeC+
GJ82KzGIu7HP19O7mNSq3Obg7EOWwwRroYit4fOP8t0sEG96jk7MOMJ5M2+xmTQcDbNdxb67k8UE
p0jPXSXaA4NTj1P4qxG7ooalOrC0Qqk577E6K0tr1lgO/TSdFZTzY9ax7GUe0UTOO9Cf0dq7nem7
3dDWo9XKwK6wfRNoPMN+CAHlYjAhveFUxPzrBrkxjKPQni7q2yskXwascQF1OueD5mOHswjm9TLU
n2Z++1wnqSHcM/nP7OVmSfkeQUF4eOfuqmwjtI4bQ6auJqZ9oDzIOtSdYKH5lQ3l8Ik66erjrR2M
g5VUqywOr0wiCDvparMibOYd1dbuNkE31Z38/wrVjg21X1gpzvGSUT+ztHRi+yI3iwwQzPU+uCrW
OP0SAE4cx8HV9wFUDwxYKfasKEY8bxns5g/nNKUV5u/3U6+31gY5ERwRKh0U4SSxRh0VR7S90jWk
S7ypb9nlbL5n7lf+jjFqDFeiG1ey27Q1uPi1K7rWcGBXy2Jvy7RAOuwWgBzRX7xtvSfa/jQcJ5w9
y+Wn9um4RwbJsnwxsEdYzlVSKLdafbY0BAzTZAmsH9+/WgrHJqTPGHmbMrj7Iurn2gF0/tKR+voT
plfhyF8CwrlWGjt0onZ8rZCzFA4ToD3dBGVJvdmWfHdf6ZmB+37x8c614BIz63Ytc0u6PBTLy3BB
ZRvVObJokDkS3DXkZS3psVUNnSf1xF4DNWQdpeLOiKFqaUDMFqodq6a5Q5vTHQHrYg5WfViTFqz2
UPblRfxcZeTVFKhD6rL0Ef8DadjOAPgSI0OV3sslN6DeRtoubspB2GaaiZIaGfyv1Nwbn7S9Wsxx
5xe0kpQ17HkpTkS1QiLF66akp3VDBBonWKcXK363R5a7nxip+IZUjuN+rpBiZnMSiPbsTcwOZWiN
0OjElspBJJcC78N3hHDEozRFjFKkA79CN68g80gg71VRZDpmw8YvWciESlFUlz9UpDcrTqmRIBrm
ASXs/hlazR83IcgjgwSs7rGAV2uL78Ubp7a2SQ8XLNHqV9ZjbuD6Vn2ZUBh969Q81tjxjFyfng9A
NEMVXH+FC2H3FYdzOZv+GnaMYiDv2ZJwFb/BeRY53woqCs5oL6DI4FFL+EUi8Dw/4qRjUWAUDoT7
u1Op2xw/0DjYc8hwcVIdo7CcAQ+BEUrCxovMaDpqncD215m7Alzys/kPDzuNn/ntk2dZ3JhbCui+
9bcJEti6TlFhVtGwQExQ8jZ0ces1rN6S21TkXMiMYywi+QrJLK3CItOX0Rlz8M0uu4yt+ZH1k4Ls
8TINz4yHzErS65b3dCfAXqg77RELl7wdwkbhKWOtj4hYLUSV/PKnBOhc+XhxhlvEG+QCsLNl7/hx
AJHc+ujyN159q2/Ig2IkW1t/X3ldUtn926e7LQABGkXh8BT9sTqJHxStGFWVzNxNkymK6AeifAsM
zXa9DPWtr18EztgBrXQ7CQb0sTmOpnsds/9pP4Wfeu/yj89cRvrlIDkth3dAo3piklDhYIu44Uxm
FsGt2jx6du/dfNFl7yHjO27Vb8M5F0JpdHWdu4WZAkJDS2SUgd95/ZwjVwn90C5zzvsFOhjJdGm0
xmQDHEXmbq4vK51c6genCToNtT5OAL3Za1sgwMjvlyPkzR8CKtpqZUaVh57U54kqP6aR/3pUaW53
ke48mhV5XFxWyMiVLStfRkV1BK8XKSKeZ9AvzVF7PmMq0aPST2xVPdDOmF3W3QpDpR7DMIE89wwa
KvOGIMOzxkWtUnv30QtJUfHux8i3KcD3ObKUaQK7nf39Q/8+Rocx3fhBoYqJVtBv4rqy6I5a6YXv
ZSGIUgwAOb5GgBoogFdiyYkfsU9dDgRTW5rSPtYVgaa5mAKQyRrKBOSPGKs6eAfXoX8rMBcneovr
e7KIT6DBcjuaGm820PhA1IthLTyMzx4FL0wY76uwEtfBv0ARvth2GkwEGR8HIBdpJy4MNBCLxVxp
V5cSos6bKCeniudb/Qr5/PVHiH+FqisvNPr8YJvS8U6b8GKpWninfjbY1xv9oIS8uD4e1BiWpGVX
ENLomriogVbpWjLYU7P4+itEHh/GXpYb65sazVwb9CWLLwpnZjKom5HoojAfekHkKYGfFl6wUoBP
zuXthyZp1vYL5V09Zs/13IJppQJPf0h9t6PNoQ5PANyG+mXfYotv+os8gWriqdh4yfuUUCBHu5be
kkXjStFEdToYC9Yu8RQvGSMrktECxtzc6VzkdJLZ3aad0mPmpFPfQD7lqUTeV47Mdr9gdsb+laOT
1NPIMcYeOC4TyUJrJaLf461PvfDLr4+xP+16k+oZfEzN9+orBQ82fLqfIms33tFDAD2HJ6n53iBx
idT/yGx/ueK7lqQQmjtkjLiJsuXGRVaoFqYwAqWoydIHx3xisXRnyi0BPAqsDBXrqe9q54bpkTMI
iIQLY/fxjDud0A45nc6HMa1dXWQaZOm6CB7urErGrqNmCG2H8gxN/WqQjt2T8BVaM8RzKOSVB7mP
viXXP2KvirPquZwRnBfp8uLRqaJrdcaPtw/CCLj+9thEdrnvb2S51eiDlEvkLDRYoD/KPNJbRzhn
fH3eyT8igU9vF9c5/pkjPJD/DTY1Ja2Q9/LZu+vszAn9eIWKOBHB22ePFb6GmmaXQyvsTrhhADPF
3sq9d02elu6GIffq9ZXjQOW2tWGAMaLOSD30gzYW9dpSUkkNEXOgJBVl6fkb1gsabbDLEWaTzHyo
GKJAoUmb8T97Ek9X9+nSnflwaw9Bm0AjTMwVJ1yLXxW+Q9gRBwitjbbnHiN8WLTald5quWI5H4cz
dooViY9tnGWEYWy+PgzweIHGKslp6BSIwApgVSQssHBWI0HQpcRP26jlFYYCtRz4md5iFIQl5uLH
yltrSIBZUwEEAdYq3Wo8yvPnS7bWoVR5+rYMDyxlMFpK9FZG2mCHipTVshsE2mK8zS0TtozkQVLm
BlYve4+YdJd1+AqeCpCpRhEWPG6zVO0OfoY6zWQfCOKyBEE87VyDuPxZtaB+Tw+Eyap0i1qQMWxd
oBmzufbgrx1SAagBSGSTQglCXTRzHo4ufGkWG22yeecIFIL8/eKM4C2PzAWvn6kfpEDmXyH1J2lF
vw+NPWpleEwLYIv7HXmkpw/F6eOe8M29ZA+GlltxlrNmfw8bnguCBbdc4RzHq7B7Xf3E+Sg5Ru59
2jmiepFEHzZRVRevVSuS/+V/PVRfXF92ks97F/ijltUkzMjQ1wefslk3tG9rzP29OmGj37YSmyFC
9/iyIpMwJvC/wWXUbMkM3C8JavxJbcMLAVTWby+8ICzXUwK7xYNCt75lqy5SuRwvf7bMdyQ2p6ZY
buUzVS5NOw04BuX3STEvhSkFAD9MWvfbYth+KrCZob2dmg/armRFpUs5iq56Lome6FUMTge/pdID
UbvVhnzgUPM/VTvnHGj9J9/36lWvuH9xveV/w0VZoJTSSyBUESnaDehGd3OlokKqfA166i61kksp
Ma0v6Awb3P0GP7i0jPsGHA3b4btZ87f/PJ91gpc6gMuVEO3JSKXWQ8ztjwj8HgbibH+nlRwc3zju
AU2Qx7fzD01cDvHvuN8O39UZK8ZKUbDmOJ0q47fasgj7uPpsT116FxBlZxQqy6fcwkuAyMdAOTdp
8Z0k3qQqZIK2OVdk/SwPMXwZroHYxZFsB45K/nLBEhNwhdRrDF1Y0actiDqrwmrSLbergl1Rwj1Q
HpDqdBR7PRImVoW+A9lijgl+bFDImkrim327WD7Zc5Np659TtsMX4DQThdSPDIEe5lUKu+8Ll33O
BIr+jK4c389GJl5y2onimssmxXhnYW8t6voqRTbSccyTLQyFqRA1XUvkefE/q4TAscuXHZ90/8SH
KWfM39tZWOxI0cmX8UoqHhMUyz8sac25iF6VTYd+CDZo4MyFNhlQEK0lrTuG2IN04kVkDqZH2PT1
DenoZ4VBw11qkol2289ncGEdwWYKXYdBl1VOEpZBN5xqJRWx6EEjraB4UnRwVnro9KD13SRbdYwT
1xBW8Awflw7tdyZ06dEzx0d8Kj/c8AVPnc0mPFyPTOAWDyArDYp9M3pkl3xtQO12MQcN0D97l+tf
CIdG7CHze8daJz62uDKzUopM8Yb7fSNveX26I9xpaXsOrYIW3E2M1Fv6JlfT2Tm13IW3FI+Vk3IB
RxxAb8y4R4otpVr6MdooOhgzax99u1sh9J8ec82/QzEdKqaoRu2y+OPzg9UR2aEY/ZYI/4Wr6VfF
HxCBhoKMbdwVHK/q1dRZSutzbfPAeBOL62uUWAtMnmLzVeJhxpn4mjggbbvsJBeiyos0NGOJ1KUv
8yor0erhyJyU0x/IIlY6hhzJGM/64xjVO2hOBkFU2/Vu7atQZQo+9fKpX9GRU0PvYN5BnQnJT1OX
blXcC4x89FCpldY5ce5kIz1LryCaFGzzwK6/lvz/zg5c5AND+NqM3rHSAUK+yR05cC4bH51+yQIb
Cy8UBqCXRdnla+GTsswE+Ykm+2tHE2LgLugV7jf4NnHY/iNrSCYK41aqc/IFvpkjTh0cSFC4vyTr
fk2Uo6m36WJCq9RdWaGzNW3eCY+HZTZFrKqHnXu6F5QvKNEDLNl5WxsYnLD6hvRfDZ4PdHEelwmE
6uJBzPRD+phOuK3D1HGfCR46JRzKZpxOK4HeQiaeFkzSFAPv1v0IdskXnF7wLMuNvKDg03wa1OZU
lIxeXY2aKQownjRj+byRtc+BlzooGlI18YM8B3UfTz3/z9V0aUVTjzxTxxLnVBDBfUAnENHf69f3
+MecYqZ2Lx8mh9AWcrg9sXF+Y72hNCxMUzdqkPSg+bxRNHAhjB8ta0LpzbH47OZPbXOHbCduoLxp
Lw+vWdJYNAoKVnjwRKRyx0oi77zJy1yM3lxqLTphce4uaJbL2X0QAYLzmN5ndwBJuXUQ8W4E7Ctm
We5+CfXxn7P9ccs2gynjzARMJ47G+S1yQplBFw04O69kU+Gslzzcm1VMdT1wHxgYR6hFnFUcm0/T
lbsrOqvKcFmGiHNNq6HN8orb6x9jE/B3URkWCssFr1+SPqhH9TYCI1sbChdV1Rb/SbZ9H3I7GM8Q
Uqz0JaOxtTqa+++uFVAUwU0/XFVAR8wRKF/eEcXHUHLcl/FUt4/1LfHlR5xoxff3L13gpclp6Za4
uUXFvwkl2WXOKQvJFJaHEGojOn5U3UZhBrPfpyU+IxFyiFWcoja6VZdNz2ogQmwPboDBWtjgis5i
7clr4ByxnpiQrPKEIO2EYPf6Tef23gJOhc0trpvYcHJX/cQw14Y5YbZOOv5b7RJ8OsMw0emSFdFS
Db3AKUXoJcmNq4q9Jvu6LD9IH6QdCCfJZboNWjQwMNBdO03X4SggpAxHfeCHbUqqz4Vs9pwebdBN
ej3yGt8d++QtNKUi6bmhQV36CjImJ/5/7I7zxd6u5hxxk5cdHS2+EpBwSAY18kJy9MSnkJBUGkaA
sZb20ZUWyaUkvxYcHCBW1hgWvFU6dBLoVlzIMT0woJRAMCm6Mx8s9yY/bGngagtdXtibVZrtzGJ0
007Mec5s+17s/CVpZ0sphp8NsjHFpzqaxfr/okzHvAb1av5xNHowYll2gn2AyPIiaMTZSRYmVoHh
rIHNhOl2tGOKj3ZlWsDarnu7UGrVGdwA30ndOrrmTiIvYKsncvKJkRbE/Bd+LBFzaT5tUYKsn0JX
uS/Vwvkjt4CNXsRfYnG0olbLEQmqVIsH/gUbkNXujURPipEnp1ywsDfcYUq1ROj9RB2KfbjVHH3q
lpLp5MB6Gu2EIX5jmiErjIpzLaDPQRxOw02IhTm3K8CdrmhR4bdPFWwS3GV43NZKuuP55A1575Ed
sRyTxY+4/9ak3nA4xf6JA6//fe33xndF8+DB8vhAVAUjnTgBZjEkf3qo/a9i8pqWOYAfBeLy/3mE
2I7OGhAY9lY8XyovW2eHVUGVF3a4+26akz4q4E07kefHo5o8RCUBOT06/TRVawFK9DVPB6zvS9K3
J2bSWUa4EkZvmcGVtUsTt8ONHb5N8xJwxcIMQF39F/h3hydhL4+Bu/ZhBim0vMK07v1EStg79cWT
kIPml40O1b4/edR0lvVJ0wmloMBwKk+qhNkNc0D5bh6eoMpHCNF2P2R9tuJSHUNdjOYk/31W+vDI
3UPpvXcuLiEspChByGb77dsUw2u6xkphSHIzTpjxGE3cK4EzcGt+gzbbPlUEHhkh6n0S1eY1nsJZ
bGHDJVjGvB3PD7l4WRqOQfH8PtDLT383AZp1/VS4KAlgQbiy7bJ2p6oppgQwePji1acXpDt/YD6L
GXr5TvV+36++oxVzhY4wF/69JsNdQeU8DQcrXW9u65+8I2YBQNqIyb2Zh8PcwkCRbuj3KMXnYqxS
6tS4PI9SQQrfnGfeTU28FDHG3NYMw4iPhBzTVrkNxRyMy9B3Q8iY9ku1gOZC9aMuIf4o6Ww+ahtE
lwNpzeFKidNJJV1E3Tr6oI+BjwnVNviGHwMrReC9DZNy0vwASbjGDMzUsxInAWy385yh9F3R+C5v
L9m5/a+Xiz76jQdD+9OQlg8Z9ss3M1GPaLmkujdJSqsfMCRPU+KHi90oHpFepENRjKfWDR4ix1vt
wz/kOv0mM6ctzKjfXLmq6B5TFjxkpt8XvTUQ+9LemophwTN3GjgQiyM6CBsHUxrxOrDmoiI2MBVr
2tqs30d6+GVkxcFinLhQMMIaVVTtwtckozr3NwSOI8tA0pKnJJlUnTgKTLCYPSi68pUPg+6qN6CT
8D2vWce+LmiT2kxH7C6TZ5HAZ+y7+yoNWSXYOl+fSeG84wxUFxLoBZUu5DMbuGMxfaK6bLYA7zwO
5HZXKbQit+5PoxUfOot2bK/O7C4laG4Iv7HjGCBTUNRcZMtSN/GV106RM0cJbsaZU+o8+UNmbbhr
+ATo76lEm3Pib6opw9p1D182nn5YwJoz9RbbJseNfAm4LNbudOYuZlXCXw/lG2RJHOiNz0w9nR2j
622jluPGTApmGjpTitLPcCqVFapc1NuTB9OFO7haFZCHQiBcNgJSTobASbpb/Abflq/M8Z2GwWn9
DwNR0+5yrij2GDumyi1wKCgDPXV9x+FmeKsyEwH94F54/4ZbUqhr6eQzK84sIqj8cNeNowajYkKI
yCsMpAZGP+JRG8B+ETi6MttzYSUOclUwVLyK6rQmOsBRg8BFr1MVrVcVy+tHtRsxVXQv65x214xM
yeHWCkCB6wPt22wEJWlXZ4ibRE37YMF0i+6sNg8VQt4AgJGxJzb9qY47GMhk/x2ZyWdFRryfIq8p
nCFRqZmTbTqX5i95h1wzqpKpa34JPMe1mI1D0FlHxAxlwZohYVKqrKo47qAxdhCoT6ESpElvEjra
1TRlAQKoHf23J9uUKdLnkdCQQKBf5RnzCV7Xu7+DTmj9c/6045INtlQfJ57OMpj9gFOuS8bxtzY0
4KY40VGm7gBBhBv2HTVUWgXsIBBbLfwBImqtGnTenVicsRA4M0WCHuko4EYZOCbqlhuOQ35PrYIq
CIiMwdmcJseFKzI2+KMazUOYkk27yXAbjvjhBYXTOuYW7M2zSp/wpDbHwOSXtIeyEh3Cnidmed1M
LDUYCShqWr6/0MJp4YZYKZog+5ywEWrzQtotwh+R08h+q7r0Zm+EL4gDhxugLcVjAGfk7uIS4OXV
0vUzp7kDgrQSERxi2Qzq92txRpErkwFim7lWQC8t8gJL4Tqse+jmAIlcuMu6rapVgnqVQoJt9xaz
p/RVchuQhy5ZNirJNRw8+lrLXCLfUi4ZfQ/ns8vyqDClO6ejJ7/jRIwDrzQLFHEI7jkzGmNDIL3U
LRmswSrt0hsBHCT2jDKzhYWoUGuPHgKFwSzyTCQJfNYmWW6nnU3lJPlnUWPuAbZHlSOUCicd/EUK
StqvB6tQJupfDnN4nbLQQRZqGArnnxDr33b5YNbR5xLkhQ3dAZkz4KiymBYyTwrtO8nink2Rm60q
pC1yuQODIe2NKed6lopg5TvMOQXd9R7EfcgSVoICw9IYI82VcIWWSyR6l62qmE/6wj8X0UZNbNBx
skkDtc+bcHQItlPbDOAVq73FbgAP4NMZt6MdFAwlgFwZ5xHAKLvsw0sQrjLLjM9JPrnfQFNN25yi
oRoItUYHaWN00ZKHtTID9lD8TOp4ubtk6awsYK+xMcp0mwCHtjurKLb8Z6z4ahw1rU0l0T3a1/8m
3GOJgLg2UsyPF5WtTG/u9Ig9cGQTOsP8WiJZcZo7aN97JQay6rDtCFD0f3t4mfPOjCqHldwrjpwa
esMUrwh8HWZv3s1AN849Cy5aW5OZfistJlhVozr6EgXqUbQTjT6fDLt8eviLGIf8Rak7Hq44wZrk
brVf6yXmf0Pz7bZDzcve4YB1Q/dc0q1HduCivQ8njyKuvLyZvYlmARmQ7YzTNBt0ZTlywauHHrSp
uOTBwQvLd9+Z/u+s3aqmaVaRfkmpZXTPb1H3DgRZKU+uVtwKsWjCeRhjVXgz6fDd60fOcuv1L3uQ
xNxCBBe9ZpoS9bdzVxXj0ei0ltz+OSqZjOKsj5tCwMuJZ5KhxkLp8ac89xgEeDEX3AD7K7ctzSSe
GpjyrOumBi1nhtZ1IS8t1vvhF66BXfDXxC3UZ054wlEq9flOsuXsRf7faO7ZzvBlc5gfnUFQ1zCE
0khDWnwruDqyQvvdclF9wUdUDM4tMjiQmp3nGjWkDts1sY7LH2+q4Qgfxr+fdt6DcQ4HALnquxTw
Z2dIOeby9SKfh4ZoxxMN/jSv8AwYfqpJLSZQFxA0/lKDx5/dKDPoNFc+NQFlFLKzc61JddI1YBSy
YdnsaiAqo8l6Jr/ZA3DF9SrctUMI/wftIv0fLN+15RnKu5awLL6CWv4Voi2cWQjocMLtb3cwi9fs
FPgZysPbrElIdMTTuRcxFsr8k3SWIsdHkyV1mz35GW0ouvIY4EYZChYTDLIxnrVUYyt5P7nyEyup
c8kBEv52b7eQDUsJrn9ak0knwgMU2bVH04MFs1h/SAnMzmaqBLj1TQFXOk68h/YBfhuv4iPSmu0Z
EWTTmLD3p98UTpHnOsyACsEQGcTm9nWssJxnBUzk+8VM4A21bU1NToJgP3CbaAYtlwm30ZQ+qKX7
yY5CodpclEbeC3OiTWModv7lOsTqEuYTov/dZKTEooOfVjRyWIEMrD+1Dnm3RFmEZeb2bjJcbkOT
lC71PL/W8FzZQJMdh4EN5gwCcCu+RwpX4Rs00dLC1Snqv8D3MB4Ll30v6vIOIodN+VPLJ1JK7mjC
zV3IawjCONi8T1vhJMe7F3tz+DpYnD+KtqML9wQBGBv0J1VPSCvTdMlXraVJHdJF5WeClrfPY5eq
t34k9Q6THcI2o4COgs1O09cCnxFWEM1xhbMOPWX5NOr640Rl0ckdDLANUwL+BaWcSroKeNc86c0i
kdriz3Bpn8mPb6x5BzunWtf+HPNP8uIUmaDFSKtj83R3HGJPWrGCHF4/976+zk+jvXvpq+Snrpz+
KCICHqKeAUD4T2QMxcWxAljeydUwO0m5x/+9NZrkEQbUT/QUUzr5GvpmINYqXLjbr/3Zr/sQiKQ6
iXwu0z56+lbRmQiZH/dn7OHeFjFny8MyOaPBzgWxnIf70HNs3445Sdf7Us3vJpUMYz5W/yVPRsv3
QiGjr0vPJTAWvrwUcZH8lAclZP9PrpvjJPjPjnaLPd2gucTZ8eiLZalLJ3wVPYs9F0iT4FSdcp7t
tOPJ1ZmUHWALF2tpf23ZPVbsb1l0Xh/z7zrZSv9Lk74t6cyhK5Ro9BvQiDYMHiMxzQJYeGHNZ6ys
8nv7DfgrfWJmZ03oa8pO4i16jSQn1r2h6GXOkEyw/bVtZh2xUeMFKM9MmSfdjjhvdMLCB172q6Pg
CfatM7OMwvWBw1YpPfXpA5Fs0vPaCeBNzP33ysKdYi5kATKAC7t9S9GEEQgK9XRBN2H2YPrMoVXq
uClnfVHSpLGnQzW0PzZukl3koS26p8U2q6vdw9IOFJzH5vm6z71xrx6trqM5u9jGy8hakA0CLS40
MX16Dm/Bwih6lnFMaqywbAaPSA4IgJHwlFze/Rbv667ajmCcyUctluS0I0SD4C8BxBzfjAl+8TYi
rh6Mt8En9CCrWqCXBDbQJBH5W0uhufnrAB0UFRutFCwRa/oqnGrTQL5NnsCkBcTseiYjAG8X+C9B
W5kyK215W90eIZmk7Ge4urK5JKjrRknFgZXUi+3nRBmCZtwbYud5vckj2yh5K1GsF9resLUzkN1u
VWVfKrX1LCSEFyVhuY34wsmTfE+CLu3FdL87PU+TIKWWqC1azFTJwMumVnwT9kYdlYV+//0bK9jI
1THgiVMPTKadF6533ZsVcqT+4MOVFWtEjoC3vrzZJf7/AUYwGa27i59w4mOJq035fIFNbASPYNGW
83Cju+jN22gLqZLBdQf4zwJef3edEZOUNKza6KjNC5G94mQQl6QsdV89X7RvV6TvZKOiX5rj9ZxE
gRv6E63hN0M89UaP+zvBLk3XTKtuT8qB8AMZEElc2H5W9zfpCsTjjlkNmJOM61Bym/HWHS/4pTMH
N1dQmW83dZq/hckDvAQXBPLf+datfe/zVhmCTqKijbiwDvayPCorHHkSS7KfiocbsK5dZ80yPTJ2
ij47yJzC66kiZpxEbUhrZRlb50+BbUEff6KZGZtp/ky+xelSj0uAJDX+rfnguYwObkxz7ej6pDlY
RPKY8IIUUnCX8M3mtEVWW3Cqa5oWTjUiWTYlcMNtiZTt3s7jQlvLDTMXZYWZCTNj+iHngDS5mDEa
ch/5XlDQ01+h3LRtKy2f8K271A4r47KRasKIG3QDLDALdU9lHvVBZ1yiu0IIEwuNWAIwLzu+Y2Eg
arpoOZfQiDpJ+PytCi6ogstHJQIhoTBFJNYKAZDtQnoa03nRX3/OwoKfJymYgRRykXmx5vTGOgdW
6lC6l9XHQCgQcL+r8/MEZQJ6vEn+biRVgS7IVCRL8d0lVyXgUcke10/+ENSRY1e5v44vjCwy1OIA
XaxOI/PAFY2G5vIDpU18RkbGrzM5IzqWtOcepetDsglqe3SVWHJgTreZUswg2wmoXzkqtev8IQvO
LtpMxEzE3qDMrCFxTKFZWxajvuamiAwiHnBFT2uRwOxz116QbScPR+k6CyXG07Fxb3Lcjf0h3C/m
VFGZJQ0eTQ4n2O3F05hdvCTRHjh7WNdZW6+03ajbTte9Jzj9zQvzQmWvJj9XRu69wmgEXlOm5KO7
YXduryxIWNV/sH/s8I7UIV/whcBWUHV6/2CAEiDIM2qtWhY4DwU76ZXLLQboRwLQqXWn3pqoWtz6
HBOb69NVOBfBjSGSfZCMej/7524gjk635pZMnrASqW3H7ixKMnSaf4KRlHuprKjNli3HXrScFaKN
sDYkG+37a4vukp4/0emkXdlP+eCl5vAXtec1Pxp7G77qyksTtpZ8ZNyCO4iO/mweHep3HfKmJ+sP
tuND/0b4NY6CD3CA9RrrYiMvuzr3TPBLpyNVbrbW0oZDtGDNQvoNTiEbLP0Y5+WbpM9Zq5NmqpfY
WMHoRf3+E2Eo0eLFjYe2uLPfjd/tmvikMb1dZzzi1yoq2s4J6Hfk/U0712CZ5CeTvCjBPyCsfdNp
wXcEDiiud1z5exKaWR8EjQ31RfWekPsA9+o0dlwwgsIvznGBg1MR/nk9ZvDb6jjfQ33UBDByHzYl
Cyhq1DSMVuh7YWC7dDfPh5nr2x/KuStAandQgnwB1CCI7yFs/LlnSmH26zYtC/U46uSUs7JkFb6B
gnMLdMPPjkk7bqVzWztdHWDXgdKA7tlwK49HOWU3RWpPeuoS9wfkrcJp2ygbAoqcf0X55laa8pXh
Fm2glVZH4wnRKjaiu/yHrXuyzQXodqy4f+i2iH2zMgOPtJQrqbHhE8kUudjBdkWB2qJmja126opF
gRslcfboAWo4f9UF51aFEPyMSAE6ApSAWTAOTIoTaIdPoNlKYumK7Jh1goyf68s4vZPLJCrz60eq
PH29Ub7XtFB1AnBOFNtmDaMg1j6Re51aZMpoBOJN6J2DP5z6W4OsEDTJX1BAG1EdNVlnglEDTb3b
wut+H++hIVsiaHBE5xTinFUG28PT2J40LSqp9x42gv2jup7yK2yKj65zrKLy7aLCKgYrhUuAnW/D
9Hvt75ZfOJ9Z1xovYrsmOZHWutB9ziIMCfmaGFnRT/8lfDuCNJ2OnvJG9BX3pvwHyHcWwOs3yZEl
kt4Jc/VujEFij3+ZTtrQb8ciGIy9XYmP/qq5ODKB/ubjR/Hb7R/ZMe9IXauG25xXEfL4sGJPsWkG
3kwzqAZr0lO/MEULTLHVyfNpAEGI2JP1l290EoMoVqxqoH/9PH7TCwySYE259ceaB3fpuJ1xASAE
If9dsBRGUTNMdeAO9sq3A7krohOQ4bnKUBusjQwIqPiY5yWJNJulAkePjC7hjLOiGOnhhf784FF9
GT4wQJTbiO6kKihYxGgaJdNdShcnOVAUszBJ2qwZ+3NJkbNCW6tF/U8IxmdnlZJYJDiuoqP49QT4
Ha8kTWdk27CKh/8PC1losiM//6zHT+As8N/wKrgrJxcc6oWSw+Zcc8DC85FzDttNtnKxFglzLmro
PTPZwZTZYKP15uUw+mXnJn/LdbcE2zwtE8zrGRpk2dXU1RnAE7cQ9V7NkCoPkW64qT0RTZYO0QA8
JgjcLTOXhAzSGfi7NO0CD+8uxPWwmh6FjBW/ZpBFdERWbdL0EikBLmQtkunVFn9KFM3DF2CpF45O
u/wEjLyBlBlrolFi3Wk2MD30ALtF0xxhvnkReKNfnvwidkdv20Zw2G/j6whpLFkW9snhELdi1s0K
8oTARJnLuAfI3uIA2oSWr1DO5fYQ8Vtr1rp35XJ4WasIIntxPgtDnV5ScieRPymeY9Aqo5ynzOaL
MMuu6VHYVQzMJC6ASlckcvjhi8i9gkiXEDvzsg/IP2Wy5TysUL0q1aqH3JngUMBJ+p7mPMOM1fQ5
3Qtb5pWJxw/GLyV+gdFuQx5ih83/XmQ67Dm2OWbqm/kjDWiUTXm0kGqimaManr1rlf57VECd4KAx
gwb+gadFAdn6A6+NY2BaG10fayu5c6nWC3yynXfUCiwXWSyv3EGhx2qMQsbAwRfk9tbtQ0wL0L89
eJQfZUnW4gZuGlYuNJE637fw+58ORM0l5H90jkVbJFzN2+xyJDXd7qRgrbq3OCOQLLiPZ50zTogQ
qDFm5s3xCWBEUNFnQ6XcXLLgqmVoR0xG6p8u/CnZs58OO7WAvs2ldvvU1jmCWMPLWK8rRAZsTZux
FJGwGJswXKg6TkwNiV8I2CJNlCoddNI+Jg1dYBxuuVW+9hzrYopZZb/DYNVLgZF9mHSKuGfRqxX6
wMTB1WJiku4d35iTgwEDjQ7/asl5iw7IMV9Wgdn7D2nNJpzw6+n8gcteZagQ/U2qKr3rnw3V0wm6
3zRqoRCOqWlIhzDHkMqgvp+I5Qi23WPl1LYHy65b3Wg0BqrEvyh3zwgQu8gTxJl/oa8QQq0jQkiw
DBaCzipM64piV0ZWbCT4AAYTm/y9DwoNRFw2K0hi1o5Xb8qoD1y4XKByIUevmiqOJ451T3gSENz2
jyo8ISkzVYGv01MslyuaDWltBEjS09O5ehS+wVviG8Qlj0Ffgn3UF5d9ZprbjF4/NvRXmV6IhNHM
pVLTfQLLvCiAYnW5w1C7+QalatUoZVoKrPOl/Orc4skkFrRN/IfHAcrfzx65qlb+a5yBfyWR0Eds
utQesUwIO6uTN8oC3OR1OxQSs3qpNWYCdVOdyU0oidRFFdhooWWAys0TpCHSGrC2AgMA5jejgwZy
PrQbJ6bJXjlJM+c6JFl7a48JDPJhhUMZvfHJrb/6zrQp0crTpljEoTpVCmqgpK1nQ9j1z1KPFF0b
F5mcsHE5t5iuynJQ5f6wydDjZSeB1Oxzmw0TLgVQW8VHoESLtbzV1RFo1g2sY8zjo5QH55H56V9M
8kNeVMwQCPZZE1b+JzRyns9pscOEUXaA7DDxKml3UmFmJ3+MeHNu+IUDlV5M9/GONVtZoPzNzhte
vykpJvhYhNp4JRoEVOWF1Rmt8gVqceBCKFyiBqTCjgMGH4OojcGNOhxsbmsUjOUznJq0ljpjvaGe
ORV35JtZSbA3vYw7qB3VrNxydok/Td4oKN9/lPAchxL9/4bK67eCF4DdE6QRRODPya0lbXHV9/j0
fNkiI3HvJCOtkVK9ryqN8Yol+QvJn+/buPS+MAI3AI2Ol3ga/xZ4IGQeyjCVucuw79ri4SLTIDc4
u99IEy1QbCl/0InOHNS4BBl6HwSVwJXmHbvKxdpGCUI5iCWyYub2xRRKAdWkVO0O5v3+8lLKUIor
Y6nL5VRMQLNjra0cmgjdIWxaATlGVTOJaeP96oAfS9Dh76s0iFwRcxzxslYbiGnja51WOvrTXSyK
iySJAEkN3VBoCdBKGZWmkWCGdGsXbonF2rMZ0N5xPYmhdS+fRQwtXukf8EolDcgLDRR17cjjjB46
Pu1e4BdCYcO1AE6LXb7YRTMmH0t6Gp+c04ilTnduAydMYCpu49Cr04viE/ETBr39QLwSfueyKZ95
6wZmSUg6zs/0uYM92k3cLXKJU4dEDvTQWJOL8xweKYU9BaTQFqCKsmXv84cfKDsqpksUDvLY8koK
0Ae93fBdaynK6hq1Ia8eek9YuBxO9EOs9KinTs9eWbfr8n7QT9CbuUu8D5t7JuAeyDVTX9/vgzHS
TJ2dlzLJpDM20JgtV46P5lv4FINyN/htT990XvdeRydZPL/10cRXjvkZxO+O92LnQobpKqCWdaM/
z4pVYr7zBeGQqeZhNe2e3Ax0ohtgYFBVl0IlVnbEc8q+UX2Dw0pD0pml3/ZEm2TzSgq02CRt9Bbh
8EMTmETwz9hk/WHka2vF2cFPMWHXtuSqRLa40xQJecgYW8gKR0g0JtCcJlp3XXr3f7SETpf60sXO
0A3EA/4epnH73A6m8MQbJn8iIiXUeKAl8RKM59RW46vAohKLAuZVA9iqjQ5sW169S/io5DMd6IT2
+pmZlVg3m75wGMQ5tc/zKxGyEt/xqsrCxiBZidwyDsmba8zzY1ehzF58YJmqQt4OPYQ9p6BXA5q/
AhAhvBPlZnVk10VzCNtXhuiNnIZmXQ8ym2kI4AxkQc1tOiU639U/6QtIUQspYn7KUIPoYl6ksvM4
JqG/pEtj99fPYDd19yKSrSm01nY8I8MyNW+6/oJhUoD4P6qyzbkFQF9fDBZ9VaSqETa76mMIkmFn
Y2JPNbyulsoMrV78xsk0c787TLXS09rBim+q7vDHvrrVBSV/5XhksGONoTjnpb8VGs7w9RRaBJCg
+unipCkNdNY+ri0QRJqi9eFIa78sazzsvOvQaaikmHiO9P/uU7Q8lGpEzAZKli7BNnNrofXmGuol
z/O7MglTKSC3en74qZnkcwhkKYvuDv5Z7dAJTPxUriny9m6nmYpKKJsM/LP/58DcMfn/4oux4eSu
XVms2pmCxplsv5O9jX0Dp1kx+WMwzeNOk4Thwo89+Zy4lzA+mJv6b9ohn8cyGdQJRDapAkZuBC+g
g9i2EVkZYRemMAswL7M1FcZDBd9k1otX++VlWd3cR69N+9jCC4LOgMCXxuoNImsWFLAt03J7DDyl
rcfmFXqyttXJs6Qgh18Ox+AzHTqWedU557VTL2xTcV5LCx+oWphL0jl6/tWvlrgVzngcSHU6+LmE
JTusAwFWqM2HspswEbllE2hhqWLZ+q9fJMNx/5c4vfJO4zx/+d242Of+9VX7lHpvF/edO8VLuJeo
NbJLnjaSKk6VD24lLSJRifB6tA8kusi/AXpCmYbHoJF43YuC8Wxb+Hxx2NNHXchKOcx0Pj6bo6cx
bjGDyZh6qH5UlQtSHRqMHxaAVNBS7o5CYkzi+K0kcM9Ud/tQ+RmrV9ZW8UjpJgnT6Dw/WTIsKNnl
NZKyrNzIFaSOGgwdf99/nMAwDBsjxJq1xFkf4V7lmFU+9BxA6hRv4FsrYT40c6/oOjCAwvfqzJzA
u1vaq+wnLu6si6sUgJtSxn4YkzUd4Ey2a7pFirn3rM4TBSrD3zGBUVP5eb5Lme0Zjt6VDY+3fba4
dlBFrKOm1d4gBw4hgzVvrtxl1+br9dY8SzLJ2Uv8e8VTLZbzJiLOvYopSGjcKdAx/OdEa4CAl9GB
ki32ZNmb4sF04WSS7KJk5xJHoCCAdBhLfIPeMw0xPl3DVvyq5VYEPnHzr2Q0Ixv1wqQ7eRqzigHk
JaHbDz24DAuDEMYtQA0S/50l8Zfv9EJrTh5T+V+VME1yqPyD1zDR3dCbFWxNoVvgqEI6urrBEGI/
0TZQ7BAaxLGf5Rvk6lAW1HbEUiwu4TDD3ysd7SPWcCvNDaqJaNZELmHuJuEpkIVvWkVr+FtzBZmy
dGJO3T8qm6CvxFfIEZKZnvxZwG8nwnBwzXpQP+ddweMh2/NP1z/IvDqhVevsk7cDd+MNI9OA/yi3
/e+GKz/agDD3cEFvAeT85bbgiEmeIQyVvruJYL9G2G0YzKhGXUOqKqWv9djOnytecUmHtMDKssvY
DbPg0gsPMvi/M3W4Yn/V/p1QIik3MhcsMU6IyiCL2J8Dr44mo4KW318OJxlPDctIZgqiexSI/DTH
t9DYxdU3ZsFkfMAmJVlBOQ57A6jTocQq9SQPYU1F+P8/cEEIwDdA2bETql2RR1+yVMQpmx/2v81M
WflbG3XAAm6eLUGfwwa9HBZOAhyxHMxipAXOChSLCeaiZ8S1Ni0RQ2bxH/4ZktEbu3Gq8kZ4COo/
B+DjonCEUwQAoB7B2i8gFu3shhr2Dm0SbhTZK2REr5VH2BA+1yb7ohYXJlMvKj2OAk9IFGQ+dS0+
jMdxWhuaw+LgSLVUKQ6Vx8xA15uIc+G6GRwm1Q0VYciMpZmR17IrOo17mPSM2+GIat0eNHf8vw/M
27FqDl5dhWoGrOCvu1sFkl9+cEpMJcF0egSPUtYOwjrOeoeHf+JpkBP14xxsHWergY4vPp5AV58M
IxSlfRJMEQ//qvWtkUORpzzh4MsSdxsk6k1U3lknsCU1nnrgZICcZsLZIxK3mGBTnnF31Tvf860T
lNyzUIlCdH6wCS0ffo1ROWzxNEZ9506tmV1m+7XeJQkHRg9So7W+qN1k+gNRtKZTFyfiwmu9eMPP
g8c4DVibRj3XBMGrM9HPoM1eX3Lt5TYXmjU2Z3LzA0zPDc/XTnjHAUS2A3Oexq5Dw41dBaMqGGsW
4SCiDO0PznEpzhT8fxOzNQLyhjXzmUXv86UMCRqdyHDIoXaSEyX7GuCfAkpWxydNRYxmsi9o3FUN
fUZK/Vr4jNYSb2P0njnT51p6AUfs4xY47M5kmKaZJh3lNZeDN34CS+Z/QVPM2aLaY62jv+X0LVcl
D7Xe+MKL0QDwfoyZGaOUt9uw0Hx05jbFvhji9Gf+J7KOCsJjpBxkJ5hqNmvhBdRUvL1063U9qKL7
8cbOXEtW3UPdXuiDCDBR7WxeKWJixaW4t/1rtqBWms/pGBjJQG4YlFzxn2GpqyLpL+RPk/G4ocEr
Xwjvlf9O0RmEVK/CE+SdTx6dl+oFYxf0QKeWXbTwzLKb1lyTzjg8LcOwLcN9OHG8YkaTjJji5ZHt
zRusQ/kRgeSFG/ZwT8U2mKCMvj3LesfxZ5Ccaghe4JeXftelnYPEtztMO0s+O4xkl7j5MiygwQ5T
TW7PcKDq8MQbniXgvO+YODGBcXiy79eTF8RMqNBdyi9+CWfIu5CxSBP0VNn+VHigNjRYImCPmomS
NzLz1b9VIY2Oo2+tY+ybfayZXShUNsH1koG9kOBrU+vNYtsr300s0AOw4atOfP9dQwnBQuxsPK+n
hK3ZSXL3F7HqpsAP1s6UlH5sx4aQuxtFTEI1+zujKHNZXA39ae/QH0hkEwxCUOCfPydiOFkYak/2
I1JWRwrqaj4+marJ8lhP4xAZ5SWdBc44f7r6CwRWCimK/xs/ErTPBhYhDY+c8Lw9O2ttHo7aJVIo
tN27sE5JgWygWK+Eejez6w2k/VU8fy9vlr85P3lGKYaenuXUSZi5E18IsfywmZS1kak03m28+mOD
BPer13KTU62816edAP08TkItkT8aWCmhmG+U8GzuHIzUL73XVLmodCF3O9uBy/A3Owqxrziqx7Hz
/Omefej7ehgyWqV1wfU/uWm/1AuOyAQc7+1AOfaCuSPMILQ+Jth/bdhBcsjJWOc++09RHwJpD2oM
ti92Nn2/dqBxVTIFgeEfgjZhxTnefyUQ/HzELWHwYmOwFkVts6Z+4p/skk5asep9spDnE9Qwa7wj
fCzSQqso2d8ENgO6IzI7kNd0XCi0dngpjIwen0lc6/82NDcKDGyUj5fSvXgYbbZGK23gTjcQvDmL
vugirI8EcYAu7Aih224ry/9iMfbLkFaRHAF8sdOZ3RU4ooZQBeRtTuHMxZ9qOvGdvSXAGjlP+TQx
z6OtMPp+aM+ryWuBAs+hvktcQbJ5LIFcUPFMuLrfACnVBc5QPW+nrSd7NlfFSTrXkUWi8NeJSlin
5ZgkUxm6Y8PzaUgLgAwhmHZdSdB5wXqpmVyLMmbH8v+3Z37XZX2Mb52lhLDTEEcOktdivJk3cU9D
v+Zo+9DO+zpfbLUf1Hl+G4rJJKtF7ImLJfG9Ht060uRuhmG4NZHEtPp1NmjKOBuERYTlGE0haVTf
Ohixlg0HcSEt/4D0p2cKNDfg6VS2QsYLKZuokiar2l1Tjuq3fKli8PJviMXrj5MVWwX5U0hxcj71
w1FdTi1bLNIlpVwd1JmFVHuXz9awlpXq30ksWGaK4xhUeUEg5MFNpvkK5cdbTftYmV7bSRf7Vcys
AjSFdLUkjEFYMCk9GF7/qeh/ov8/PUJJnwD39NLuAtB8gspGwCdqW9gPIZRJMzdQhPlcxTW6Efyl
TLwvD8+nOHCKle6na/Mawmxc/o+FjwkCvNdsqIsVnTnvoSC043TL9aAKGRxPWZcVODRwLYPDwtqv
SGun1xlX/r67Kdeopx9rRrHtpKB3L4L/xewnHIHWlPyAVgEmYjdypcnTRDDtghOFOZdCc+3cfJe1
IMFda4gOfOyMdMIK8PwnMxCf3tz9ePtsU/aCY9SyfZ51NvF04nOFosYgoX0eDwd6w3etErlHpxje
svhGbjr6Df3oSu2E4r4Vpfpn9N2/xF7QAJysWauLt45EPR2MP8HvnV6mJKAD5Xsy22wwvxjQCe2Q
LA+tyuZO81DXQo6f5Hw4mD4E9L4rt3vBRLf/T3MEUbCUQZu+PDMObjAuQwIwX8OyyFgjcGfGY///
b0XzDJ93tKOiFIZ4oDmcxsbF83rWJ8AOrcypF4K4WM/m0eKhWVDc+oGCdwNiLY1/GQI8+nfWlXWY
8dgnf7OKo8Q/dGNul3vTjOyOPGA77BaidwkB9GE0WH+Ywv0kgGgRUavvSxAHGRsq8l++kK7XX1n2
wID301uzYv7E74L8OiJYPc0UWxzOwq9TOOlAHIr2t0vhyTuqr7QLFAe8YkKa1W7lNS6zFOHUtz7o
gY2x5dfiIwZnAbDE8qmJxx0dBwTGSjMJnNTWeCbnIWTTdduzpKQS2ttjoaZe6XFNo4jzN34rBNAT
HFPrqBuf9KSwX3TeDGbZMaE9h25ZcLLXY6V0znWCztGumYrXpJgLZnWPI2L68sV/alYKzmnjzAq2
4EuhxrWOvQzdqv+mMLzbNYJmex4I/6O5tKa3QmTANE97ujBPRhlGj9w0NUv1z8NgUitm8MMZGePt
QRko9ve5u9abmm4T7D+Usso3etRcSQgu4K0MYtDxviFIFZCHfLxX7ot2iVaxHnwX2NADqHrDrMHH
C3m9WzMSqtGTt7BNd1mNh0uvhUXjRv2pmx/wjGAiomZdxCWEHkTnAVdf5YNmO3YTvn2HYOlcz7Rm
leMoKCVL9wwkqeLA1aPTveMwdSNU+8EDC3ADMKxygMLLjwyekAjVF1mHwatcb+auH4LqdlE7J35H
SWz/Y10cRxwoaLNTEqqyhyhyhBtR434uoNfW8nl1jU7wyNvFtKS/eIp7uysae9WZQFrvtETB2Tj3
Bg8liXhcACbcyudY4ALfPfjiZO7OCvokcdF+WIVSk2zrcF9DkqHQ984GMJLxo9O09UfnyY6tlfeZ
QX9bZde/107B+nhoyx4Aladdd7FSXCYPVtuo7MJI3YJAGHGD0nCn+T5xg+VjrWWXoLWpEK94StD8
cHdm+2e3PrE2Iizcin4CBoQ10/yQseSek1RkR2MPx2PiAkh+OKLD0bSg48BYvluOjzzyWf/Y1l68
sbx4tepS06MApobk7TxDTvg7g5PBb0oO8MBm5s+uiPdsLnqYJX4IencFh/+heob/Xz91oMsV79Lc
yRjtQMizZkZx4HeQf0AbJKM6RNDuV1JmDNMCB1LQjTcoNpSKnODGaZJa1LOZTTHAABe1dgpXUYzD
Ob8M+8Klfvw3AdF5BAtVjolXf/8p+LIGXzlIH/4+VZBk/EiZxFloQdAjeU5eSRJq8mt7OQvdgv+8
n5LEd2vl61fpR4vgGTwclg3CgyBaXmNkQRW9E8WIM4fnbHF0/01uLNieMPOI32k/7Ky/s4uN2q/8
aXCv1wCt3g3pOtymlGrQl9mNokJjDcsL12LUfSFd1DtT4gwQ3zN/NhG3QLFCvHdAJKeZOFzmlUt1
0tGzcXb1tH4NwPnAQIJVE4xIXrmU0AEyQ1cMfNL3AQFcCqeS6wb00/RDUyLGMbVfCntwcQmspc+T
0paAs8ZUNYKVf/6IPsu4MQVXbsdgmoBCNIjVX9qD2W8YJbDvIQ7YB+R2+uAGiV2wD0IpZELHJWY+
Hne91Vld/4D3aMm+uhYEWwHKCTlQqTQHfT1DE1HkSwjiALzYPcTnqICN1u4AqDtMwURbGEfbinHB
BgPTpoIRqIAVu2tB9R2YqQdXxux/DScdubkCn+t2UWVwL9ywfhSdh+sQdnX28PFN6xQSZ2xnH3Dw
OMm9P9BpvuwPaZKILXgA7HGNPO7v2LIyo0QhCaDQ09atf+PYpwqSuHmY4NZL7q64oItLwvKbyaEO
cALJ9wJPchtpLdr/NUVvWY6eYWpEJRHSUk+448g7i3HHGzFvbCUGQ6gd5Q1hAH3+HGCN3dUehXoh
a6Fyo2TSAfMLUdvhVRLymSZIDOS1fjXdddYH4c6CwYMSoH0tj4aGZFRnuN2FQYXySFyJsIPW26BZ
MhoP0BDCjVGbRNkldKNu0Fg3A/1bPzto9iT8t2hazMNHCXIHL8rKLDaMuS1bA2FHKBjpl9AtIRan
5nnJ/EGV5VmmYRIr2ZGQF04vG3oMGb0Y15gcT0AUPiQcfH3J2ggofYb9KvSm5TOVrgo1KqZyoyax
qvYCN/JqyV1QTK24uTNv6cPHAuRh4LTI07Gs445MKGC+Bvqna6kPYGChl7tJtIRY2mmIUnWus/V9
OsB2GroFcCSo4ff4HxSquwpw8yYrjoXjGapQOxbB1rfWZ7A7TtUz5PDxqR962Pz6QMAy/0s4RHaV
uIMhDOiuJCkn0ybEu205K1MDIO+lme8Zj87CTWlDFTU9BHnplCBBfPGfc6j3Tcu1uXjarHPBwIj5
bdwDnp49bdpjUokb+8u+xV3SfuLp5/41xr7oEChKIKMrC+PI1d8GNY+/bqOOLc+I4rmAHOPskDYx
Wm/XZfnwbgxrVipe6wx1T4nqQIfiIQ6+CmHrBpRFpSk7KCBCHxvy1haaKH0GnYkkElzTA8+1tjGX
oek088tzjJmjhZW8GjkBs2g+eqaqACUOYvns8/tFn3OOQWq2HD7ijRTU/vUgbySBR94PIcI2mpDF
eByuKv9DS5mYT/XpBThVphb46vQe6EiNgic5pWzXlCbnGd7KAzZD8jtcNxsDFX7wr73jMVPUE7Dm
ig0Bpa8oZFkrteEPkZioi6N0ccNdceVOHYZ1DkzNWcRkKRb/CeQxusiRUxDqq752xjhvP+Em3I2h
ImBIbLyAQM1bJj0kjPDfSpIik5mJSjPUPicq0BOehuuMxKdUxT9SudCraq7JsHBhCforRUUo21em
AmlDqGiZ6Vb9C+pTQ7URkrGgTnkyBdYKJDQ+zTf7sfmxApoOvLDmTrbn6I/WMRs0y5VcZ5QYI4xY
A/Hb/hFEpeuTmYHesxqztD/BOjVYoD6oU6vPYbdhKZVaI7nhf6dEk/xnaXrl4Hw1AU5wdjlouh1h
Hfoy78PJMahKkYOe0QhfvnMj97Cy0+9TlL2gk4JC+hLa5/AAIW1CL/zu93z029ejXfdhSJ2ViEWu
NFlhORImUIhGlsTClrWg+axtHGE2V55B17GnILRgTsQoqIC9x8uh66OyODEk/PW7XwcTCnYZyBEU
fgWa178LH8AhJR4FqEPVasPuIAwkZ11oW+KiOs/WcoPykhtkwBfbJsDsjdoE0sIXS+PYrKpkbO2h
sTqHBbG9Cf8h+zfjUfiJ+l73TDGR4Mpw7diHVhr9mNP8hXKz8Tb8PAcoyXO7B+reW4hgobDUnD8t
VV8KTmJt7SeNxq6WZuoAinDfzPnIxypvb95p5NnkhavYuyQuSmhUBX2TqVyIx08FsDjd6Kf2LRcR
9/r/ZtjGHXkOpaOId0oet66AH2JF36Jg1HUeOGsoumMTN+73ToXv9C3kImYtNEefI6be1RGxtayz
yfD8GugJuG27LJt915r+N3UdDx4LFNfp4URfVIK19O/lAmqb40j/VsXPzwUC0tU4YCD7VhOk9AYO
0S/DHHTSCeGgq3dh7T9js0iZMiXQwUyWzw2QmIoo13LBKe+QLXBn9n2l92tK33gYd7s7oIVmyrRi
1R0lRrOPT6ITgRZiRzn4HVozs+WUH/Qr6DRnVy4+Hl9lLk1b4FMolRia97ngxta7C0s9sXN1xW8V
JVMpHe001m339LpEFqx5/tmezus1LSTyYJfm3M/SRBjwnX9600GawCDgiybyLiaYC+n2OXLuII48
1VC5SwmnM1MveKuvwjux9acRJl3dix1DXvL3hI8L/tXTgOKV70kJvvtguEIlWD3BDXcL8zjz0cAY
WbJc/tku+7Fdvxu3XACa1eydgnuPb2ettwdpcVyyoDYY5FhKG276LKmiFkW25ib5RiVGXgAkEKZJ
9k4lxJ1IdLSuJ9lWqrNIJdK4kJrPJem44tYahjWmOC8cCYWJDTB6KPAHL64iJqd2XVKwEQIaxq1j
Num48vk+cQI46QIYe/HHgK0CPHnpROFutyqxBmfYj9Nq1xVBvRAtp1K+dAQqmF+rPsX0FHu6CE2/
3PAABGu4Iw8RzEB0tYujSadjShCEb6ElrvmqdDjkVXI5k883EiKUUZWM3jqTBHFAJ/PraWdXKknT
9UvHZOz76SYn/KbVl5Ha1u54pVDzEPBzSit7EY9TXhDtxDU2FEYhQicNoGBThqGLdIgBRy8vIeQ7
pwHRNj6EyGCu9XMpn+uEAXf1JmV0RSw9pVDXafajCH7Hx/PWZGnBRcy7WFOu7i2cjQUoXTxkRac8
XH2Of9LLyAfAYOf7CWt1Rinu9NcNPFyfitPTfJA/XNTcF50I0IoHLMhiECHnoV6ZzlRVKajDKv27
UiR49K2vFjjIoASW1zafEAA6HSnHnSsHS9SZ4lcNyA6siDhz0OsCOjyZmi4xriE4WSzyQHlX8GBR
FNJEeh+Qx6Zts5dBP+RxzYx/ppGlB5oNjfc4PsB34XvfdUpZQDZSp0ELilrZA6vtkWOlyV1CNIcG
yJauWMaOrBqV2lr9fbVTjqaTqQRGmO1GDhwEzg5m+Jh8DEwduwGL/sEKbR50liPPlCZgtrjC4XSp
AjPHw1yvuk9nvI3wAz33wsGUJlrQu+ZGp14OsXEPr6CwTa1NgnWAKIbNKH0i0aKlSA1ySNvNLLEk
MxElOZLgE8pfMH3A8mmK+tDM1vBEGottscn4yqB0K1j3swOMMU5XMPVvT/qycHRDZVHXQo8FuQ0H
0rsoECsBV9lKGafFAiIpfZYtXLKSUGUUWEcIdqjZit5DI3slG6/Uv9IQtrYashpOFa8AhR0gP49O
EBkFBxnq1j3blw24WBHX5a7lKVkQ2R44dIEqjuYe890BrQ8AOjl7o7D0XklSJfMglJt3sj8TQDpL
fN3S/XCQaNOXEnDZBDQxar8Ipdqf1Dv9jsIEnzbIHrXfk83q0eDzkQZYuBX2Pml3/ijwOUqY7K1s
SoOkSGJ6xhVJwFxPMjViz1Zj6RS483f3ONZ+FnmA2awnH5Pr7r3guDEbOt7z/7BJMC4fzIaKDxi/
JFACstDo+CzOjXJqy3wwO7MfoT3GqDqyrQ9OBcNkh546zP40TBbV57dIpoDeEjKl4ke08I66rFCP
AXJoluBmsQvpPg2fN4JVSR4XVG9DobgGGVnhV0/WikPE4MMpgXVmYBcip8Tz6Jj2oxfPSU8OoPaG
JehyUpk/SS2tK9VSkLhLXsHSWUoe6GMFec6zGoraZ+3hVQfdrpNu+P0Iusd0++zsDQhoGCIRiAVf
/Og21pe78uMplAHtKao3kc7/mPVdREthEpHAy0VqEe2sibIC0Qv633CRqXfNEU+5K0iCPBam5B06
6ipAMI10tLR4DN7DfTQWFYQgH8IF3PZ7HgSXkpVUJiSimhtCOe/57QiXp1zoc+ZJvEz2Ri57bvfd
LA4Z6R1Aovogi0MzvMj6U8espbJczJ9J6ByOfzG0eF4hM4fIPw1V7yOe3q5tYIBY/NfZ1OCy3mq6
ev2i5YUxRVcLn2GLVlObq8BiDY3eOKxOfplMWE0yEXnq1z6KDDrjvPLYvy1IO+WhJ4/0/YqMZwmf
XIHJTVxBaTbT/hoUEzsblGh1WfYNYoiEfWCOaKaNC6pj4AbKjbvLlFnGyB0OMWmKkG6cqa6eVbOs
TNUSG8eaHqffxgRx6locRtAKsPdHlwqwUbi64zWOSt2+/Ie/aSULzGqEHT04nywnEN8ISb2u1u46
ivafeLeczCnVTlktJVzuwWsCAtshfN1sL+maUzQP1IxdK3VbeXERIcc99iB5/IaZaAmNbDpJ0irU
FouRjeYyD4wZG9+MBzEno9Md1dU5iCiR6qskieJgzCBY3eZ+pceVeVMapUqYguMLVPWsfT6TjbVC
8yvAZnshItAoae1s7DPU6NhqN49vESSHlXfNiJzbuyX6pLmjEMOBqyfJ8f9qffWEmVYy3ObYfH2V
cjkiLlPhCMV3v7Ky4R2YkmNYyEBO8vRCtKr5A2WRIYKgRlvQVdp4BSliYzlLyJyFsr1tEaKpH8Sq
HUdFdIiXC1l6e+hfVeCWZs1C62OiwiZJ2pFwX7JzSt4Pf/Nza3HwlYxDoWhO5luSQVYsKrpkqUtr
lWLcxv9VvG4+z97k6QYFy+HfApMnBlDjUYDHkxk2wUTVbO+Vq3YCaNQZjzVn/7ME5i3EFNUc7Jix
Uqmh91a1PyhMuF9Zj7CUsef6S+RlUi5qgRj8PgEcn+00Xx5cnR06fZ3JhSgJ/lktPMCdd6Pxlgoo
YmDSXcH/ga3+/53B3Nz8WL7pATkoRI8TCe9BuHn09eZJjKuUOA7aEBstj7DVKu9Df4YMiMb93MD3
iIytno5gsk+rcQwVoVSbLK6GUnnciZFGUB1MrSdWKlFuwphVlz/3b0EWF8ziNS/rrZ17JmVKe5fP
yKyPGz3GNpqWVM98jUh4zCaMDjWw8Z6zA1mjlNqkIIoB4UBz8FuvyRv/A/1wzLKeUJCo69HD9BKf
QekpqUSrdMzhGpyZx38NJmLWmNRmY9T2fFa8Dj8fD1hx9YoZ5B4rmsRcoQLsy8RflLQjCDi6vF0X
jdG6SoRjdv7HSh/tG1jv0Yv2AKexVFEuXtbGwPVdO7J9odCfY2afSLz8tcwH5q6NDua7d4U0svOp
QUxnpNSqwDGSFeBHqn+YJIPhuRRAx9EW2YbdNDe+vNi6dYNpxbx8gOREjVDKcrpAGDxyeAixfnHa
NiIDo58nujHYN5CGBzorqurTJSate9n5vzPT0iEZh2Rp9q1snqa96Hm9nmzfztW/JHgMTL0bKScp
RPpnF8Hi8FTBoRbQcgohn/iibDCSpGpmFyvJeBPnBP9t4Y3ZNl0XJGyVTF0iYEkmSo3LJoV/17gC
FsUXOI5B89fuOWGRs1j1ffdbjNxmS3KMU5wyrwvsRsmZzRFE62x3/vq2RgGwWT/zJSn9ntHARBjB
B7/KNFRFJCCl+V1kbWw76GaReNen+CSt6WtJcA3sLzw3SsiP6xIcH8p/UVb0fmqllKJ3ljCyKeF8
BKdNZEg4YGvWcIMrXHzjbwXHhXPK3/wnjdt6VFpwlmmMhqeoCQBlWGSautMzpMr8cSm91DYDeX8d
/61bJ//eG9zDeR4cU4/pV5Psecl1fX3AJjUB3fxtXhpLb6SMMZulLDQgAiXekTJZDCWO1SyEkahT
kj14cw0Jx6kN/RPAwKsq9llyib4jRYXbJVDbWM4mr3djL3RZGv5Bgcw9iExdxGT0bQ6qo0szW+am
+wASwN1ZTgX1Urq3dE6CjEQL4mqCkWcSndjtel1vO1mvMgDC0vURPB1kXmgNo4OK+ICgAYusRv4x
uL/yuUuBVqpt1H4qHbQ7Yc29BJwrD4SOeFmLbEZdULya/c9WLaqDw1wcfh8AmjbQYm+GLgcivbq2
PnvO3QnzGz773Sm/mcM89P1EjfX+aqPeM02HU9nJLzSI4hKli2VNe/83TNYLmBh8qZ2WBn9Hd8os
D46rLf3XAnzXTp+9xJKUZRLqZWBj48Qv9TI+yhwPiOoC1rRA+FCl74tlxGM/V18h9iQnHLP4b9NB
pYr75+5TByKAV4y5ldrsJZMD8hCZe8wmoDQf4VDMVsaIdpLxEY9tWbm4JYJNB7S/N+2viuNEKt2z
bGmSxNDycvypQk0myW2Mr72eIwyq8LNgQ46ndu9pOICFtmL6II6TWwmsA6OflYh79SMqMZQmEYg1
hTs0wrq2W2ouKxOd2iDeHkDqqNmTzx77F8HUFK+rX1DAs70tarlMg0W4c0/g7JBhPhYPkIT/ZgPs
csJcbST4yzxNkeoltW9dc6vmJmpUYMiprDgzaDBVJx/HFC/R8BUff514S/iPEHDoBh+YjmgKVeNz
ZNkarxJdDNlpiX0zDa/XjSChaA2F1DIPkEj5sdxI24iWzO5rut/9oGdn0CZ89K2jTs3Nt9aoz8Bw
uYExxghZQqhS+7/FnZjkwvipxpl1H3s5W6O60zVGI1twYGrdfs5DN1JvgTFHGgCzxu4kdZClrFY9
hqmPySM++JS5teFb9slsCqZzZbp0cNotVMQzteoZLDtwnMO8ylzrXWNnwq6oAvigV7w8PzysOvT2
CRviAJfPZ0nXwEjwjquZXTQs5qEgY5TGz6r0RmrNPHF9lL60XhyOWD1Tjiz5Jdc06Ds4znEIH6bz
ZxRG/QhsDnI7/IOWsbMbEWpdRkzvsoWlg0cWTib8EdGnsOHtyfxurxF87BXmg0mYLuczeX2ihNLu
q9TN2vKdCcVxZhtdYTZ77Y9HeZ7hdt+cb7/UwKZl2qMtGIPfXbWSRJoKpvUHQUmzUW5OnrpmwlE/
xGYQ9rCfOmUx1ye6mzoDcTyrZTBe/d1IMQyLsw6dyG7TgBDn3dgrsta6JbuNzJeOge8rMh9dNy3q
k8hB5wTyCHG5w1kcAPYQnX+9kV/NZN2Boz9j83SUQAjrVGvo3PiP4xhV+PVXDQG5YeROqCgyXvbf
TK2/6r6tKCmthajaX9kda6IvFqGZmn2f40FQYJCG31gT7M3a2/gU3GBPBFqIq5aeKM2ff9cAdPXn
EKUlMEJS+N915J1oGiSOWhMDX+t1aLmtOSoQqOmOF++ANVZCXYDG5YIAjuHGCV9hpF4b83J0/lga
qw4tX1azsECTomgzJPOUnhLeiWOF9b6i+tMQP7vvh2EMJPZvmg1xoixH1wpQvwmeap+ZWFE5AkWV
BRCrO4Qg9Imzt1JnWBj0xR4Tdlxlypbdt3uynJVqvrHw7+MaSKuF1pzBdg7dlnIx7fxfniA7ugr8
yVzVq0ShZtrxXuKoZ82mKdlYZbkSAAryEU8me0+ocY/vBRjzHLqeT8vxlC8ydkpi2xtP3xU3sp0L
Ila09kHilr1YDvhFvzJXf824Z0WM+ikA1XiI40VkWSeeMzj2/bhGVhCmvG8tAcI07lKd3dUQwpEk
nW6S9nBHV4K0Il8YVgmj0HKypPa26Ufachy0Y28Z1pG+hJciapHXvvE8OAo4cFmxV7jQ322KfH+1
s5n6M6NzZWjugES5PA71tfxNH/RX22AL7iNQJ9jQfTAuidTmA3IvKoCfrK+mi3MFZGV1CnU/1xaO
wTZQijAU3cY8bSu1daf4qxy7bnDQe1GH9Hy0ywdKFwkNtQjvRJzCJotTnBuQX3MnVwy9N0pVWKVh
2+Ua7nvj0mtKHi+kHNjoIBaZbA5HGwnaWrY3joQAUwBuSPhT51+puQVH+Mahu1p7r/VDi7Ycu17z
Gkyyv/sAOCZfuMIAj5tM4Uv3YU0SfEClrucaVRfOEoSwV3nXDlRbQMlFsrf+J5QNh+WPKTYEn3f5
fFVZ15pL/CDA57Lo81ztDNbdtZlkGBHmqjz/pFiKuDVib+/nXehl4V7IOLUHlyCIBo+gCeuWwB/+
qCjuZecbAYz5u1rnxSDqQLADku8q+hWqaYI0UzTUv5ZF4XP3ncB3LzBH5ThdcpgIySyt3PEeR1gM
YMIE3+Mx/FxF/t64cXPuT97mREV7pm4+i4fw1PJmzfVUTQ1fYNzTRkKgRYN8NNOV6JLM3qdsQG/q
CSd5H3GVGx0ILQwKWw6LArrijfj+lp84msz9yZhSlcS1sEAgNpO6Ln+9h6RlUp2MZnbCLrvKoeGV
kyAwCqmE8emj66ohXDyhat3gn15KIyiW72mhui/BzPECgynmf98bLRe3hpl9irRgosvO6p6SE5PK
mUrJhIQVOCY4FUE5fI1AIjxaMcq94J+OK7gtT7mSHzZRKsKB9PMtxGyjmzP20h1PU0b8yLwO8qVy
fFtRg+6V9GjkQ02EiCXnOP4tDieEwOJpazfzR/eFj3rH6bGpc7JBYVE1PmJZGEmQTFlBxfSGQMvn
hphKqOaaIO0GN84/Oh5yFbcJA8PYaV+bxO7vjNVBx9dCSKae0oqkcZiGS7rbiqPUhX7nTyyWfz2J
uXyloPtZBnVc01l/G3VfM5hx+r3rggFOAtOUG4hjjtC9peUYQGn/0ChzPO6ksgiHayiNgI5Po1CC
aPs0p7GjxrVkrt11+hQWuvjQLisYV9DaofAyqw0y2r9aiksgJBONSu6d98GroQBVLJtc8x8MHh2f
SQ78kprMwdw7rsyTuxNq8PgVij214fwgzw+bz5kfaAWRMSIFboCYrcusO32j+pPPlh35BpWT564g
ZHZbXF5NYaKi1jhtQg3u8LZu1cT8ohWija3V9p9LnfeJGTiHMED8SxDQv9epAdLUsvnbF8/qCUYk
qhMz9A+kMWrewHIxoeq7v8hm16bilIAuH0OIsj9DPQIpWYQd1ONgDWwm+h/lHaEaNJluTPVCpNFy
Wm3UrTQ2DKCMzKt29NiFbuXZSUqh1wDVCIqHMu+ebsCcY/dchT/irdrZ8QD9oY8mnouWJniQromR
Q8qzllB8PCRLEuDk6u4i3jP1+Bmghu3bS8xjegpm32VvsQgkcHHAoL86rvu1V2UO5z2eZIut6x9Y
tqdQ1o8vim40fBAYZsviIfIK8larMeWyIeKsfB/ED0ArUjXjJIW9DyuJNlzK3zyMJex0YMSb5arC
C3SOyuq6tZEGkfQX65/bJ6pM8maU5rpVEbJHvXu66pYYsmVOH0mZjwsAmSnYVLJ5QZuRc+9UxpMn
0ix2Ig7u7Pycbi/qRpfnjhpj40FIl70f3hg0COylhMHV4UKkrLyEgGvPOfO/TuL1jp01TuZH3tu7
9yeIhc1B+9C6lxuzmblkARIEqy3RMBfvTcgcuhMEkRcZwtCMllnzlYEJmAYvTYT+oA1mhkWswJZ7
4G8/exgY0LLP4RueiOsWhKJLm5JCxCopnzJiHlMabZu7MLtO8Q5XHJ36648EBcCDeR16lwn0QKYk
l7n05c1+bKXDv7b3WXm8xE4aY825gndX8z4llRsF/FwMH19hYJYNhf2BzM3Xx8Il50dJm9YveewX
6LA7bo7s2funL+0YZtWKTI+Q706TANIFKw0ZTWR7Qj9zmqkeulEyomK03TdDA6EI9LcJwsYmQja0
VfeFxJ+CyYEvtMsxU91BV/9P7zQrrVZTTHEqxvGmhVLhYtsvNflHorRj5djtE6S/xdKfuqima4M3
kS0MgATjyJSMhYlKZjOYIuRBzcOPU8Xysd1dMmFmkiLyAdipa+Fmh4EviBgu3elGDq8Xq1CXETcx
VgzC/vZ40Z/DcuA1eSXKR5Vi1b/3B0vBM2I6+U48Pd4qf7b290VXrKaqS0lbu0GyDGKWd4W95Zn9
xugC+/20AZFpQtxYNFR7SnM/rSibVFVHYPHeeuLIMTfqXWLmcq/w8rOuhdaR7gVDQPnWeWkgS0np
5cCWtFjBWZ/z4umpgytXPS0VqqR+OBbShVciXwIjmdGM0f7sCV3S2onTDBPXF5kp96lOaUnNfK9Y
S7jDbRhYO+fAcgdajs/doWDq4FjqWnrLRaQnnpITjtGrW6SzCahGqeG0yX85EHYwCEUYhyqnL2N0
kk00LykTNDBoNZO0xIct3iUKFHjqtLxWtq2jZdDWsjehnGhGV93FdVNHNvtRs19azjPal6gJLMjJ
p8pxO2ovMLOeG1sHArPczes10bSHeyHu1TgkGmwfZBJOsnExFdB12fE/Fz1hIczWtdLBvzkqfq9w
5rRKzc4kSe60mZyZ8Bhn+7SDBLHS54WsSEKZN7vP7IGOtTMvwwj1OWfWSPr9ri3fyBJGZBnlj7tt
J03doYdrLeXpPAToYXxpMPObd0Y5RE3ZVVxj8trL56qHOCjSVFB8jbtT+MYf0FCO9wrKoP4Qdd/O
J7sUEStcZfrYf/iCSw84Hzb14/T2Q44PSdwWHGfPQ2sKk5lphSCyrlzJOwPd+Fg3STcu3GRmH61S
vVN3yvBOBQtNNxZ34Py0OrrweMUlxs0aCeqPRrwgd72MAlDcynL43MjHBY3oqOqp5dqq7EXnzWEK
9a7eHF/6+BrvbaeqPeODe8m7ENTW86XxHn7/bq6xdim+dSq5UJ+a+3T4X+wUJzQ6amTzpsk+wfjS
XHENgZ85X0hj+Z4W8vAbT9/AiClMHZUVyuyWWPLtM/jvsCZK84pxdvow40V8kf0iXgNk4OwVO74v
LQZ9gIr2e8KHMQLUZ1+NcgZPlOmda+bxWkaWCqRyVttyV2HveViHYMpExxNVtNjeZnoQTpzniygL
8cWT+Nyvf8DTWUPyvURvWZZq+CFwE1TbVA+MYY6gpaVA1GRlGUzH+uCg8AZxlft0YjAaQ30/1Vq9
dMyJNtO7DpHl8svqcg5WudvHjsqfc3dq23DcwHV466/mQRV6b7M0U2rZdVoBrZB8DhrWmv7mrXa9
l4TZqwfYYuuJC+0Edh9Y+sZx7bN/3nBC/i2GsWc9vTNVwdY7jut4OwJfUvwFmMVnimp5Wf/iBHBu
5uTTC7UWlS0VHXq4bKJwNE8MhJGwOTeqdxEmUTBAbbsMOfkmFunnrEXi3Pdj6StAKtjw2lC6DAb+
du9fffWJz03jUkpUQOXBhLs5zm/w1hmY8jPmQGFvyeGgBfRfBo2zpusgG2+WfhELffH3YmKWti9t
EkWxiKTeu5kXM4Egvl99lT9mgUZqs2x+XAnb/hOCfSNsnP60TIWeB6cAm5v5QqrE2Ggm7ayCMJva
c3Gv18eNXdHnZupyPAUK3QS0LFSy4YuZKpMVctgeewWFmVX1A6u9Fip4wVEdOU36GivWydRyuS5Z
WSmhFJl4M8A5ybkgNkdnUrxDDI2sSYuviTa9qfNjyA8SFH/SIpuu/3PGFlSoMQWInSPGUj/Evin0
FpwimOXw4Dh+0aZR3BUyZy76RaL74THibwHdlofecCBpopsyIzUfqQkI+VJWrxVCnU0O2RSyr0lv
0TvxnSbHXn0XGdkhfr/vVqq3HTgz2YO0UezUDioYmZtZVPjQK3Gdm8f0g/qKG2xgr/fwPEVIdAbw
ALDMLhUywvAGETQ9pq6IMYcgSA4XBPFPvQDIIKJxLNH5e+y2/rJrmQbopv22s9aACigWwE07rlss
NvVaifjCP6k7T9rBamdLJMrgrzzYE1Acs9oCD03G4PIDuiM54Jkv3c2cfui6/+lrOlNGgQOSbCRl
e7+Y8vOiPymLu7HRMcev4D0xhs9mWFRwf48QyOOv01KBtr7DxILyg8JJlwZjPf4Rr/Q/oFt2rwD1
1iTcnfu7GuHwXO3hERR2+QS1ncV8t6fKGyDvoUsly7bvM2yivng8i+BtzMjqlddFUdr9OIxcgZfC
MFaJga7BcWo1UO5xalDLq/TfehdVRRxlZYca0yskxfYTIKzrrLSpGFThyTEqRcxKwbWuxxcxlJWH
g733Kz5zFQpGNRg+YdSZ70x1svfEdfxiATWAZZpOM2YoLlmNb45HbxcQugBDjHGdxv7QoPEKHmFu
KVGFFpBcHF9yt6wzRxwZufcFDb2RVohXloy/sW6Y4G9HkZS9fbsQUpl6ZDBzsQKPOXXvCXC8vqsb
mFRr59+UVChcSPpd47xOXQjfp3UBnSGrcXc61fS5dhtVPeqNHsBQ2xK4jmsg34ylBtWuqiYjDt5P
ARILxUzBhENP2QlVF6pAWqyWPME1y21jFz03FWNZhrv+p3f4fqOKdgfowmlNiiQGpjr0mwgjIReh
4CrqqpDh4RxBvg3ljvRWBSw/xQRAZnVjKbojYqKN242RhlS5ElOlevIGw1AIjvtpMgilvRbE36hW
SErhMo+Sum4NAT+tpQekoQhN4GmAN4KpcvDyUkz9pljUGrR9AIPLF9Io6yXOTYfrwvELUCUrU0b4
JjN0BqMC6i33U+e0QF9rAkPh4T3RacOUx5Iq6NMQzaaDrDpJuCKyybdChXwULk6zHYzSslFedrLz
QvOyzcC60G8PVMCPFxbNMYtI9NNkH++aAYcwQm+A9fewR61bO4MEeQcgH17jIGwzdXb0dzqyhKSq
tA8VitorXuMBPoOXR4q63Kfq1CPvcCMTFpZi0B1IMvRrZOSOzXHbzAOujhVSXuu1U1oCH0wBvOFL
j4Wch5SREEW2A8QBpzGGGBRYUznVqTYETTRkz05G8A2qX0WbBQhFEkawx/YsSHgqPID3OA86z7RN
0c5t+ChCrYG2zvlUn2lMnmEAPSKnzOsQHtEM3JhG4+pg3l2CgPmsr0u8uqwRdHHdJLvAyP1nLWPy
WGDPjiBzZm27k7K87xa/xtZM64IyX7MIipuDiSs3J48FdDVkNRCmkvCM+zyoDG5WAilaifZ9NoQ4
nFlG6gKVmGHV85A5Xrwt1sEEkH7QtlMqngKdwpLlIPfznpNNbw8f47PHa/lvP9ze+rqrtLDOAfFY
kpV40JWoHeRbngme2wP/pWAzz4WTDao/H544HJCVnbr/n5C9BJdQQTESPc8A6rMx0zD28A/asljc
8QnWus2jF3BdqcUtFgmrnYuBGgUFbzZR/aMFe8gHAGvvV1Mel/Ya4wG/6OmvLbVoLX4OIvEO9c3r
nw4vSGRzZoOPflCldPfyMBaNQmkmPL2nQqgE5dPl0j9RV//eBiYDfd+0w/N12k9cJNYk2zkXuoIc
u9Z1/cI0IIkqNUMlJRKIojvvkOeRBug0O/yzhdy/IpY2TLTKbr/2eyxhtjn2U1kI2EHiLJC/HXXo
tQ/ncTPWD2nIygbS70TgmBzfo/BvV8CaUKK8LOG1sz6M0B4KaeDuQtO0qcZwiU9B7RipO13oTWwr
W3oN8hxz/Y1fYP5rsNkZUjWX0T4SBb1axC9OiAlkj4qnJCZHJNVsv278sIgX3J9JnWN4MY51PJOY
S01Ajm5IktMIS+Gzn1DVOr1HnvfpfgPUvgdrMGXiKetMMpwlYuTxQektMiiUaybwL1YUEjmnAOIq
kcaGWA2FYK8zZ/SFBAXI340sSCYJF2K9gWbSYF/UCVomPQB3eH01Wv4dM15Hqrt2Oz1z9gWekiG1
qc5XMUqkIFLiDZDOyO7mo+IUVLufGMEARhIeFrvi4GGd1OQT417esF3yIFHVEE7mgorISfwgLd+/
Y7cX/cQueRkw3krPUFCSP3ohhMf8HJ67F1xAiVHuxGTXd763vZmOidZmF2PZtHPrpZpIiKtXutM4
MAWjrvCmgfKiQ/AVI6V5hHkQSFBqAJXNW66LeT5FthhuoJ39Aog21vYg6XvGOdR4MQWlSsw0RxjI
qrRzmv1os8DvB/+sN7Z3gM7KPreGsJRGmjgtSHYsSSTcT2N+N32GNFx63HMyoHOVxCa5W5XeMHhz
i1n4qyrDWAcJtebt19aeh9+VC0fgEW1nXUxIbURoEoLVddUU4UUfZlfYNY1SwjvtNK6QeVDzXdfN
BCdG7kl+AB5ilTwOqY088cEZJVaYN62doUgVVxda5I35Zp8LNzobHv7XChiLV3IidnNhGVIo24Mq
YEPUk31TGMJTE3pW5uSSilSwJvZKdutU6xbvrJxSEQFWM5gkBh94yaIkmO+vrkX8tOI3Fn1Zqu7D
yALMw9ci1srYLnob5ptqaO/iD0eyoEG7TqLUo7lBp/3gce6I2EcXRLWaKh1+i8VZh8BDX9H6PFcR
F//HfkWmCIsSoZzTV2VqeUn52GugtV7KqqjQ3k0h/xiyO1EGEHDtnRiZSz54u3Pk727wXZLH8uKm
BnU7Z8WIdReMCmm8L88876gFVqM/yUS8eD4jyd0/8d9bFytW+guhEF46wgoGxHrVK3y0ABIMlAuO
mSTABw+CRUWQITXwdNqttcYCQ8rBx2R1Mt3AolM06+rcc53wyC2kEAOihtj3X25y4DBfMWQvT4S+
wXoDw4V+3cu4mriKz9+8epvN6ZNvaNOcYgSqdYFdJRgG9igZhBwM9v4p4P7U+amsetEL7QiJz+I5
GSJW+MCTTAQwMo0mINWyZjDbQnVVmBJFLyfeZUzZA2Yoddqlra/87vK39uWhQ8ve3+GVNfRo58qA
yMvxo1cQXxhWMP//bF5z1uI5psspfJBsHu9Zjsn9N0+7sWVNLqfrsI6zV/6w5JmvB3QaiDFWx0AN
lHVBWgU/fTG2fUZXteQtpvTWmqVnhMEdGpYfwbKKA9BA9DT2Rgx26wntYpAJcWoAQQIp1PNJE8dk
st8qgBlIPMPmOqpjoEw8/JI+roxOLM+CoZlAz5NGAu9yvsEO11nxRLSNXAOOFc4aXpESzs1VBXSt
qcdQtU798U++scVeXc80+GpFlpbG/3dhu6AKngr+earfKy5dk4VSJwr1wxZLrxpwjG/dWx8P1JWO
h99riIz39noYQ4YZnuEVDbn1ic8OpkoI95WawXonfRrLZxxOVdoEjMBJkFqWhV/z1WzJkdq5ykpA
Vf5bN981Sn/60zSQ0a4UlM7nU46ElXvEjBsbA5XgVRtHQyxbXEC2s0WkbTN4lHZ1GKRG1YxHZCqA
sb4y9o6x/cZ7cM4dk22dECaFlgGzqsqeC9MDTacE84Qt/t/JDRxk6uWLVx6VHNLb4/w9GDPPRFzo
ctSw3Fow+zHlpmy3sVra2xXc5gaO8nFu3Rdi61oNd4Lv0adgGxmEFYqQa/1xztH5BLgi4VBSXhXh
zB468Y7HCFsA0nkJyPGDKDVNLfds0/Xq48yeYT1E/HDw9kHuEHL3xV7i8DwBtKfH6RylYSElKLRf
5WHEUe5l2M7bh6uwmLjFnBwpHjkogmWshOcNh7NQWX0E0HnJYGI9tURblJrKV/IfCNxHeHyNgAz7
HuxuSkh1cOyivLaee1IPFhlQ25caJe73vt0bXmGxLlNHuoBvjA0tJJbdsGPbsK4D7i9TTOg4zqLP
h4x1U4xjhUzhSllnSOx7dxjlWrOImUzGOSZE7WVD/WCuTQuS7noj5YKGqvikn5hhNamCxvs8kl5Y
Dws1JydlwwlMz2QlJyk632TwwaocE2fUzwpZIl9R/KXG//dwCBYOL9XDVbEFWwiEFAUv0CJ+5wLB
xgHiKdOgbscxydf2Ft+ByIix/vSTR93Dn1ODuvWPNEQWsB6BWMx1tWgnvek/Olmw2LVVD8gV0W5u
3RL0ZtZu9i1tvills9Oe4bew+Jx3xVbTGDujKUMzGMk1r6gApTbHx8v2MLge6rmVUTqJPsGywBTX
IYE9QydwczW+U+4ozmgg2EcxuyUjM0kFE73MQi5NkNLnZXXLqBDGeAhWzKaAEvU3Hdgr/bg5Yfyy
+pq4jjTfbLL54Wu9lzKXj0PVXXVFIAfbaRfyFN2SigBEh0XaWKW6ZFAOvsEHj0XgfLh8Npg7fYfV
ZlW/vPMTMGE2IxAEsIGAghqZPoMNsGnUOe4EroaYwIPOI2bs2+/WtIrbzIyEY7L/E826zLQZwm8O
4UIWJF6Jg+GAyJQ+pIVJTxnJmvd8Q949MPDgfjPlxpIttIeAfcXc7zhfeI/x6SciMKT0NrjClAOm
qBOTwh8j4x+mSR2dL3hgSLDAEmKzK9AwZ9M8N7qPAfnnBO5A9JYCY4mqrNX+6vvo7fHFbZV4QRHK
UTHnWAhMffCaO3A+XocwH32ykitSi2d63Tv2onIfFG5CM3OgOToNGND6eIldvE//bENgfGcQP12r
EOPqzqdPKHSZ7wyRhDPbhS/FglBWbq9tVJEcu0aLxsNdmS0OIsUE2JM4/zRVZzh820r5dpx3SSUi
hgLlJJVmURxQJr/Ha3QnaIBj4MBNEePCobc9U7DKMNHhiHTPtpBrEcXNguEI9UJz8FeUS6hBBZ2C
F0c7rtKRLRk6A7ZOKcbcqeDxkd3k2UaVisLCEHQ3V53R1k3P0CL8vSm0mYH5/ONdKgfPDtWZlH0N
/Q3pNOv3enypV3vmG41xCxgY9+AGb0ReXaUEJTHuwOeIS4Uf+SiMxJPiVYelDa8e48GkgcH09Dmf
I+jEmsN7oKvpTpkxL4VrHoYn3kPpE50X7gWlaH881LAZBSzMQMfFiD3wUk2BnEkRjYVtEWC5xHMa
RtrTj+M7jp5dU8ivZvx7uYhIzFImB/QNPy9aK1Fbl8oApPOBw9fDuJcfqK4hCg1JjfbIUT0gZJdW
WdVUlrzhVFk0NPqk64ZAaqLsDVISGDayVTSD0NbUOFXnN4WsKh4fa9ir/hYhOAc4QJpX9uwkenk3
S36yUCsM9krBqZZePkpxP7XbZA7zKRUIE1NtO2RvfZRrEd3T1JjWi8/kJTo/tCdg503A25MpALfw
m/22uzzM62WdhEB554wMV+ZO+FXLTw+zA2lxB2z51RsoFuo9jVe582dp8smNSmvkNRda+KBgxGXq
leG6aQleBkKUTuv7A5h1DwjzJSDM/EJdD2rFyZRIxk9twN5XM4PTuyC9H3cL/m4IC6snMRhuT5Ex
4huzZxGQmQzJ6xnMWjFOsnG0ELh+02k7D9zzakpAYDHMREmnV6zjoVtxUviHWcoYCWMd02WstyOK
qyq5XJxzxI91UIAjwDDvpad+VaE/sJlpsdjTSfS9klfmTsG08s17j2WcPASHTfud7093LDOJHNU/
JtUMWPyNZnqjw415EX4hggHhIsN9nK6xupD47v1Ox2Rf6vRVn5W0DhswHlblVLvhWGM1IF6MUjE2
58YM5+hqQQp6ZUN3NZddkTrEUgyAfF7lrtxQRKx8Od4Pxms2YOqG9MiVRttg7BgPLCsa+rT255sv
NW20sxJQjP1tNYEeJnAUSYBe+Km/S/beq48X0y1leI1ZvnBaez2MngMUITDcYHf3upEcJ4KkQCoo
/nzKZF9LD3ZNAMhHvrN6uJyIMtpRpdrERuzF8wpKEJV86dqr6MKSxcxh/lq1+MGwG5pwvPwwql/i
zWzFplHtUXG8QRQQwlZCH48SwfbZHIQjqyOzgtrFBYCeKvhimZjyAOSNF4RzRmE/NQ9hHB5FSqaI
+b+EevQWx0Qg7TbWlfzQUMQdkcCwftxAvVXoRsi7OXwOZqXD4sao41RbRWamlJf6tU4jwNVl+psq
z0f5HIX2kdJdcAXLFC9IKcVYpg7BBXQAy7GCyY6gLi+1+JsNinsh4Vi+5wiYen5Se9h/KBJM/l6V
KrCuzUAPZoFUMbytl9KvCZsg3zuenxRzHl2H7spK3IrwC0Gt41mJEp3bcRybQcGyO7rUAO+PJ8aO
qDkN0vg7f5jrk7nm0405tHgQkgzOaNWOAQEOOQEFJJSOx0mHe3ZJzXbteOz/5PqUSH2Y+bOQpn8Z
JN/VBmS5T9l51OagrTYORtl63jCLzvGBgC4+sEeFbfB4kKP+4P0OyXM7zFIYEbxI/mkwAw/+/aLe
s7qiT7BPqbwRwy64UrqvuZO4nJ6kGk5qggqN/xSNcblF+2yMZQ+0GQ8Hweg+nX4ttj7bo58A7Khg
y1o0Q3/sHrAeQh0OvR4eX1Lle62l1SvsSxaazh0FIn01NN1ssLQ71WfqXu7dG475z684ACBUZoT1
loBO0Be0Zi2KteK1XfKyCwkKQMddlxFlkTxTPO7DxEEShs3wuI7aiZH46U350LHrbr2rjt7WeeJb
QJT719qCHGyM5rKEtzxm+2G4qKYsJKNKjb53P9bIUuPxDyp6b8Hc9I3lmC3/SyWCnJ4rxER17cIo
O8b9vdEKGFi8a9umk18fA00Fh3yhmCTtBr7QIVGopazcVv/0alZIokNVdtelFEwL6iNO9bvIsTDg
6U7NoyB5FH+0cfmayWf+uBshB8azg5q80/K4Sxppwy+Z1anmhHItqMvq+VZZ8Yz5x9KsPwlciFU7
Q1btuGI6jOatbirQ5n50VW04+2j42sOGHC+16gV1Q/pfnH++hm4SuJPzaGi2rcBA9szwM47FByhf
vsiC6xidllybaY8OikEgkuazycaKj2WlJ9gZOpzGMC186kQd8c6TjO9rc5sqGkFL0g6cZG0qmDjx
3aWiRdM+/d20h2OAlKhm7g2mNlgWkxB+pOZUpMNk9BxL2K1+SwjcPWnEXqyZYcNlIV6zphPBaMqN
wi27brNMviCB5oV86M2sPL3105/s9c6X0xHX936qVmdL2cKCht5ARtWz11wPatZvXC1QkoHGCJpI
v5w2mnOwhMVGDswzzxL799GVB0KA7B4a/7eVbAa+UkQxE40ke04SbwVh9EGJeshi7kM2m8LA3nDD
2qSBTMUf47UEwmh8/iEkD/yz43SkTnuY032JoYBI9TG8RMMNzBpAl5y338os5a7TPiyU1Gb17Obr
NKT1mmatpHW+UvgURNsbedozEn5zOyvNzkeEdyEt87RKSpGrgyMtuAPbhJP4LtQvCQOw4u51RtIO
n2hRXy3egl2lKRGL0yYjr7SbN/j9jim7okTiXx2oGs1s3zTCccnB+oQ3mLIbQT3Hcw3jKl/Z//7E
XImKgHbsn4jYID/Pz1AnCpZHOa1jtR1uo3sWBG5M0ah753TFNeqGqaSZBin4NuSj/J3gLZ8Znxu8
qL+L27tZWQHxtIman4AGdRTSUNUieE+f4NzZ3/lZdOMZ38+v87L3wsi8kSgU3NZ+thGD7h9vWgio
wCTw6Sr5NxT6fTH3OwwQi8i18MmX+KOrBMsBYxuy7UJOFTaUCbLgWG59HGGKToHVWzqsj6U3ep9N
OvKQAxCdKzaLm5f6jVS2DxSt4rX7iZW6as+K3is8Z5XVOca8Y4o8Yo45SiheyI7rn9DJhnmF1x7l
OXvpfMnMX0KEJMVGNTS7G19ZyPdS/PGl4+WVM/nKTfwizOgHikasT6zXBDNo1qp6dmGOVsJSUvQV
9TSPcD2Qg9tYv84TnpoRhIYT5kP5qKQEdINOYH1LbfKszjM0HB2pxyM1MAHrGmfyOEhI3JTNRN8t
Gd3TIY+T44VgUvz4oLG7B37X8W5SzyqD//vQUipiOIVBiRxj2wwzpaJAGOveZtKDrexilv6tMDzN
eeqk8XOrIYtdnSkUpZTbFlWdGVfZBlEIISkTt1A6+yq6Qns3ADdYe1eHV/PZEo8Fw9CP1+AV/oF8
OKBYtc/hcJt4o/5p8u/QjUd7e83E54BWrY5Esxg+8JD5pFQU/lb7FVjeu0ksWjYudJghBgXR7ZH9
H43VWkT3WFLlSP+02gjgffcqyXD9TFTqTujd2IzfeM1N4Sef+S1fwJagS4QFfUaK9/7DMguQowp6
wHUH1SBf0XmCUMcjbylTFvFDHQK02eb5Z/m7mTFt3+HEBgEnzHqIxKrVOqa5u/NiLPMhoHbMjnTD
tatjOVHyvV6X5y3A+DuumI0WnpVzgQuYbpCzL2AxF/44BNOslLXI1lUJmBWDmqT0Hdn/vNJqPm/k
ibKRfhb4OZbdTVk+mp+psWc+rugUVdrU3CvRZhu7cXiiee/p9amRGIENCiaccSMzzQJU4tt8jxsD
BbEzRtDjmNnBP0Lu7RyV5mz0efKkFG5Fqfq8cizH4wg/PcE+qQUkYRWVCs09ViEl0dVxBDdHX+vx
dr8mdJZnzqb+CnNyz8k2vefFx+7clWPEo6dxZxviGrJBZHX/YQ5NT0aczJ4RfsjkZtOZbHkCy71L
WBwNNBGm68qhhe4lRGLO5MzetbUTolMZHAVXkWSBWj+v0DBaamhxHQc5yBqzvz0Vco+/jMw2dP8F
lUtGuso38tEvN0wtrQpIW2ay+Dekqf1spSMheEQYpWu3eO7F8ebZkoFJgNIs6b1tLcu8Or0egOL+
nM49QmXLK1akEmnYVXMiJjUXHYuXRBKgv0LNHqdQvdvIyjDovyo2MD3yJMJd0IM1T1rK2yV4RPCf
qAry0cH4Apt/mpIS8W7k7Irk2X1kx5OyaqconQ1DdvUxvMYIbDy2PxqN3HevyJlTHZrZbrc8Y+m3
73nKBvHMIgP5fBc9lfcbIQt1EuBqlh/7Puq5nOgRA9LdsoDHWcfmdacn114QGvjcI9EMz77mpqdr
aK89YM6ZqWNFtSmg+CHGB/5GMiGCbgC9Jz+URVA0MonI+gWIp2+6gQMSKfk4pboTDvWq5HOuydMb
DjLqv+Qz3TuVe5AoSd1p/9jAUHZQUsmDP2gN9vP4em0jWnSjEPBDpMCrAQquC9FwjoXrlfjK/HV4
4qnXdodyvdYqq8ffBK1nO2rmD5+7jbXhbzOW/bI5lKFsM+4VhHrjFHd+tDeXLJMXpEaZ0ZRSpxFO
HImpFjk+MzCNaWsd5hW1BNSzo00X2AO0oo5Xx4CLs8JBVjfNU4onPd8mvbUfCB1sJHR1iyULYLvs
+qXRu/HB1buPgIWwcTAmXXKXYyqJdF+4wYUF4MPHNmmQDJfx5XqpuC3AFaBmEJk4L1qxnOZ4SKeK
cd/2NiHjE1wCN6qAx1K1tlygsj7/LgS2sumqaHSTkKh/g0vk+niVuFApl/ENI5bzy4qvKblzOeM2
DEfEDT5PGozj8NoqeMoeS5FNsBQiOATib0YH5cuCskqDVI2M7jSM1gXv3MqFpIiGMyvAPO8aCs4l
JM9DChOPxFyw0lIbmi7RMnVJokPV1IuiSpkTPQHRoU8SFXZ8MVvYRNt3cU1qN8KWaUZZP1TCrRVy
oZT3FRklKmMCCxHuCYLN1jst0vY31q1DFmkatGi7ZdmqBUpNNdPjNKAscbCL2eDw3zY+IHbGU/sF
QfjmyQSRVgL6A9X8swh8mlGmj428DOU/Ye9wj+e1ghgntyz/0g6Hzpe7jWBJIAN4sNjV3wP+bUt+
uEm6JD5T6RNT2vdK7E3ZS1IyCKvvOBQqSL4hLO1+Ezw1Eb+DMbAjN82ys8FLf8fMdWIQbHGIyG/I
CpRBs9gszEK1Zc6abisItGCgVkcbqgom/XHcfsljrrqSBeitkBbkBrr7rcAmchq5lh9oHDlaQAGm
Ts1ZFHLuQ+VCFLVOj8fr3+mhaSJHxscfLEghj1QnTwJ2JX/Ewa4xFGjzZ5ph7E46/AeWDGyGfMZx
fXlG4dGqwjKRCG8zxqGGkzjFm7S/JP4OrO+y+1ADHIPKuJQhjKGcAafey25EUa9JtFdKGUTI2guP
Qa7CU3XTdTzJ/5vAEogggOp+ZxEDFtBMcQ0QOiUaiJS8cOFAEJwPT5tDpwSuEKZYjGRoumaiX8aU
NRM7BH350c404rzd/PqtnMdIpmOQb6w+d0aQamv7UlqwZzL4B5l8kbP3gE0yav96qfdpUEAz0Ttf
PLSo9SqkT1WGn2fYej+aQOTQXkPENCzGHfe1kFPTwmif7namkd4H1POuj/6XNqrwQ3CWyd4Gc0FN
BPYwQnqb4GagWARs2b7HQJTwJOdCb60eXKnx1Poh2ylQbVS5uxoEvXZNAjooF4JxoVKUTWgWxEQh
+FApg3gZlDsLzKuFAM9GQCJDhmgNSxt4b+oJ8VsZm6cIvGtzG/0J+uJBclX/gQ2pxCHt+9lWcvPd
6G8P0T0DfRDdTFX5xhUTTTYQqoaD8xqGeU+G41zlozmYkanBog5wg8Bp0Ytdffq5Qhfb3bpo41xz
4UqR53TWdIVRI8nk7UeJYeiTTAh1n7cp2QCy7H87iRl5b7dlEZE2REswVQy803lrrrzMbCSlzo6E
e0pGYiwtNxqHdy8aJWlWv4NLASZYR02a1FPz3su+ZnU8pI1ilL9XPDXiIBACmroywNM5/QnxU+FH
fBtuKQPkNFZAEVmZEWihq/RoLBh8TbNgfCgm92AaKEV5DuTBQ8CiXWbY/NaMbqwJR0++LgK+Pg/Q
YzlX5JtC21rdNFJHHjS+9h3kWb3Ak1Cvw5mjVyXH1UQCHYaVWjsJDGicLlVGhI5c9JFwdurvrbwJ
8AigKaEKHdaZYflrquibIBzNEWmj2KuY92rxT88RatRnXPeE4wX9/UdEoAmvcIRQVoUL2t/mCs9i
DSQvA9fY60+FZ05gQe8Aqpxy35Q8ShUZXPsv2f/sv0BfT0pEoMioIUY1bRS3kdoCTliMDQBD/Te2
O348u7s5SPMMOaVqR/bEbBIZAWLV2n0pqt9x/6AjUHoGUbrhV/VGG+Vjt8bkp4ReAYiGGDl8zT5F
3qjiM3s5qj3WNlPYnhSx7XZwkkpNvYZjgljMvvYkJjtdMMYHPuzfshfwmWxdGVkmCxhMeE5TOr81
9iO83OZyAoAV0z0KpXZho76hdO2div5OwXaTLrJdDNp39euss9YXPuzZJ3tEix7ViDwqnqGBg4rq
EC2ebQ9bH+BJX3BbCgweeUCUQu6oUH0fH8E2ERLgxCFPyYJZLxmlj6eluYJz1l98eN1keUOnSzfn
2rE2da+BKIszvWGHsP7WIrDxALK+9raYRuZpufCVtRfzedVfC4PDBEkW8VzBuKe+TJX/DdtVfS9A
EYUaKD7EI1+bqNUX7vbyFSIVgpCpA7nTQ/czJu/2x2EymFgGRaTL1ahTFUYoH6rVPiqhUYouLcQT
xgrACAvdOTgALFSPps2Ayfill8f0Z+y/0dWEeGOqNlw2QqG+PSBcKDULGi3AoJuJKzu0dF7ov9XD
Sx34ul5wE7rSwUwt1Ftzlsk1V0qdlYH7s/ZmNRa+ujzudo6uf15WfP6CW6oAJ1IwPgm1sSPJrmcG
nt/IIXKeMkowYE0catsVsX57lYrZy6aBEwt24wH9ILDYN3orXOmvU7hB/Pz7y2afyGcosKAxlFu7
zLwDBEiELdaTK5zzjN3CpLKhW/CPLDl6vJf1HRav/bDxeujeNL+OUEIEfanFSZe1X7luTeGOGo70
fqChXOsuSyJIawVpxacGp+jmj2AaRa4G57v7zDPfzXBukvJ+6BJs+EKu+SmQ8XR4mWHRaavHKQyQ
H7NoRlNAf4v0onn+LxjpJSiT0MrmlxkC/OeNkftbCxlZ//uVgAe8ZGGL9q1L3n71tSoQW3Fr+k3c
oFw+JD/HzFAVJv9qnPpNKRlvPgCWSRPc/v7nWp8dufF0kC8FqWLUV69KFXElmhBJDvS/oFKGCrcM
w9mrt+4LWmVp/G3gb9SBaC2tjT/Wd+jX53F3h2n0Cuw04KR5L5Tzm6/fYOXh/qiRSW9fCVBx2bUX
AWcEyBN4eShsq9Zx2jKhbOX2d4qffHqAUxkVjJRyhP5F99gK5kPsJD8+FgZtEs0O0roLuTjEy+av
bhNewF2JZ7YolXmRAer6Sf5hKjdgu2yBj9pH58sLyig9aAHHVQjLfoCNHHyjfhZVUreyBPowNb6M
LDoimFDH9ZOUhTqm3wSKO9Tbz/TdbhQSww5ttDuFJIbl+UfybC2a6sbXjiZnjm+NColG6XFAyviW
0CNZjPivmrxFhEMBrOK8QxqMC2QEc38g1+qwtUVRVU8/cqVSmd48Fa6b5BiMFfFGNzy3LZW819oh
r0hxSPo/NqoZg+B7G19ezYVuPfAo+C0kkeZOHo2/hRWxIJJIkESXx7HhKjZKOaxBcUFKoGdQ2HpS
/KdXLGFci1y2lW0Mfmlsrq9Fc4BPpF9JmJkkCVvna8fyAymy1Savil27raxpVBGu6rNY+ed7A0aO
oy7bOOnEvEcZlBint1ct3BMM5GGZilIL5PWePzVrsqsSsOYoC0ETX586AweYhV4tRcmugj1l33n/
6pAoLANn0I1+AO706ugSoVjLgqj6iouYtcg9AFFZ6J0yHj0Y8YSXXrhDcWg5pwUyZmC/6C6uj7iP
HSySiOe+qYwM/f73v/Onle1goEwxGoE197F69ugaL6glpagbKgfcsrOYTRjnJhu0v+Gckygdhf4N
cdppO3I7P5/40tkhSlhFqBM8bS+dUhAoaA6ShQhVX/TxCRqa1gJGmcuYWHz6pHBMlHt4EjJpT40S
FMCsQOkZW5klVeBCbWaBc3q80gIxnmIiXlwnnashkncp6rg3pCu/loIWxSICUkizLX/ZSHzjPp0z
rAfxFpu2bOcaJwSq8TOPtx0wTd9ds6x8GWWWPzAV+E5aLWNZrUMO3/rpSSdsexUi6ierD0oAg1yt
0/ELWrH6leVacraoPpBtoCq/x1vkSnFdsxp4oRzXvZhkUgdv/axK9ZFDkqWzuvbF/Ddk8X9EwyBB
OstA718ctzYV8QzimpY/SqLLTdqIpFMOQtSixicfbF4qWTAwNZhwTZQJqrgnQbz6P17vtNmBqxE1
PQdgWgcL/jkNIYufttoni/H1A0CoVUuXn6CHPMzMeQjoUSnsQqO8skbyAm3FbPY/PDhTDV89yW0W
DwCGG2DUFvcE3LvgdBWbgek4Gr+QetOZEGg1Ngin0Yhstc/mzMus7Dj7SIlJdZ8IxBGJEZuBhtQQ
ijTNLyv2qTZtCEG+0du82h6L3SZwYDWWUEvnRO7EnyoL4Y4ZwlQUYPRN7RTu6udsNcX7RjZrd2kC
qaiU+46dCmj8KcXdddjr8wrNo+d7p3V7NMU6VYALQhA8tEtFzeZ7gPmGxWR8Vnp723r8BeK3Etby
tpsFS1+jrMXphUr4/rU0jC63phLFXaikiAEdfPMsUlvolMZjxnaB3FvLZRV0/lp6yoy9LWgGOEJo
QJwFbx+HDZtjt8KM8SP/nVXQC1oY5vAMh26/vh/I4lfIRBr08/QKjbCwv2pvPUMgEzSpczrOkGzr
C8v/1C6tlv0ZXrVCSOSwbLVVRmFAuiZ715thHswUX+cFxWUekt+AYBLp4rOpmABzvruunJeQ/BZz
gvb5cDcsqlxhlUuBrtjma7rkYB2qyLVbitWRXRptYXCHlFRq6tmxZfLD6DF2gP+Ri+Bljw9Veonb
7fM4xX+kFqYIXsofxb4pqv48RkA8Y1MgYD+BttO2uYLO5ls7NFy772K1SmNbuJ0AILlS0hxPw4pg
6598qoQ1VzGw1yJR2UyQ9DdUkWghZWAteM4921N1I67z2mn6CWtW5tUJdY6UasVRYpWU4arX6+cm
lPcmNHjoOa+dnFSRbNfqBjHJAipwXRrJaI1SuqLsOYAR02R5OR69NQwVezADwejqX0KsPvKp0htl
O9iB4cdHl+G8UMulcmmmit0Y+o4JKegtW5+/xUdALxhpq123IthdB6bQPFdidFEaubkj6c8SzUd4
XS9cJr+ZYhjPHeHTx2wYBB8hAYn1NqC+MUzk8TtYuufKYSLtTUl6jMzRhJWaDEAePj5rU2K7ti8y
VgLrzewN4SaI86WyS2/HW21NdBqdeRDA3SvRKnbmStyvahO59TADRscgFe1HOiPxpIhnXUhoUGgg
adGc3Z6rQEyB/3WjarEHPqLu02+iJJ6g4uIBTgFABdt6xgXTOeYUoxGQ7xH9to2E8wYzG/Oykjxk
XM+JFOfG6KrfpugJ7DrE/a7YhhHBqv3UR1PNeZg54q2wCd+rGpbfFtkqgy51tKmM1MOMJTsJFLXB
G6i6YEhcxgkY2Bc3lfjJfkhLiGys8Lkgcjtpohaq+i2deugyqX0BTyd3MuMpDYJGZgf5wlRqqHOf
e3bCWGz/KyQKuE3c7/dnlkekxUD6mGrw7Ng6ETMsWr/mWkETvH8uGkXj52zngIk0k1POOEUsteD3
nVMmhWkDMHPr+r4pq5YVgJZzAnnRMuy+wWNNgufEYgQChvsSG92MjC4+ylLs1kY2o7GosmUNq5J6
obmHo1rhJseeUBUS/8FGJcBIyXe7nvZ+hsQtXj4vshyqQdGtaYasNUWvLm3kaFae6DBr8isz6r0Z
DBNFC1GKHbc0sDKD2Mgex6a5nogA9QdtV0h2bkKd7CO9AyasxKJn7BwcUWFZBVD2wTKH/mYzq5qn
sYoC9ltLnxzLZYg6ucRHehbw5uhPLW1nOpYXZLu8ngRuFkVt+9AWpCTI07ab+xEqAlNc+qW2uSqm
DQYmGCW9Qvl73uA+HpiM8Ghrlr5u0kAEltY57s93e/nbwnItrVQMRG74qNBFOcTQVdrHx/lLbA9V
3+qxv5/zWltvoxy8FiXNp9ZvKMRy5Nb3FeS4OirwM6qesXsS7IUFrC+/hBSJe4NcF1xYBoulHVb7
OHcYCow+bLDAbsjiDC4GFQanfJXgBvrHzDWmqnWP8cYw26gEgI5OHEFqlpm3KfBDyF3A+LF5dB9a
wb5Msg6VLxF+02IepcP8MarBu8GCg8yVWB2sYsfaGabfcLBFqGsdEM0PC+6U198pFKMEvo3tTsID
r15V7TL3E3WF8hjf7iygXHwEfZ38J7KiGhLeSSWDAzNnvYW2VqxNTzv0c3z97taTRvLe+V9j0BdU
G1t2QbWkXZjP5n31m3gOX4UnpGnxzSdQcFIs4775WozaefJ996qrJIOg1I2HYxgam1hMOmoN0hVB
iKlADN1MijhOUpc3sad48VNwQKz7LEc5TlII5zZ+16SZ05RLn0lM4dWq11ZCbehfj048scjpD+S4
F8gliWlZovtqG+WAYjEyCPlmVgzD1/5eWa4RKzs4Wv84YIuVmbTQSMxqJmlAFY68aUMWS0A0fBfb
td4l3UJs4I/RBOas48ZMb4VfltRwI5u4gb1TASW36W4kpjlOnjF+Hu724vdZnu/5wMF/lq0JhWWu
OjyqpqNflukoiE3rynILIK5c6VvgthQG+nAE2msImLKmldqeEpT+2Bbp3HS6dHl39cdSN08eQbUT
Gpq95WUmj9oAPENudxSv9xjzzlGf7AGJ0XUTIWcWjCuhvmbumvfEwezJj1bCIT6mYfLQubS+GPSL
G0/7KM5klHKOt7VwDQ9giAPbX1Eh2q1eeTCNZzOJZRVILSPa+mTQEC7OYsY0tVKeDveeXo9XZ9Lw
ywuvd2KnlOx9kn4hR1mHSUwHbkbr8XGMqK5xDpcrHs9WBoQw1MsDnlMcJSn9O1/iC00VaW6pA/lD
BhMWEe2s2ARhSEYUta3wEB0tU9NtEs5sk/5ymGwvIuStmd6GsoDhgu20uSY7u3Ej7IjJIkd4mZ6H
QeeAmImuKV0xiqOYlgcCSDcclHQii9bcO2afzYqf1BizQvQhC/iHzEu4C348SEQY2vWrGeTwlDLN
BkoZa69y8Q5qDoBDUWqfC90kuyl728M3t7TZ3rW6b620eKY5S1chcpIdZKh8YsOigaYeJWwdZIji
7U3HnXoE0GvYRGxyPu48dqL1Dm7tr9rqfLWm0LSQy7LmNTDdo3fT92mi73xnD1SWNeU+vStu17t7
zmVtsxaWGqQyX3yuVBFxHi53Tk4b7nJRLAKOQ7SzYTe15EjN4kFgRdJiA1rlHfb1dAmXgg6rJsKf
gtjfTIkQGD2wOt2GcuURP8evSZ4kBgxVC+LXgV3yEN/QwJZKGRin6Es5qXgudASTXhlIMOIjGUKl
/sXP4fs4+W19+eF9Cd/ypPuYP7r2XhHLo8tdBL2xZnHmtevBMPwAlWwfqyKtyuXL3XP5nZtU7Pgm
pmntqCrUj2/YtijUmd65EH/gHtUUwfwYNPiKpUr2lI538sDWMSWpo5k83UExhBJ7Wqqxgp4r0j1w
MUqp4HtLBQ7tM9pCmONOpB7WaedPi8whpz2eMd63vxfQJ5tMqNPloRjyeGmkcGL2W6RNmw02cyoo
wtSTKT2Kp5sZc5O3OdBnGRHknkbXtVIR868A6eXYCERjb+pGk/dIXOwtIhMvdWPD0/DebizkSzC8
xoNhcxQ7zEZ6Zg3jptDFpNhu5rqeuyGg1BN/MN7d3k1BhroD503AjuzIZDBJie9QNv4t2cxWxzCg
djkEtOTfvSvqNy7XHM2ZePjrWHzGI7/kOR/ToRR3GsNF9ZaCpKsvMbvfGQLTWZkQ9VjAKJZXaZVm
R0oUJb/M7SZAzbRXinImdN2q7cjh55pcZuFKSN5RtEVrdW9vY1Il09cz/T0ZjEBNE0u6P7PJUqLx
2xaLC8cZhpuU811HmjWjYANJWnctTu+sdq0Bn4macDpGJI5oJNznFiKTnS4zMCMPryF1nu7RhNDp
D5FuuKkob0i1ac2vyap7IfceN594zpCWdhRc06rLdoGxgf9yJvERg9YapsdRr4YV7QHhIPdrlF1P
tN0eI4C3bafXT38aj58A6/sRVp8bo3BuWYpL8DIZYL87o7pQJ/WE5UUzZpwix/oPnWQbrE8YbDLM
reI8kVeSV7RXF26T2afxHAnX1W/ED49xHAX7y5q54UQTFP+v+w8pTOcqOA/5qfiVuX7MExTr818P
8JQ4meGi8ymz7gTbV+KYneFAiIJAKnyW9RGdB+Y3siSMjO2rH+4jeMxcAJNm8wjBZHYoZTMpyn5A
VLhQuHLkTkUcdLZk8bo6G9zzHVcERznvCQxPXgwvLIeqIebNngb34JKMhB46iRsDUQodw+Xvgjep
oxQ5L/31pTZSp3nVATfTHD1e9PQOSoDTnZordT+kN6c+ExXNpgDRWggtdtiG89qmo3CesqZtiXKZ
yaDTrJiqtbJrULVYuy0sfrFS7ggvRUJ/mjnp2aQ0pyv+8exXznqQ+Xl3QwucDTHZ236wKhVVwcnr
W/SBXJMhBIYljd1zGKvwquboiOke8cl9yFFTAZv41SWtmJQ1TNZzSiCsVtplShHNJSCdu3Kx7S+9
IX8n+x2IX/2jfXPPDdI1GU5apjtx4CgtjYrxfLd0pJjJrrbgSCTVp3Z1HufPIjuPC4CCR2y1rDrE
n78VC1bzFU8NRCNS3+mrJC/bi9fUP4IjVh1pe/+dAg5rs+beAypoMxYNvnHrg8sG6zJTWmGUl7Fc
W9btfI5LEkNQLOe/t79WJrVzKDrRgZwGnbTFWsDUrXqqIT4YYZqNFBnWyIoDO0PrdVsLX2ZGjED6
5ZJQocgPC9Yl8XaACFE/6c2ZfxYiZXfK+TPCCVkEgKZl+DW8oostdw4W3W0RRE35ylElp9TMdTUG
hf3+IhXFFnDaUKZL0aAeseNUTr7LcVk3RqPmM773jsMtnLOdcyIM2Z4MNvyf9rkAsFEkd55efKZ0
WiUINILmu6pJ1nbkVGlt+omDHGowv4VOdQOHZUiTduplc7G0YAkzmWrmAW7jk93f3RcmkiG4G+Sq
3/qZF5Y3wqDfcn0xfFlwtlXVx53ByKR1H8giCy6CdZQcnykSnOi8MxTCdoFC6ucklU0I33dQBRyX
Pc/gmFhO4HoaKQBWgQ5hI2E+gDEUUu+Lu72FlZzmHBxDJCvCMtr+c1hRN+stewPJBFH5zE8+JDhc
dISGG8ZQyy3+tqt+A7ZbH11tdOECrFMxuIjY1lxgjy1XaUjPhygRZYgPEpiQU0QbPcZ7jZ8ZzCu/
7R4c4tgYZtU6kanhYifzljSPQxHRG9/kwKWBNYDSGZAgGLUOPIkj17ZqvoJ1qx0w2PvlaQVSzbkj
OFFGmPGJ5kzZM/BVWilOlZGaWnVlU81PF++6gzepnq9gd0PTM/HVt6BUina7R/EEDj1biOI/6nWP
sEtbi3sqqQ5jZ95L/xWparPNmnFPOc/kvCfSe6fJLEK6KF6EusHYKR3BPg5pJLfO0DWoXGjuLp1X
9BtJ9tMSK5SluIVg12fWm3VdGrlg9Qb47rz2MA6Ck1lDubirwsZnFQEbifJPLV8WyoXMK0Knkf7D
2X9NrP7crO2tjtKFXtnoCpaX1Nh+4ncYvIfNLacalR1PJCmFVanUQvcGM84IEu062pt5xePY/cgQ
4wXUfXCRombVirGGIJq6Eaa4cU8IiRVc0tAYZdTqI1SyIXCGSiDIp6OpZL4BYuZWY5fUWgndTXT8
8THdySWBiPrDBN6YSWTF8YJVr/+McDlRiXyDwLH4SUCByAsZurHPa+chJNj9VC1ifi2L4uRUuljx
No2tPPtLOcsh7mOsDWbI4YXDYeHORrmrN29e9+jV5aUjjKZ32cfHuuYofFpDaNTDdn4a90Qg/3AV
gIN/FfeLapuDJHt1UM5fvD8dHo2Bf9A610PQ0sLx152zYFVCP3wM56DYGWIUgOmI57GnOPJAZHXW
25CqJ349jvc90aggNmwbyQB0qidnA11fwCkjCl1FDSNyPFHhp2lOnZZmkxzsDzxqs4uqtuSuqXY1
aTwpvA0zmC8CzxwTT4cdYPEsuVPdzIUukO2hAXeOIVvzPk6YxZAkQdluwtUd4CCWO6vviPDjypy7
xH9nahr3SZyMektmsNqtMKrCUC9JxphSM73vwpX2I0bBGx/klHS51GUMM/ruEIj7rRKu6iD4gcMO
Xagaju0IyaflntnjtyHCjZjqLSqoTrIryykHP+w5cr9/7tHZ7VoHtVmasLrCNUVLzGOOs7ghIgX4
AMdYM0N1dGFWbS85o3nI01Wn/fgrZ2rYWPQl1HyplzBXBtIWf3oBOzZuGMiPmXQAy2zSa+o4nsqU
1NRTnbs20bLnbn6EqwzHpTfCv+zZ9zGBKroulClWsuffPuxy4oCjvMRUfslOXv0kuOOFMVnMjmPF
SWnoWcfHFQiI0wL6lHFyBt/DRgwc8/obhdNth0o002jFLcB+mGIZBrbsyqzoFTm7JpBvb/XZ1awl
RfDV6sNeuoGyAJCi9pqAUKsgnBDJZi4eciGWmBAHUExs7zZ+yIdHbrCTICx/HkXDkQq7OLuMXRiD
++jSPeqzYCZnZYciYZk+2uI3fai1H9c2+gm1BhDE5J2SVYqFoUC21voQ2VTrb6tcxOHi+7y9Rf3w
gd17yj5u1Aw0KU0gh34JcptYZbCX7PG2RFbw61HSXc3HhMZ/iH/VjecEpxQz9+QXqNLne2LjgdZT
2IAO2Kd+abn18furaxHUj8jYAemntJNL8LpcrP1B1lvzR4HW/3mTn+voTWCrrbodonMGarH7uuke
NUwoMPHHur2CuvgPVA6QXFGJVD+8y2haXHQsz87QMtaVbnBqydVA0Kqudos4vwvcUy29EOXQLStD
3jOCHeF6aVD9OByFt1ITxdYDBa4ir18PxZAcyrnLMocM/EhshOnNcIvEFwAXbkPKlZcUMWdu1V1z
U/XqKe2qpKRTcsIfnf4Q+cwH6bqhslit7c5ZHcMdYvJBplXMPnWhnZUih1Bz6xvblEWyFaJ3yiJA
YndxScJt+36bFghulkz8LNZQnatWYmTV+JCOLrxQJ/CMLtzIrut519/bpMjzjqxGBC02OE37DnDV
jjhG6FL0Rqds4XZWO2yB6DKdmHRaS/EgbgnmzQ4RnnRVkUOYnrSXQXXlYmonW4ke0H/Wb9y7cLnQ
aeDgMizz5WB5GGvtCpPBsZfSWvrrpUQfjcIhLIKWaMIteFQL6Jzb5yZyPt3B4zlV1pyHgWyfiwfT
UxYvG8LFBv7dz4n5NOnVoRQgtaI5uXDK6mHKEU7/zSiFB3GJnshYiUClzKnu4tLvJulMqKSH7qav
oYAvyxlAmKZldNDaHQfi8qzbJkeee6gMzQ5mLnLGC88b6mTx+tPGlOQr5KNDpcrz46Cscy8gxZf2
UnUxIcznn8gT/2ner/Q7XO5rVsVhfdvVLH6fLp2X7ViL7fbGAxUHBU5n4PWfiA36YsK+yQzXxc1B
RflV4TBzEIs9v2YzcftjCrACQP/qRbFIMmIgrXlFNm1VsomqD0UlOkijhM5fcP0uWx3T+4iM0fHP
AayUieOzNqk8unLhVnojVXbFGKyn2olFUzWzQeWO5WESPJPAZKzi15Wy6iCd0hLrLYeSnRnKkupb
VjGmSXMK/vPtNDo8TIRSGUltzT10hH11XN3tU+NT15KDQJ9wmZ1ngZUVwLUJI8K79z63j3mkpHq6
EBaY50gXgbLkFF5G3a3K4s5a9pwK78taIAde2GsgjQZ6hSlOE+PTg/I19Ts1W7hidkjdB/nsT62p
SFkD5ECy4rH8OrzB/TeOEeJyUCvrZH4UTjcvLkutSQ+GyOEM+O4m+FXJ0HVooOACyy/c6mN5eLFc
fEFhctOQh2JkMRM/XWfXYEPflbMBIVxLLZKOtZOJAyCKrl1ksuM2Gj5gwVuZsaMvFSdKnXWODu44
jf5ssIYkClUGBgjHuFzAEAiHNwDINx4agtqOeB73D6TVWSckosEK/T37jBpLK60Ddw4ijP1/zxJn
0NMdA7kT5q47b/kzIzgTqvGLb4sfLSX8MdlkIKeIS+htUdF2pfhuFYe4gNMFsW3s4cxv8z077TFy
rmxppBRSeKA/DmEoYousKZxgPby5FfEBguL9eJ9TyS5EfJV19bmWGr/l0l4eHvjiKXwrjCWwfYr4
40UhZO67PbfrqYeX8pW19OGZowDWS5mkOScHvgmB8IPc74NJ4j9WfUis6I91UWAbnJUrC31nJwHH
tI7GGYIU/5Wo3/DvAtvmo+8NejWhTwyS2bz4Xha24rbgpGW7QlfyLx2cqOYWHtIN7NVXD3xybE4T
TLhjq8v8q62LkI3GoKvc7UeOWPBrx97SLo1oVSJZZipTDPo13L9Sbfdz4PtFtfB1cxDoonA5VT3G
vBXugRosRrLHkbAZLEeMgQnyaRwsUDYEOaYckIj6ARz92vczpRsyehLqPWd03tCg1u+tv0fWICHW
6BrTaFtfHvYTaZXpCwCJ7t0p6ydGR/vUjwOx2fHDL/fZQ9uy4mBJ3fGCPgMpk28Z52kybuWVhMjb
ZARVaMmYijVwtsoNN1S1i5UPfR8HESoTbPksHF7OGYGtCd7GpBN/HdEwt5cHpykwh7gNnvySjG6o
FiUW0uI9fI2oretUuO5/Y8cH59mBc/GdrnbBNXhIb1fvTatpgPJ6paNb0SqJC0jtDL1zXVhVS7SX
icXstoJXUwQgn22Fcd6nAEXDh7/cnLQFoEJkIVNtWx45/AgMZ9k6DxOWkOL6+a84YJwqxfNRcYyO
+t6KVt6WCffEoyOCVCHT7R5mGHU5Vbsq06qX0naUl0mb85mkyJeX6Xv5y3oJZJu7VHY9unH0jQJc
KBcFlyfIrYu9Gf+Z16o2yUJNADiqw7re1U9QOykdSX7MVwH1dPpNT3joUQMYJl//ZkNrHr6L1O3J
mIyd+f1Nl45CPF/vav0nMxecrezYd+45RlS3apqqfgIZS1lLKymVXwUSgzmN6O1WFrd8Hb39vx5d
vU62Fqcn53yk1vjOo/KA5k6fOk6OF+u+3Lh+9SvNTwC+453jFNlDgC7LPqNNpTRapT8/X6i66rij
P2bvmQE17o0UP4rw62elgAqh4WF5iBe+0dvUPOO7hKgAbjYSahDBbYc0ZYQm8cKHaoJC2tySkXKe
N9fJJiiGyZYoD8qDpUgkfd4TuzTRBApvdr2yo0ifVHfug3ndX0MhVcE8p6QPxDUpyKb+ahE1AjK1
Qr8qakztJv3dgqScElKvCxFXtblE4/yy9jU9p8zRMZVZIiKEIPvQw16ln7ViSQ8Ga7+qIMwITk88
QmS5vQlXw8dj7xhq/UvvSwB8Y/yCaNpcb7pgVwsAgfBhYJXSee+G4obz0Ay5mjTQTkIYGCKx/9NZ
CbvwyJjMdNVg4c+IYYhn6Md5K3r6RYjLy+oErnAFchbXHZJkKSTvRELiAjbXAcr8Ncd4JgfRpO9c
XnXZVjNbHe5oQ/lH+Kb+0BXAIH75MgCGaKA3qL44f3RpGvPqvpDFcRoq3FTmgWTWI9P3qZRdb+To
ht0+qX2LpA6thxRQ9oCyLdymdB16fQ55P5kTjAsceiiU8PjUCs9BwdMgYy51w8kl2JeXurAdYwmH
TJU0oiXPffnv0NFtIjpUMEVd6vNkZQSHtKtDwD5NGSnFrJe3CQDmA+IzhF70S3hjzZYqSp7eD1Di
ij5QijCzx5BUkNTGpsrbpqros0RI+1Q4ylxtc2WiCVZKwW1lAayJz46Vs4HXXvHGFgSfb6ctpCRw
m+3/5i8qMrdWaA6fTusEhCXI7Q2QU43eRGfUGR9MO1c1RVBw9D7B4LofMgzpIba09j1blRkkNqZs
9L+GZ6YiSa4TD2FV57Uv/4BfM/jI+me10usunaJpbk9tki6gSXjZDgUHhVAhVr0XmlnkQxpYsqde
wmt3WUQrKFssV7uwTjqLxv9lxRgj8AATMUIHNmwUmvo8a71Q9ChxLvNN6IP6HpWGptcCfqieCqK/
IKjf039L4wzNxaxq4CxOKm10Ht3gbHs6MxfFn9ob9pEy8nM5mbDXD3o3Fh6cfmPBVENP4auT9RjL
QQMqavakpqwBK0u1w2GHbs9d3vx+tl7ZWgN4J4ZIMqMkBYhiQYUBkiqvYyXJI/4ewQw+e39Wr10O
z687N/p2Gn3QJTQAlgPjjdt+KRKcefrpjsb552266D86aqVdnV9GemUqcwbdKdVNDIQS/F4mKO75
L+dATnumdK/sy1l+57/FamAyEDnCqjYPpR2296LfE641sAcY9I5U2u9egCDSGhDUYdcycXpIDYLP
qi+s+eqVPdCWp5RAS5TMZc5JNKuaa87yp1kiYxjbWcuIX8CmZ240dLsRktkZvAIF0k3mwHa1uo1r
+nhpxW+fmMkz0bBNvWE3OJ4dS6JoDvo0ag1ZNfN8HPf5g/xD6pBkWP16bR4MlOhxhxyYu++Za8l7
0l1I4sEKdLfGKbupvp43/k7Vy/KHV0IEa313u3tMG+aUotOMhAQdZ4une+YmHAKHt4EyCxN6c1L1
vK3HW9e0hjXjZNfIUDEmm1B+GhUHkdLAlSlKy+usCDC4krWxxYRARjod42afyQ+z+Pq8R63JWpbT
KU62msJEMwXQuzMDsVcfSG1s9TTl949D6hs7c5mHzcP+41zp4oRM+0yqY0b7i/c82YW7QHxHDiHc
Hy/gwUyKom4Keor2kLPlia7cl9esuQDN9/Pma5NYqbSSw3GK2EKKbl0/c+ExFDMIV0JOqcQMrTg0
Rq41xmJUoHB/qzxKnW4uRDzxU7KflOqbDKf3BT5fo0j4YIgZs3WUlDiENdalnIK1Ys3A8+ASEBEQ
wrwcZ9h8oGbH4q3NyJv3bfRAlV5pSCNXhtLdVvlcdDyDVLDZ8CYVb4Gyf6PYwgjP3tV1PFPlVB4A
hCG+lo9no97qH3dPq7AIIiAu9xH7XvnsNc8Kb+qYxfZVkr+I3vqNmYPubAPuiuiIuStOI5iiDKPI
5sqXyb9IrJugvHF7g+prSxMNOtuDtnpuXb0lLM2QvPTnjMyxUjJPEWmUWXKJscIvt58thlmJvuj2
TESAaXC9QE/0Tq1Txrcm8LNS81z8BMNjJcOj6LZRU3M8A53004mobh3TLSozqamzf2jcJbPcirXX
+bX64WSG9af2z8oRuduwKaw07fVOL1OBi7ldzthyEirVX0aOBTjnMFbPBkMRN16ZvrHfudlt4QFY
iOs95RYT/rqznKStxia4U/H3Hp2Ho6I3O82BMSb0r537Iq48aubH96V97tDwjYQCu2YK71xamw9N
HmpJY6o7LStqoKxNW4szko7S9RC8n8S1WwRfxRqLcIWopdom5Jefcrd6gv9cjBJipdugRC/SsFMY
fW8JgtTEGZ3qpwdFMekXSLy8kmRROQSdH1U4v+5cVd90LbvVSLut5SCb5fXe7Rxo9KEOK/YFOpA1
2+ZEmZFlKit4hG9M+MGBSe3ivQNuItF0O6rdTwzuyxLPRpkdI8mxBUalSltz1oFnI3tmxifn2nFg
Omr6jALlkKAZYlSyXBIKQN5GSQ3O4T1dEJPIo7bPCYAQuFM6ConbCvP+uQUAucW/NWH9N6pNCsIP
oRpL+XKQ9V7Q+xSfjIgIPzg5afhTSCqCkVRkxVmh8EYwRgJeXHPPx5Ij0Ld+uqF74L7lTVzNrdR2
7UHNJczYJmjcqOj6neQSfOp1pgaKW57nnBD457XyeHPG06plm4f0Fmxro4hK6Sxk69Zl/qMK3tmT
zQyshT0+xKU1pKyBLozMs9EvQ+69pRj3SmgeQpF6pJqWsSOdN6TfqCIwbPOhCcMuHujYdd0HjTId
wN7bCAbNM3lRs/j5RYozCnC72OpLpsVJP2ShFLGYaIta4GRt5RBN6Jo5EV1ek5CvrN/TPp1ID5wu
KClDMusVEaSDxV1f7SPW/nQmWzkI2BSxVYvC/KJ2UmZksBA3a1MDPpQVR5wRZRSoHy8E8vg4OCc4
vfC2S8SDyLI7P+9rY2NJVQNFiScGsR4Ws0XI9Zg44Mx1uU6FbJUkt6Gi/8UplSgyBZlxGNKHZmMj
fTk6yvst5+RDcwt/h5kdvZY3Vh/4/LP76Mv36EnbWsHXIy7nWvplGJHxTuyiSyenKbsQTX9Zy/sp
a5iusiw8mh1724UfJsdb4zhZA+mQ0L3vgVdZ8vxjWPIsvLxRdRkRRL63RMz5fc4Yfo38bbPdRPkF
voqbJHDdIHgBa9C6f7IlLgz4oqiE4Q2iR9GHmMdEHxpJjWZ3jOUQVec8cfXDYQcHj1CSlPND+PmI
fPVuwED+KQvuYd8aDhiYR6cgRoIx8hPD5PrzSpdzMrsdm5RnA9qpXisq3qyVEmpPlvSzYCXDI+TF
wnD8Smb3oa6N1K44qaFB948N7JfRT3gujgS5IG21xZpwEOFRyDSQ4YKBnqomf5pwCnf0O3bluQ2L
afhbIQTTjcMQUR02cYjUIehluM8wGruYGJ4tabthrvNEfwuKAemOPRarvcM69SVb1OUHYLvcZeGv
d+o4pyg0/tc/a3tFAyXe8pcjW26HtwCx0w7goue1L0G3OgwGuB9xv6SscI4WfL307wM4QpQkls1A
rYQ5180qf8W1fjYvvhoBzZjT+ZKWSNlBMQYxMS4+PrK+DB8DSJdldh0dNjcWxXqus5OWar0bWnJJ
da8eAnyo2yiaVsMB0u6dzxNlPfnUed7Q1L3Nv8G5/a2136G0vIUBxVRDmSW1mWkkNpzylcQJkh9f
KL7fIjFuz8Z2u66FIojv03g/X2q94hIOJjPexcgYdA5wq29agfB8VBufxTFP+X3tpp8VVBZBsQ+g
WjlkM4o7S7LRwHw91nHeoLtpnMfQsW6/ns/9jtlB77cT3PSSdIkJ9kMZrFLd5Gc5nBI1Bz0I1/7z
cLx1V4pDshTs+FM1q1yAWJvh+5+nhWWRrTBxMjig50BTMU6HCNaCOCr9sStyzG/CBCr96iJHBZlV
eevxl1e21TX5A5ku22WrH8udQUsDcQPy9ad4KZnYdW+5QsE/J2VPRXXbbPsp0GAGEveHZ7fiCzJV
WBldKM1AjeZNBUefah+np0DciATFOAzKH4RMDcLS+4GNgPIVJnOZjwMIdTGnHTXW17B1XdZYSa8M
VceBUQyipsM5vA+7ooJNeZEUnoCh+Z2GEhzj+Eeom7znxleA9bs+5X4VcabawKXJ1MzeL8GH8Gfw
eRHlRCkyabkP3+dImY9V8likVOK/cRnXmreYRkscmUjpWW/pAoEk+WZUOzjikp1O6b0rBQ4sUIwx
CCpWI158YGL+5Uht6+nos+FDUyX6erbpUymkQj78miF3hHEnIOfNElDE41EKPnVo96tYfITjY1ht
Xg8yV2or2U5XqXYTohcALkr8RHoLvUh+uU7e7uPrkmfSs8gjBgOXjaWGj6z5c3c+N68O6K9J0Naa
fMvn4nashp1GHcwMq0qvGkmZ5kdIn/EAX65Ak1E85p2pgS1lMnxQ5/psdO1hoMAYztRsIjTpkzra
bN8j9sUIsCfj9h+hKSTkaH/6Yt83FxDWdN4itLgDuZMtEAajlbQzi8oFIHXQ++4IhabFiBhJA4t7
JWiW6pg5zueIplok3rS9DIVx3+sDTigcnS5aL/lk3nUA8ROtFeOB5H2BLHBRNJ+CcXwS1uAbgMoT
zscLkdqJpqBpRrv6o5wsgzLzmDC3IceLpStR2FzLlR1c7HTGZ9w9us0ICr5NfYEYUNCgGxMs81+J
T+MeMuAOwp3aKMSXOn2A+M3pCergCmvQJdXxD2HNLAfu+GdxbebFDEFXujzKJPgFf+nzDPakjtP1
6cp1ICwxr2WC+P0wsHoT2VQd9Y9Zfc8YhfLPSGrLkVAJDptdbeGPpH4mVGSOuJNvvSDl76GYvJmU
hZAODfBseBaMHszK+3n05hh5qZXveReWoNMP/5a8lrJReiDSHYMsYc9HVIyxYUbtFCJX/cPjgFqD
TJbAT8+Tjkqn/CedAsBtYs7dEFqjANDdwXRiwmpjhNrKcWQKcLFOOleO6qqVso675GHLNI2wlM//
zTJ01hkDsXPYWBqQROQu26/uJY4sLYxueWiO3kW/8EksTAKrMqYm9978aRymTuQKWAW5NXOEsb1f
ReX2q61Tn9FCdQUaA8bZpn6n2wLNTpRVTUjvGB5/4RXemboA41rgBLN5wsik+ToSE4rzml6v2D5d
/oZCbLE6BkWH35zFn8c4Om0rhZsIHOqaETjjmkCj0dEP/d4FcfJ7UzBHX6R7uEnNRiZ45jGzB7K3
mEehGPWp6AWsITHglO91lEo7QAIV2zj5w6HLoVrEWNm8T59/EGSv4a8eGV/vXsbdEeWFhBY3V1oa
fGQWk5pn2pFGdcvQ7Gk+jccCGm5CD4iq+J9iv3iQb4ZbIJVukh3r1vSUPHbot9wYtsOhqd0ANoHP
8+MFWxPreW38QhpM8EDomUydkhBrKU4or3zSoxX/psRvJa4bnxxxXhuhrmuVC6NkkMb8SeIBYf5u
RaJJZIjQ1UNM+CcJjuWXnGIa8hOTaKfhTvM558vwjW9X6hLCZIZ79fyu1jDe/k9ivZb/nnq12tpE
MrZPEVu7a2KYqvBJVL7W8rl8NNSJiSE9e0SGDcy5c59ZjTyZV8qSmFZigLZrrTCJ+LFhwhCMlNXT
SyZs6wDZyVVoi14QkaETbUy8RbVJ9Pc+zduMq7piVzOrNx/Cifz610HV1tlKqHYFxruTmpDHC+Sl
tdgPTrbRIL1E4uvBQmwUp33ZB1qldFvau5Es27IOdMGG/OchQ8q+78DtqzAcDpRYG3R3uOccxzgv
Ra0UZWGbHoWkMzgWGvJEROKJN5Qc3L3wpxKQM0sgEvglOC4Ab47FbT+IZlS+094ycw/GRhpfOjCx
HSoLUuD1AvZ/cEZHh9V8kyloyu4VFBlzedNrWf+rZOKiYUrd3XRCrhqKEIk08NeooYAZ5ItAJ6vF
Ze4nDuwXEqTMbKwRUngQ6URLXIJynUq8F7Gs7VpcCPTs9UoBvDZVuu0KzHD4lSsb/6tnmo9+9HSa
A0iVRBxoWD+N4Gh2fyT6QUAViAeYopyD6tNuB6Yr9FPIri2Jtp1YxUBzitglbHKWzWeHM0pM0Bg2
l62HnO919ouQdEP9U0Ghu4jGFukMlMFM8uu1W+DWhTcMCRo4bGnFodHp0yOv2L1ac91wvtedmSpL
FJY2A1j5wH7vjryWEGPq/aDt0shsMcU76MpYmsc3C+MjHHfd5GXtG4C/+gmplLQHZeIU52geShZL
or3exXjvz4nS3TUs2OfBwVxRDIqDItkee/7hcoPCJ3YFXavcjXddIgfNVbwsjOeAeNYrrVD2efsn
IAu9uGTGhzjkunZKVQ6ezE3QBKB1zFBH2jNxYxUgcGtd7t6KinVC9fWNxCPs39aoMppE0BTvXFjF
vj/wTCzPgPh9FrwRjtmM2hYQuYfOyqqWR9+Lp79Gdg9sYCWhKJmwyyRXSquNfN0UOeyytol3N5HO
N439kldeS3VmJb06g1Vh+Kd2os0oU3tSjIphLWbluddWnHfU5GdMyhwtxE4HKEPy+z4Bmw3CJun+
fqKPkawuCtYU5/loR6UCnogQRmRGE1oO6g7KO6aMpS+FJW/HepYX9pfMTCAJ8MiOYC9f9MesFEMd
8LyYQbZKZxrXRU42sP+ZDjWIbTd/XdaZYLcrUJjYtQLxw5eE/UUsncrCJ5GVbCoR6h2TxGUsagtI
jjJNneUP3wtlV9EQa8+SCyAXrXt8YL+Tgi4/p2kd3eDaRfnKwU63taqqL9IvJx1pt89btVc7KiNn
kpai9Iw4T1YnqhYzZJw0ak6++FQOs0yD+sIqX6AvbTu3s2D7U7MVFgssBisFx6VRXgO080oRoz3L
DUDlDxUYDPdIypUPHvzs2/3M4tKEPrG3Aa1f1W1MlPY6C9U8RyrqwTOGvJUtSZebuNSiHw2SfKmT
QyRp9t5bjbfX9ZX5xaM9lVq4MVKTLQu5+CuzAUEjVnkjbp/A+zJsMdKjw03CYdpKVBToWJ0oE/Bu
Fv1em+uxAg1AqwRQvsnEbIwyumFbjF1K7VVaVFNpYdu+Sxlk++9xMVT9vtE1lCckT40cGgnLD+O7
79TvKrkwhJpz3nuGery2DsLyCTv6HG2TTO2qXRkDG6l5ip2RoGl9u2pjPbZF1OPjQzKinMREWhsu
zMTMeo8nml1E+oqWl5iHujgX/8DIfuAsRf8Q8LHVXbewSSHN5+IWpPEz7rUEzJ7x0E5Fv+Mt5Mzb
WXkBvwZEbsczT+Fvw6tE7zmClXYY9oAgXsnaSLzD4j3MJBV9hMez3xJa7F/JbnI0zibcsngwv7Fy
ExKdagp/bbh15xn6yXRJTnqsancAQ0B6ZIz5hPbB3Ti6H0gab0PxY6aPRPQkqdd75Y2zm/9TX4+t
HgFW4Qn75Ig7fN/EVgEMq08ymI4Ow/8xYKyyGccbWL+wk3/QboLTWH8pzLVbZibYq7MHHR3NjON4
w1jQbfojgBeZLEsrBE8fMWvdmcySY8l3l7ccfiGoMCivUhAnazGUVDbx08qL31qcCJ1dRn36plGZ
HVel8Nv/UrF0ToTnVNQaIXwBldnp17US6MemlaTdy2D4zRPcpJKqBatkTI+zB2DaZhMOGYIP7Tuc
x0n/Y2slIKk+0nyKUSXp0sFree5c1psu5W1/9HOxQKokAEpySTc3O4n3lk2l23/L4XZp8Ef4UDMi
3PQqzh5glcHWmD2+72fuKbhV1YNEmGFGFf0j684TN7nvN7Yz6WQOX8BAajcDwNP2Dx556Vz2MYEq
ADEVDX2Jc6c99E4hCr4glCvmZfxsFEJpyN01+UIH9IqEtpiABTcm1XameDaIwpzoF36nr3U8eKIw
QbDImeIadI4mVhdQD5rYua0XoRzqPA9O67/43ChD0hlfACcd9+V5B0B57xdwxnPKPlVScixnvWgO
bJnfFNsCvLVk40QtT6HcGZCvuzQE54RpOr3r8vpvoYE+dYLCoYF5PYve/MTIz32oAdttMM9zdIac
U6slBV3DHG36G1AC8W1MlNewY7iqD2YZUVPpmtgcfOZ8+awCrm3MTNxd63r7qzy5O14Mi3JUtTVA
cotKWuwrf76GJvk3QiqQpFmyKKqDnnDFUtZLsfPiak1TxIucyKke1MiMeIu8xsbQu8id5JQN9sKn
JEWOpZ40mCGIDp1XC6f5KKMAe0GjNVGGcUJ3UX2C3m+bYBoAFYgQc3X9jFFU/DhxUg13JkXsy/Cg
j0+VeU3KNg5grXqPbEUnTYZsl5SKWBnKOePLMya16i9WYouqldz7aTjkXke9uNISBPhMpzyZGZny
wFAtQr3Kgc4ekDODTnkoyQuY9dj7jg7eywBhBmVgdwm6mwhzFbU9T7BsXDz7qJ1jbo5Z5pudW8v4
htxYM1eTqFu9t4DNy6SPMFEG6bdGjC2wBPRqR0T5i0+lNDySlZi6T9+PjV7WDJZQL9e3NOHoJNs2
uxepV81lF6L68K7NxDsA1MrBOCanfgV/usvQ3fTaFfSBlM8Lr51p8vT2lv0g2AYZK2C8WUfH8VWq
/qZ+GTlH5L+iOaTrEn/TBuHcnwmnZr60/K+VE94cOFF08pVlMzcOT6U3cx2i3oymQYqPjJGjSFv1
s2RDev6naMOYI2VHfNhPKhSQMMrmIFf5QcUCRhvhlfxMo8h71BfFazIOZRwSf/Wkwk9kecAuoDGO
fmcyUQVuQ53xzE6jhK0nKxAPGKnEMXFt2K6JRWjFQj/gNdwbFsfrtx/LBKgxy3dR1CYBLYR7uqq3
0l2xVqNnE5BHpatono7oSoJ0z1qs6rXDK5Kh0vTW2TnC/Fi1nG6/ZQf/xDcI2kFOnfQebFkwrXt/
vUEVD97vRCWFnnGFTJBHfksdzEWkcUECE1W9OzoKFDtT5c7BIKKpe1wcKXK0gxJ0jgeXKIOOmB1w
nf/RGJM5CrGa7OmlJ9VEWdpqJgPfqrdYLTNjFWqIn55B/ZVCRsKH29nAouQ7BLRJOfY6VQl4oDvt
MbcVSj6GO45RkTthJQ6IqR5pKTQSYxGWf7Rr3vU0Ka3qouBXsvPSKtOGLbOzZePg8FXpKv9LV/L4
clBEUTBX40MoEESImBPMfhqTf9SkmzjwLXQX4WDxmsTXf5ntNJqKLT51ZhwkatuHktYQSW7hQ3Sa
68JfGRchB2OBX/iAyvjkWsYh8ApbLeNvo6vh89jE/kYce/9Xw/R3gefzQfph4IPw+tKdzwe07o+W
KShyx/VQnkkgf5k6iqPYhfBMgDT6YtBQLWOUNvnXP1F+h67a6/2b0S5IYP8lbXhPGVBxzxckVCXH
KB7GDtNIiAqRpDK3tFD7zDcGt7qTABe0ygnH7etA015qk+g9mG1jniYafVgsV9vjPzv2tX7YFTfa
Z7JLDgpqhRf5OvwuW5HPyq1AER7e4m7xEfs4SKBn9gLWNqnFWi1A7PZNN9tM0SjIbpnAqQyIbkmI
1EvNcvzTMnJxPMPDgI/ni9I2yODqyzY9j1IVP6Mry6eoY+cm4xnHmCFrrEIh6Ps3QIBb2bky27bP
VWNm2YFw7/Vcr8U7YlTEYDkY5Pi0SlmTTX6pVbVVsh6/Qdbn+8MHglVXhGi5D6rVdvDEThiAYzBs
6c1imKS1IYNFmvH0lb2uFfZ698mSeFUV4hf/sfb5nzRhe1DaoDm/6KcUpekZHb+bsSwI/6D+4J0J
Y/+5hRMnX9t/u/PRskoEmRuLRjToXnAx1WRhW4/3agCbZ9dHXskEIqllo0b0PMY33wi4qhQq64Sy
FF2pJvV5lIdo754oNTLgDk3oxjbNGOYogUR5cPJLK3KvrkU0L3nqvyWp5sjKj5bQQMivyreZH1kz
Nf3gQjSJl/wxNb7RUDcomOxvT1gaop6Ev5VgqvoiX7YC4k+kNrgG0rhtu34EamdosUt0kpDTwjEv
ZCwU5KPWmNpYKSqiqFT/unCbY20jcOBoekRDrjAdqPlQEzyhQjYvFXKGeaXcU2+HxzRWzlBRHwGR
nvl7sDIDep7z6CEvZHM8zCpUSSKkNTBap16QO1gkJmLqFP5/kM26ljWfMs7dBqzN7ijDMiO1wcnT
myjcuKavqhsPNO7Dhm4PIOdbsOCvoQkFV+o/+G/H56Rsp0+GxrimedOODcMwVeHHCn+P+3hYJP/2
crhtU8rS2NjXRHsHf2pVs/w7taJiUK/R4f/jgvl9JGlUZWWOmn7Xx4oj73UXw1ysTvpEUBeidBpq
31uLub54ImfYC3v6KjKV0Y7HwspDwWtJar2vOSpuk5AcRuDncNLUdE1psPZlFtkxUiAx4W3jv3e8
vvysttwozDu6y7FLGk5zCQh3CykI5M5G7pv4cqLDXIaQctUwHItoGIgj3jahicZpy0uiSGTsnY3v
VG5ta3GCHgjP2qe1g7Of4wTOxwl58jgxs0f8naj3UEYYmMXpp/tQGHDC5rUHMgnupLEB0ViMI0Dn
xgwwiJpGasiX0VfMm50LE9pX5ksZIBZFHeeKqno+dpk1wDkEQqaxWaB2LXOQKx6GhSd3QA9Rkwbx
ZN7VaYg5z9DfWUy0hXGfz8EpmAEarX8qD/DInuqi9ktLfETwtegAPbfQQiPhmsOuEzstHkYAgaHf
Lt9F/jf4KsV9xtI9JbquoP+zrYgyB11ms1DXJPK+qPbEiE06URmnr3UCWQU4DwSWRZ7KgeIo5UmF
NhD/kkwh+L3P69cRqdEVGKbNghp/b66BTHRfy/qp/L2NwAKL6Q5DB1nMQXI9o3D0SkJnzEyP/rrN
9Mrc2SfX/bCZwUxCapFQcAIxDdHdckmjslMzoCbr/jxQb+C5z5Rca+vT0bpX/h1ADUr6hSv5y7yZ
XYtUVtBwRbCeGFyS1CxlyC9E0DbwalCZc+levWkbKX6zf2afdgzVZLD6NJqERr3xIYHd3tJVc6Zw
sMgMx1W17DpoJLK226JdSj42M1sfgrSKSRZtbMoE2op47DTk6nrhTAhVDgX/8x6sWuj1C9O1rPh+
iJixQlHhVqOCLD5iUoAfEYyH8ZQ33jFcgv7Umezb3dl5rFkfIuc5ibU5JPqDqejN7k5VNS1mI+fN
qtQLdfeoRWv+Db0P0owcJhv9Vr2XJLAuwLLVLEzrC/E4x8LCF4l+kGVCg/vCe+Fxsq9NFq+7jqQn
2y6g6r+ucla8NMGupKigbR0l1kDnj4ClpCXgkzAvNf4b42UO7HnLlQeoYzPI160bmg2jclG+gQv5
Mf07X8riyRc5RWg408+nqFLzoPEKlvj5tl2D2/UCrUUycLe+EpZ1aWNIT2dWo8J61DsWwIsnix0O
WT8C8Yud2UDqEXx/Rll4/nS3ctAIY1oFXEmwAAwOHg20/f+ckQ2eErS//zWhjG36Ee2PNXmbIM+D
JygwB8Iaxz2inOkOQFxcNeYEaDcnY3YnwyyAGNSzorCsrwGcOwvmulWqEB0aUTIA8xqIbkuQRjvJ
ziV/Sepn2phjqRNfKsluDmCT32IixDKvdG+t1elIJHmL54z7eqLtU6mHg9fLsVJUHfcieHHOc0vW
OmWV2J8N3KjJ6YG1LLzVYlVSxVmcaXBcF94pOTALvqZwQBQNUqap/6UPcnjPMnBb+JQYfSZXXwsc
b1jTBWqo03y7WnmVxpY13+j8PbTJgEbD8g/auQ13iG62W5L9Xkvo/3cLxb/ZMkUX8edXx/xqSCuF
ic1Vab9tNlsA0ieKKxvbUaA6hyaVuN6P+tPHdwhvTp3Cx8KpOtSePOj24GZvHKUeCMe9ItMJE37k
T7ecI7EoiiQYp3/Xm4kd6PJJ9sh2z5zVvIrKi4F20ocrDU151c83RInyJ4ahBg6Fnka5KDwg/H1b
eKYGrbA6+hH7+eRyAA8g1QODKQpe4aBbaeSmz+lzwypNN9Dy+D2V8YJpFBho28n3Rpei5k4PEZBw
j+2ceBhS196BHjuAvK9qCujGvkHFp5TJiK8HT8xiz8EDnGTEOSHp2+XoSOTLGQI67m6xy2ifQhBn
20rqB5xLRU3DXnB444XYdwQuz+OJSCiie+KrfbZiSLIgfZ9VmI+9IY8h6rd5fqV+4e/HJIqe/jyj
hD9YMTLB3Xtj4eBMO8dDhje+5qAKMWu/zUh1LLTRmUFCD92r7pVsotbUcoLBkqYw1FVzdrZPKTrG
qQlw7+LKugpOj0q9aOBgE1MXjRZeUb4+xFQfw4LvexpTKZN6N/QbZL6UAOhH7kUwn20pMJY/sOhp
G6+K45ELZnR77/pV+sm7dZuUsNW9fXxbunuLYFZIc0vx2Ms+5+krGjJz3HQHgSz74AHTHL+6H4or
kVV2ZfPfSPoNSjHeUAkLkHkEVoU6e7PklFemvGeZXF9zStmP88mR0gQvW5tzoPTP7c1d0g/1IV5p
/gb3ScM+y/Xf77aZDU5IiA9hr77/7nTBilAPjxtmL2JXDe2pbRFTy9F7rpVDKbRCOKqZQ2Z4u23j
8r2PXpT4jlochGPHQEKvDO3e4/QurxNSGt99v0Q9jLBuFZwgCfQygdehMr/JU4avsgANd8JXtJLr
EvaZZCuD3RYiaS5MCGYLH2dC5rg2yBnTyk3BUs/iZ5aoKQvn6CP0k7qbJk8YIZMXiC3XlwLOT+lx
esYqGGPxxYKNVNXQeYOAVyDZkvh9ACANq63++DwgfWGfwWe+Ut6BS1QthQQSVa3Wq36grCkHdk8f
4c5ns90h2pPxdTxVq0CvEzmzC4lm11Db9xlYj7hxe0DFT5zUHiOYrZEwY4/6a7e6uDvES2VOEKBX
zORWB44DkNhxmt7a/dAVLBTy5X5/VmwK7ECJeAokOQR4fUnvH1DnGXzv3EBbkMUGK69fNjozltPh
qCP/gTQo6i6+/mLmeG5Joz8puyp8JGLxCFJSmEeImHmpzhZO0mKTmYQORqhLVF0o3w1k5BwNmeRZ
opmdzwo6iw/WDbBEa4ibjSE/q7ba8BF9KWNkRTBOoNYZvtaGhlF3bs+LTaxssve04zXHLRX4YAOp
gSrwfDaB7BzWHCG9NxucMSnmfTJ0lV8XgNLEBtOrTecLWQLge6dk043oLFBTRtDAB4aYg79oh92L
MjSIg0uU63pWsr3d+ECG1UghCrwtKLD3FzYSoPOsVrZqRER4MMxCLLmFFGECkHnuBhBx+QoSI3JH
Xx5FrMHESGsF1rQtPP+CLyh0WnUCgJVIj7gjVpQ+yzsrnP/ABqkGWgS1+srFcSGiYk/fUEpw6mWm
HDnYZzawJ8Dw8FweLCHUMYUch1JeN8CSyJBVisOMsZTUxdlWTVduRF7+IjnrIOWwqX2QwpQq38d7
4dZnCu7dMRc7Boqdwd+xhizXxR9QWS+EhSwqR3T3JjVHZto8jFfYZQCXfUeXkhVHilRVdWPrmjPF
QCfT6KPySHf7i89B7yfUTbwl8DxNho5FUBIxQ76gnPcC7WYYm0IYKL03JNjBp7py4dbQiVnmZ6Is
EcInaUYXLGQi+jdd18L0/WIuJi078AR0M1g5GpaNr9/G+PjaoNKiyNMGQrIJb8wtQ1pwqPUBDss9
lOPOCTEzGdymYPZzajvnV0DhDvmr74FM1ebCJkWB4QSOTFT0SL2tMzpA/0zk2Nh0GL90gwbnIkmR
nrclXP6d1p+tZL86bfKp4eDWjFrQZGuM9sik/TqUvkIeuYlrGRErPp0Cf6eNCs7evoEne5AqVd0v
xdIt4T0o3LfXGb5MZS7MKdlsuFjZPg1isPRfbAJN/Aznju/NOwrONNYKGdBBc8dTDIO8NYGA4UQX
kEPb9LRqz5QF6Hj4T2Fp+wB3ngh3zEfPPceONtsWvVq7PWVfQihQpF/7Buh15pMNrvSvQ7FFya84
mzLnN/rVnMSX2P2GAxvCcDvz8/y+IfPbRbgMIqf32tg/6QedSsgewXiIZEG8BCNZMi54O7EmEXGA
uCqhZH2G51gDUIkugNopKCAYnb4fxmxCKQV6pfQMlT1Wnmb5oOiMur3la7ZMTn5M2cKOZ14WwiVX
x9bseCUN2WgAQAYA0IfN8ShhhDkujH4e8IflJRvhSEy+LJK/R4zufYDsrK8MG+343tG0vdjTNF0s
7zdCohqGxFnavyn2jrhcYdVp81svAKqbah6Sn6lH6XYYRckoW0A3LQkCu4QHxyPY+f/L7x7e7dov
XxB1dbCY+7X5PWStEj27+nNP039A+ma5VxQclL6KTA6MZEeVfhqQhcsB3KoWzMq/ldAE2Hw4p9pB
9oM8v4IgFIKml9Q/UzyHkkEmUNzHHnygPQsM//EC/5xw3HB3ZKq5J4fYiHwGs8VMBzV4GMO84/wn
waEUKLUw67YNBDoAaCx0rrDQs6dlFRHkINt0ayyztbX7JBQLuc00Tw6zk7mIMPX5U/HIznaw07v6
Y8P3YTjK63jHt0iWRMmEUNBO5W11VZPLgIkBZY0fdaGCP2aP2TGtdiqpXbQyFXyX+L5FAO1E29mk
oElgYp/0uyBcXRNXfEl+ra6raGm2kXkh/ttnYZqbsvkgxriJBWnDBaAMW66ADtiQa558hEohjg5I
5d8mT1ZNwKjclRjozz+0hPpzOmDL7BawS1jHGfi1Gx6WpK3F4zC/ODHmtWu8jQ85R5MnO/qctsvc
A5ShtotyMxsHz1KnFl8HnqGy1dVr2FKar9byBz7OxB+Xr3yK0KxdtIEQFNS8Vfi3GsTQNy7cs/yA
E/z91Z/TKzmdJkgP/oUP+OdMh/Ic5+HD52jtihcVFrjJ4OslhbWh3Q1LVofIfveAc3wZsbs5oYJq
vplq2BGigOE0omzKBn7Rjf8bbed6UPcURZ4lZp2a3pZPc472Mct60lsyYl/aQXFM8+czPKjhSH0x
YAay2aJrh6Bv1lsV+WE3NG4uguoNu6B94Umf+QXLH8EOpgiEFwqqBR6zQBuEOLwzqbixb1vurzSn
IxMOAffSRE4nj7piTF3TMW+gR3S3I0TB5nsHmAueUph1R0n8DwSSoG0YA+dN/aZ44stNz0ZUsQTv
9WrBaRSL+NonDmvRboFJxWUWCdXC27C+lnfLAod35pzG9O0A/ZHS5RyrIlFTJNO7zBuJA+UD1MDY
0/qf711JW8uDdqP4lWIdWTzANoY5DiaUfrJ7Lr2PfgOoaWZfBieyfhKLtI5Gslg6zRkRVdf5nil3
ONbUcIIQ1KLO+kvhRxZi7nmnzBRG+4kXP4cv2wszvPDjsKi6xKDOjWqr4D4K8PdvsP3a14w4FWTf
Ideg1E2SbGzQ6Bu9wHlYZIbrdR1OGQX7cpF3o1dL0xiT2itFWfb/aWfy6O7E+S7VKdUeDuBjXdbc
jpHIuWxMGeLOvcv9c47s8hdmWDFtHVzjeAdq4u5jAaSlhjjrXfk/mHDhDPBWymWqgu+gdKPShehn
ik/sRX2f3bXxWWm88Qj0LzYw2Hd9Gz72HedNQKEA0k/5r0UkjPm5YTCMzI98bmwRtJqB96QO+/6x
jaMxCZaK4luukK+AnQJP1ZoxwUiAUgf9cS1gQxNHjlILCf76tWP5GKsYDdi57A2euRF4fOiRT7sx
w+nRC8+dcngctBYUt7e9pPzZ5f5vnaahItB4BHTxgMClx2n3/F52kQ8CiM/JfgfvyebzYv42ItF5
Gz9yqG3suDhYgIHsIwntQus1zVqpnu42GiTJmBBDjTF0e+p/B4NGZT5gDcSdYSU4o6U05cL59R2l
omufDxqv555gxwib40H3iRwRo97KWgdWXr8LDX5/H7AO0AyWd6vE+hTfCUYofbFs6ep+EguuSYEe
rgxvqWlUzuiI96dU6X7sejC2k6L9DLXAZv4tl5VPZIaOm/N/ZMUaf0bkmjLU2wrD4TBM0YL0l/LP
rMe9cG9OxL2HlsOtHOZ2uBYbazgZbGI5zA/BZC/pFz1FFyjl+o4OAXhq6GT0b7vETHrY84/il56X
fqnRVIQHQKtKX9ED19he+1g/5joOgpdwW+PdLSrc8HIOQE44LdszvGdyN5t7r9HdSf64fn1EpUub
bLrYmzRzBJ3uGDBPdH80JC851SBpBrWoa3QJvUVVNotHwYzeYN3uCP24V24L0WgFrwQDHhEXTCGw
n56wqcyaWYFFldfPOPOpWyRpnxnY82+05Rywr8x+3MnhLqfmN1fydsBRp5PGAWOijFFg8/Lc2otX
aTH8Nlfrm8zM+eZXobcM9C5e5iC7Arb8+rtwGoCdAZRhKo4bHQ8shaJIQZTe/slIm93837E31/du
9D7Gk0gWgpMtPzmL5CTLLrx3a06ZthOxBLfL1iBwF7ayWvwUA+XIgpHIerbF43fXxocKIm1LbCAS
TFs+EJhYZ13OUlvPwAHNlFcVpbyp76aA7J3ApqHol4luCUe62XyR/PU0OQ2mkj6DD4K/hC0JFjah
cZQMADLG+d3Lh0wlSk9z1ONPkfS+7Oi4Cf8jKYF8wt9ZxquyIrJLTbbLt0CtTnmuyQ8kpc7dgbI+
Cw7YNgG9nshd412/p/akH/ox3Hsn8yJ4womx7yWoeRUDt2KFCCMXzkto/buY5Kiwl8oJdjnlsexC
GgxPfABOJVN6vX7FdSM9cflilfciBGuSgUegxC6R6r11mI1IC/exyDuxa/DgwN+Uvq8wMyY/1fI3
9t70oMKDCwpvlx8SKt2SSMWLmC+2rqUPvKriJ41VXEGbmoHiczJM1i4MY5l1hzrIhblGybkUM/R7
8+FdDPLbKlJgGjRqi8nnRM7EcwqpWjgcjzGhev8q159Fbyssg+QVaVB35qfIGlx9vr+1ZiRryq36
WJufKX4mo3mbmRHqNwIgtb5SoacoUqSY5LX9g+AZOK48A4NGxTIPuN09vYBWkQpHJoFA0zpVSKOQ
TfUy4ihxTYsejMa/3PzbsHLSGuJ1PmZpfaozWKRMg0dTo7CediaUR7CxoLaKKKv4SnoKnJKFA1A0
wfeVFhUsNv0oUSkUsp3Af6Fo6OtU7+uJsTQJeDO0NhkomnE6Bp0sxxR5hP3U0SBAmLrZKpe8r9cQ
29PPdkDnZuV3Eed8eziSOLQkK+VfL5x+WmsHFwLqcxfd5/103GPliWB5abxHzT1b35E/XhHumsvM
XhOfdSHBvekzhU3ABfe8O7SgGbiEIUZxX+ZMHN2tx/pQO+h95py9l+yC2NqHQdkRWmTQXK8R56Vs
OY4JMGd4+ZMUtPLoBgIRp6OazuoqnRHuk2nHvP8z19B7OFOYtY1kNylqkd6fvickDYBqNOx7HdOS
jKe+9hOlpS3sUr2UZfZvaL4JBnKGBIvlHahT6g6/o9/tAHwIIZFkO5O30Nh3CQ2xXq7jsCuWZXPq
hnxD3IDBZLAeAcYrZBLqCI4s3bIY4AY9DEOsbyrmUcd4gnPxRvMekiNpCJs2SYzRKsZhkdXqhI37
cPrmuoRkvSu/d/W6tqEUhJD4chpFZQpP35kv21rGdYBq080pGmi0HiMx5CIOpJZLFkSYepbqzIxt
3OhKwRKDO03zMHYIgC5brLzXCfWqEJnNLviEgHahVCVUGXT5ntouX7bPjsPH6pfgHm64mt37EFkd
tH5FZLYeNu2pjP/Z+Ot6TCaajC68LRXsJptpqKgiw6N9PI1LFJIwHHDMYv+j6EUfHgjFEq7b4Cr1
5L4FAw/ZBrh+JODPT2GmUs++5bqMW3JMd4JilHYo0Lr50iNTckjNyHdNPtlyZnS+mU7PUB/tHzvE
kwNSMlFuL1GHVs3xuliPS2M0DkWLFOWCRyYYLl5Xrb/roxcmf1KZ+7W48B0mzxLMFmpJ5cZPKUVx
MehQAf344gXOd0HOZ/ZsbW9PfeSTcwgmaazy695yhCrKElkxMaekTnrBC8iH8U3NDFf6/Nw8zNHk
eSR8IUc/KjIab/1bTNK4X9EHA4EcfpzZPy3U4xERB9oZ5ejtglDPGaYIRYMxFnXZUR8g5YftnG3z
qqfIPUN+ZkvKcURxYg0T7RG4LBKxj7Kb7AeEldUsCUkHomjuOoLNbF8yGEkw3F1zduhcc/gY7/dv
ukE5O+uM4FC96+BXeP8BQfdVSzKFcAPKsM7svzq1cc59VNCbmOo3xKzW8C2rqEbcJhYkic8AsYaq
kdObKOhnip1wu4bs7w7n72/IT1UPb65qrPh69lTHNbzLW36X2Df/HmGrzShWXp7N5ukZNasLCE4L
NgG79EKEL0x6iH/AEfsWnvr8fQOkBWPaLwx8NRUGbaubwFLlE7IRTnV+9AxEiDBF5BOe4uRJgzU3
7AJE7tvXbsLekbC0n3A6Rp+1bU/h7IJOsVYpnI1gNoNNpyB4pKh6TN3au+lCsdVUiebeCRm24kVX
kcH+EZO1QB7OLSe53hm98GZowSyAwcnaB8WwzE2wW/QVCUSvh8uqyQRdK4RRacu03tbWyEHE9khX
C6ez3hipI9onT2GZfj1UDajBp7E/0RihD9aXsqWxk1jGVBmiwFYpSMSg6VPtWSwBX3zxC8s79MnM
EGUZmoEmYbZZOCVoRRdZIQ9Abw4AmJ12qJnIFThr+Yz1PQwkYCWO7dPS4061QPfhx6SyQNNVPYcG
jc5//7sygUvqjM24hWle80GrABc9GrFC8CC7FjOLiiCWtiVRKR+h09yjyxq5Mk6h0gRI7MQwLopd
EYV+iHcy8+ae6lKgObp1ScNsusUGd9GXbprcVvFm5b2x6XWK01F3aBBIq1k9Vk6z0VOQU9pcs6LH
b28wLGCSjeIXc98PoK2LIowp1gew10Wl2AeFd5StL2LvNmDcikxtOHTeiU8vuJNG2eYCA9A62Kji
ujsDwBXBe4a/QNsxfVhxbkg88CDyfR8ihuluiZOeDQk180S11d4Qg7gJQlhtSbVeNnM3+Af4gXXA
akGcSeL+7EngLoC8DHngHHPislxqoN8tzStps//gmoMNmsXQN6DZ55kuTDS8wtGp2sQB9rXv7Gkv
v5PS7t4J/tVpgkQO+RTyJ89+F6/Rph/n9JgydaKnNHd2PvbwUZ0iJJSHmEoN0ifWeRlp1S3GQQAJ
aV63surgxG20J3m+VRWx2KynBIgVNRlSV5WwaUadyEzJianYfHk2O0CB/165z7DJYtsSO+YkzCdh
CwMxR1aeJb6Syw5FhB4Ix45G3TFGhOQrxSIrLn3ZU/0Ja+PJvER9SmRYKGZu8gj2FiaS9ssjrRIZ
mKAfRKMjPLCZFa3rXv6MeLO4MTwQLqv4DT4tuaPQa0uI4zdnmqy+BqytwRIJdeR8Spyceyo8VZQD
CqYy3RwM4NYiogXIt++e5lOBfgrNgk8lA5HEFsdMEFUdCIWtRSCjI1P2Z0vsXrv6TZJBLcZMnklX
F1TxTrkShXZZmxZ+0FF1+2Hdvoc4z17VWTWxptBm7KVyhZYqqSJYtYkhDazh9SlcpsPJ1HZBhs6O
maMwfagZXHX59ZS//i23Uw2MMR1Op9iq38gKzTBsR01Gmy1vrJgVQCXJIdEaP76nUcoTmyCBRbtZ
omfAEBHh+YpA/Vm4D8PTCh4IMMEo9dmxOh8EZyN6v5BBa6FxUZUXJwiRH0o8vAvI8hKYx0I1q3qn
ric2UXLhdDit6CJWzktvOGJGBhjsiGB4eEqGVsuTBB7xrt3hFS/ktYnq8OZQSxF7TG7SP/szrUXp
M0kZ7hj8QNqtrx/P5627FHHHGXlTV7H93Bq5KzIfGOZDiLNHX0ioLsoUMcLVUT0GSii7D/lWnMoZ
HyEbir/HBa4SbyXB29VylprLMe/pK0mbMWRD1abHbkywAV3psQPfvd9KVk7tPwG3ERnKshqCuJMw
bLvaQYPFv8EfZ3qTlvlnh/gMBmM9mRDKC5bSzi7G4H+zsDDtDIqbkbiTqghw/SmKxGRhmbUt1Kfi
wn5US7V8YOjzefGRKTgceLsJf5Dv6L54F/0fKkeuYn9uYpPXWsl0HnEClM1Kw4qERcw8ufoC6ZNA
/GscNMHz/EAzKOuSZvMVIza7Vbzmx1arXDKcT2xHbzxaVters40Hbv5lTNldfzjCFWabjR/XJlkJ
H1RlIhmQDA/eysTawXK7nnGmCOe420FtHF4TTGj1qOzDM68GBitUUxRfk9hxNEYhqRvYNf6us068
vnbmivaPtFdQPgTvoJ5HcwINJGEqIGsr1M5ZwAKRLrqqsXSY7vjDGKnWrjZSd1hEVfqfHtKKIMsU
egB3Gf/rzAIbSv9vACgSoSTzx5NFd6lCi+BLg5iaSEPQuXZERClFOgalcVjqDnu1NpCub7GqUyyV
/9cgtizEKdklluZlWIHlKYsY147UZm1tJUD+rWkiikBvcb49x3mOuTDcHau1y9FYBaiEgoNIhK/a
vqCwZEaOTS1iTaaREZ8tbqqHdGYsZaxVscKxtNc7QwQDjsjgI33tyZPcnNZAdwRmpSx2HG/egtwq
cD1auyRGkZqeysScC0+HPNldEIPLcXO4u30Cdafre2IljrEgbPDpfhWm2v6lxWmLORC/JNzDVOh0
FezUg9mJ7FvBvOcqPSb8MJoiw5io7luMBN1OoPSHMSwHeNzTH6DgOpjSlQZ98atUq6c3Y0Hp4p1Y
0dqmRb2auI4peHLM3N97yMwEw+DYrx75NRmjuIfGVxhreoriAoho0aPFQWBfkLhKxgPGlCdxst98
RaUPTiERaeT28bMrYfWWzTIA1ehJDx6bWx5x1rCSX2gO0V/Goaqi1awbaDC1UNYkNt0tDV64HAos
SSKybHP219Dk6XCN1OB4MW9HB9NaLt7kXEBhvmgjymWMW3XoqlJKy+0PLlAx+Wk94XItmNwZURnH
BM1/mGaRAWV3lVL8Q7nvmppgHVLni7oX+QMwVbFEyu9mXkDCCHh7Zy/zYCGksb8mBUlxrwJ1PTeR
0p0KdgmRHg6F/nXOm2Bn4fyNN0YJv+W4D+/bo9pMuTpdID732RZ3fjmCWRsqeP60I1YeRrtbR0rA
mrBsKWtaf8lSUfBWJaPt/QrQ8koZaHx3/EUEPT66QAbfhztOGBTIEs9oyNx/X8y1OfUhnFnyUund
9f1inkIWeRliRYIcpP2dF4c17z+NKUAtFGk8tZkhXtZjrzb+TKgbeAXq9OzRvkhoRpI19MBCc5Hu
pa0JbieZLuA4frrg+JcvlGXMuDZAYnRlA7ilCPijkLqk292agS71Tdj95MYUgC48vJLQGo9VNC0V
dY9Uke7CXExddCqwvVNArKTTUZaYUAxS0xLc/kSUcp4FGLwgI3Udn/0/eF++HM4QPmxYvgWe/1Um
ndW+zDW4rv+5m0av3F3bUIIwmG+JAECw0isr1X9OftSOhN4M9fvaCB12oedc5rpo1/gH17Pk0mxB
MxgR+Ge5xTOT6XyAoz4CUYAEeHaiOr8xd2DRRRM47TbGu2rNRotye4JOeNHK9CQVEs2sIK3Xk/h5
qWahN1KjoSxvJEW9okdwTwvXWbUe8UeFfXsycDE1Ysdd9/NYF47BFbosLd3VdAwHTtafr7T10Df/
B8wj4C2ElwUXxb+yMsZPaWhoBeVJcA4YycwhION/UV2rz7KbleoubMluXh/SfFrxAItYDk8y2bzc
L9t9Zs+Zk9YKWaunkXPZUe/cc1aQBWpb9ei0JYCp8C36m9gbove6iYUdq1iCY0JoWVfx31YMMR8c
y1UaWpn1KbeBaHTzwQhW3X3ShbLHRhU/zF5VGB3gUV9Q28zmZCpMbAVBu9ejcjyABZYApPLjUG2c
sB+zbMXsicK2pWpaheX4MzXs/Qa56llE8Tlb4oSs21VqBoCA9PS2ABZIJdbBV3+UWACl0mY5W5HN
04MrqvX54e6ZDvRrIyIwGCEIKHdmfFpG5pqytHZPF5oJg0YA2S3bCINcx9NEAWGihDBLcJIT/04y
KvQkevSMhfWEpKNh0sCm/NmdiRUE19rA9ZQ3Dox1XcyMTWwg89KSaqqvO6fh4GofyG9h8+7nszNk
DtwH6t7ziBCcn7hCtCwlv8nxwp+2LZNTq0DF5lyym+G69VVnGkTJawaoMLoA9t8Wa9siXuW0E634
rd6Jtuk0X5bWJll0jAHNP5UCyd4Tq9H3YluqggWk4j9KoC2d3M7FiX3Fl/Y7ExvoRlQ2phay5FPN
8YhWzZmIpAGIi6lswqShxFhZIFiCtUiD+NIDqxOD5XpetOoBbjtAn4rAtXloyN1uFr7qV49dTbWP
ucljj87u53bNV28mqiVhsYy2TIi+FBtQI61qWVRrWGDNFgmh/+C5pq6j+eGIGrb9UdP109NQlyFA
lR6cRxRMVbaC0RLyNhGkvJMpBlMP3Xjzk/igahh23f6XHtj2o9Yd5HPsiawSVDdjetRrBJ5+wxOC
Y9UXZwXWoyuCXAgcF3ubynzfWmVQZ/LZrjQafOHvTeXiziyOCOKq/Ibf1XNgVDwtim/OLJBpKZ3N
OXNG4kgXWjpKiuErWxQHgA/LYKwWHaQqWniEgxW5OvWGIagVGfH8snT93LOHPPcq4hDOrBanTqDU
C68dLK7qO9S8L1L/gax+Fuf6DMjQ/qRrHNq0UcdigDxg2ptmLwX66nSfzRw4+TmWhzvNJZbFxyj3
q2HaS065fwAznNb1a480Qvw0K0AmfjbD4FsJSlIIFDCuVmlPXH9/3974NGhpkt3gT5CWVjgdKP+n
n03n5dK02eckpDmDZeEeCbbhCmxPKRNXMwhNXNS8acrLWtczCFkfAR/yBS28Jz6md4zQS529i1dc
d7bPb+605fL47k7uVlTbKF+/8gJXMq/s5NQ4yK3jlWXe3OHoPWRFJSSWonik4iD61WXe8HwVnlgN
rc6RWryio8JljjSwiYDosnGBUaxjI+OI4XsaZc8wUdBCdtgulLdZ6knpAxKsh5ZuKeMmEPeh9GN4
7MdigrixojrHFAKNMNu0ciXZ+c/P6JfAWgYSt726RyEKx6PDWoySAdgWpdmgfYI0sfFx9YVaqkP6
/HwLgYqlcbvjchwOnNeRif9DkofeHpZlnwjr1CGu6+CLdWTROZ7wxkwHFyoA6hFN5EV9eZRoq8RI
+qtwo8J/Lh7Dgxa4U3718dzBN0Wvybc0+WKr27WEhPFS08qJ6UvUCx2iibwZwRhkoD/SZQdNotw+
fg4bcAmwC+m/sicqCUQi7v+/rp3IeF8weenf0EWSqxWR5ku24OseZd6fwlt6cRYnAQ69lzSvjEEP
1BeBno5jcyCOrJvKwy4EITAFUbTTxkRK4h7yRNyegJ+IveAIsT53wKe3Pt8OFtBYsiMIfa6tAUtd
JTycJgdeCyuKHgbVGouEW3Z7UmsvuTd8ekpPEYC1+/1RWYvIA0ODq1AekSoO0adTbsdWXmf/K08Q
FY/0d81PDTaXeh3Jy0ZahS/fCaS9PwhRSA9ugBBl6sC3CBlepkWmlGqGyudMaaVQmQ80WFnxcqWv
40sYGmY5nnowf8o+vmw70WFaG4GB7PVT6oyybBlGqo1p+FVBUa8oLrvWSdW0B0gv+oMsuxfX0Mfn
uoeIDsU0sqATY63O3Wx3/unOTnilwQw84/HCzXfMUIvr8CfCe1eX4KQL3R/GGGEIScbH4UcRxety
anxF4LOQBFfooyMwd6DvXPe10nqx45d18fg/svttNVYUe6kBbG2zC7fAqr4bkRvjdRY9OVHBuvyh
gPXezHxTd7BME+uyuWl3MfqnIrMqWjhR2pClpgc2SSW4rqEoTtzdU7+oWyygcoPk4ZoWinahyGcv
72FHQUiZU7OkQ89Crs5ZcrevPLFm5ABcY2lhfRu0EBHtDp9Nam7bOFatZtK3YqHYbSn7GQdIWpCD
WUAuyI6B451Rt4Ye9sJ3yDwK7+cWREgjw7YjLLkmGvXbmy4zyxMreKqqpX5Ij7+kj2zPvQIpYQ9o
127M8TSezrBgPSRkU0N7PR1HNLMsWhJS6OjmZSfwApv7cp6jOOVfihkusXz3kwzSudW1zDkYcS8z
stJ1of8cPZjnwKkG/3SArGneIXLG7gaQnFGAmAExOxuJgexhqv2ewa3sn7zUcNgfbRXDhKyE2fny
GB6PSWI2WnoNe2BX1TqNypA7TD8EUgzHlRJsRX82tqn4BidViazGv1XiKcEaUoAZRHR0HdPF5Ryw
sJLBIDSKq8jwHFenN7AshgE51unZmE0JnQK4i0mjjaYlN7YtvBzGWo/fgD4T92vZ1KONEmlv2x01
dhXIV85VK8XPuph+GEMBh8tI7EHRVD+48DuFp7xj+K5M84UQSDFJz2ZfCKd87T6n44nGGn9vzdp3
+1R6iQ4RA6NRi3bzV0q9FlyQUja64d8N5GKhJSPsEFI+NHi0DvEb5mo0QpcfzICRJi6D8jSHNvlV
ADaLzVPDcEGp5g97tj5ASD9wR2d056p2P6y+jgZynqJCkvo5Su1RvVjZUhfAqfYcghq8XXO2zooD
Vqbd61K6rNXUa+uqoOl9ObaaU4rEw8FvkvbhcbPu0My7lbh0ef3zTqv5309NwMnSm9RiVtkMcoqt
sAOYrerUOdh4vxBIaYGQyUXnrEZ/+yfHmlNoifqAIfKqSKS7tXHPfxWdvmf9e3Jgwx6wUPLKX7y7
k4p0TmJBofdxZXItX3auMS30nDMmOmgrpsg0KiMsWz7ixD3BFtE0S1NSsK09Q9tLzs3Q6FM+YNw+
x91AoNFjfEWRJ+kVJBpKl5WgdEuwBNMYCCBtrIh8TvzsvI72xAjZpyrN8vvqSZA6Ltbgq8nWczZJ
M/R2zxAHiSyj4Ffamk4ytBo+LDkZnHQUtB0EYu2lG4JsGo5M3udi8wSdJVYkayJREccKDmImzXio
2CJRTFVhdHo/wZEAhzcYJr5Ark02oCHI8WnirrY/lCcgl2bufoMdQ2CjRQDcFR1CzqptqE3Rlm6c
q+DBK0I1Dy/m4WiliuWtOlNBzn3JS1Huvz9aXZ8yVPEk4bIx9194m/Alft16WfZufEbi76ioEX45
ZDNf9YAPAHN61w/ZsBd72fLOfZLzWKdmxksxqdNWbxj0SxXPh2L+L9qUgy6Q7boCzRQQNilCWT0x
EeypDDo/3unI88hqzcJSFUYg46/qbyHCgkFdkwUUDiLb0+yOa9z5zfZKYMJVOrn9dne+jyPFfDwu
GFFvKJHCddezSfNHSIOkT4dzWHwPp7JwVqUe3wkds+E1spzeZbVYRYRAXigqjCca9vOW3dLZysPy
6youIOeAJ2HXBuViI9yuqXhVBEnH9hPsMvmXBWEwyOkjNiFR9SiVAw3Xm3fZvlpCKiyALuk646ih
U2Y3pRlhIn8p5HerqeDbzMEOuc8cIKSfUnD4JcdipOwSXwzy9zhuSgSKU4y3gOC+SLTmEKe+XfNj
zcxPceYUx0HktmOFTrQ7mbWe1DSyn2YTQ7y4GpFwOoGHcFWecsAbWKuZTBwx1le3nCpxd5p7AZuE
WQwgkuvCbLQBefV9t8VSwAEKOcbSgMCAXlmuadrTGMRaXXxkIdIQFEwptXjJC3rC375JHQAbbf8/
GHu4S9t8MO6Tzy3pcm/I1g9B0jPVuo08jU0L0V5axOJAyHAuy7SjhaV7xIor2X1aKQrcQPYXJY/v
4ystSShrXBigCklpQN/nAqno2ZCJalCRi4Szkj4SxmZpXj7UbOG+XoigjGPZzpBuSeHZtZy25ye9
oYlFzQnTt88P9i7DlqVbiLXB7jElOlb7BXydo4galaPgnalbwIPJOAIbHQAb1BfzBtfHTwnPqhbQ
bZQCB7ylGJxLDLXGnwhGiNxwoGdxr6Jz/lThhXsf1uulobZwQBZI4LsHkcWYUsubUJ93mW52Ofe1
S7xp2hV+Y3e+GuS4VO3jWJ+0k3GAwT2Fwgjji8Creg4F1Mc9kvjlMmm9gFs/0/T8305Ex6UwfJB8
FIPy2DFugXyLDgetXYInsYWP3wPHIRm7TdrP1kym9u9BVWL/lg1nhpMjFPZbzDmm6lLTztPAwURW
NDvhrxMCy4x8wnNR5NIjCYGSCqxSLJijwhjURhRahpwlazEx71goSBnpidPj1/RUQQhVgKm3jmfR
T5+ZS6PW4+C9tHTG2FG/3lUMDo8Ok5/eLma8RHX8hlB4WR5dn4ckyDmgKRULasscKFadW/Z0d1oj
dnmLGdbGaW2ra1o55grryDg3Yu+L1ilwIkW6slSR6oGkHzZHxPoeXkGPo/gmIYgXI10AUX6azYvD
OvK/gdraxQiZnb95t69b23qaMB6pW9Hh45AVoKkmL2glw/t5xdiZVdts6CImv064QogEhbOY6Oij
R7QXZLW3Ka14mTq3MwD52xBKZsJVgB1Ge19rG/UV2ndffuFMuDjUWEw6H6YBDKboONOdKjsYZErN
yZicNF8y0rIfgZLUY0ovj/UIdIqSzPzV7n2ucQ9LYxCNymi5AhfPm5ycq9exQTb7E4M8uq+D0//i
1pcf7/fDMSa+JbEQUFKFPNicdKH58kFQyTpUCkoKek3Shte0epWiVeNLjO/MrPnqXs57UreExWt/
Aw2gU53GM2nlrVIpiFCOS/Y530H8mh69pye94ClaAmcDACehaf3M4oY5LgrVwJM/VpMKUpXPK9vZ
FOMOGb+4ifhSUVDVYLLpdLYVd5htbuBpu3QETjC7fw3EKiDDYl+Nv42/eUB/OzZmZfTAeJu/03+I
sfW5cEdxGaMN4UqWOfXy1h7AXP1TrVyk/j/tFJDQNm4MTYPM71B4ANvpuFD6RAVfZlZ/uePpQ8td
yHgNKHiDhs1JVXZsUNYieLeQ1IjexichRDTSIjKHj22JR2rBJP7x7AWvc8LkK4TVgSgrNi31z8n2
fZNtoBHvNCY8KZvIXwNV+xb6+JU962WpXhSXfBlc3RemSNy6+aGHRWOmPqrqRzIpXqo9Ha9pZHc1
teIrDbK0H17epAAFoW9icC/MI3j0bi2DDc60b3ctRIqaDgwSnLmWXFp9Vsi7NLuNccRpawNYY5Mq
Q0QmHnJGZniTWZcbrPEl+Mr1guYpBVK1BTbNIPLGZhmXfP1bE0ShczcXCCnSYEl9iv7RkaMCOil6
tDrSVbc44PJdkLGXAH0/Kv29JOVCHetEwoYoPJKOWRw3f0XZzKRmCdb4Q9Q9Yj/h/lPAG7nB3Byo
uJLHIZitmGnRUvH3tY9mYdCjMaAq2GmBlI+xpjcVLEeOrdSOCW1qU/SaZws0IAamw964iq4P4Rkz
ddgEuH9c7YUXFYEdTcVTfgJgFnEQdzw/bTwh1GLMvmWex1x5fXFcgVYvgQ97Vu5Zd1K95qGoo4Dw
RxRhSKtaWP+eC8RQ+pQnPo5JTBjjrl1gV0LCKOkysC0T+jzz7gRtynhCmZPcuzRvZqiI7oA0ufV1
njZ9/NWNI1uwFEIvuenjJfH31ThJoFjFRtLL3Ewo2TbgiPj0QrKACt0jJkWL7Jct0DEBwViNS3Zs
bg3k2Gdds6nHBivPJGaH5ubr05eLJ5+dQ5rOxBWzjGsRxlmqOrApIJMauxSNUCU6xup3nr4Vr/Go
il/Pjg4PH1PwsnmPQUz8ghpFq5F/g3UqBeS+Eo8FoESF08zDU8Pl88w4brH/Mjbxg9fLPWaceGP6
ox7Wse1zMEl/hV05yaJaJad3mJbGm5V3gpCH61xsysFUk+X5BDtnpaSjBk9DWDTDBwioNFIpZVrj
ebynpN5I/I6t+bo94AHFsmCSrA6xQCnz1GsMLVs34sqfQHBJaeW8uL9ao4MTtME7B4FrCRvQ7Ubl
9H+Pp5akv/nidrbxucQDqIx/trCjYJg9AH5tk6BNhDmziLFqrn1m8Ht8EcXACXlxk37QOFgz00HK
UrbcUGt3IiPK3Hr++PcmlJ7KKf+41Oz9HH/h1BsdArxURSqgaqY0gGCRY953f2UoiTTpMUS84FlS
rWhSUJOUCzzwYAFVkXaWyzcjhb+cOM96M36pvERcaZEm6ngVdB2RcDeS2+YE/2wulQpJfODyCP6W
YqWm062Ju1ypCLwVEvGchLuGP6Uv7vEmasE2XxHazSp5eSGuHR6c7+5D9dPeiT6eLtUHGKNy0kUR
lG+dIEBnFjlVUUJWjnWcVQgMxzuKHMcQ3qu1fx1ONQmk4NIonUIz30FO3aJvvUfJPx7WPwvHoVf4
bjS5076YPSDEKNKjFVSk9U9ZVgkAw+t5I8pkVZ8l73jbSOYY6PWe/e7UhJp5nM/ZMLFN7SwWPgRe
ZBlr425htw4ZFvGoyTEQGEoCmRix/FdLHAqmaw4qEj7MzJTlGWsbULH6ycsHdkkFROT0Wc5Hkh2E
i9Y2fOelb6Vj9AUHcs95QTQ8JxaBy6E64wQit5aLYnKehRj1AEPIDbcbOXQHR/XjcLgXMkBKil9r
FtSsvnpbaEMVtryg9KbYtTk5BUlFt9lfDPRWuPy3qLXFYnt4KbMk0gKRTiT8vxynBS4wAB+3EqA1
NQMFanlKmQDHVvzFoPvri05jd1eFy0nr9I1ls1Eh3RRvOl8kpusUoQPpSHHTrn5uF1QP2VUkeg+v
QMhQPCl8wr6iFMPqlhW4nngWxu/WSM2ozR2fCJgz2lb+l4lNFKsA+4nak0ozPSd0aeH/jcJUSt+m
XCZ8HkuLVpAWMpASxnyDPK+U1v00SzUMy/w67kUa4v9zAZ9tFaxxpr+8KsBbDp1Gjx2A/wDIk1gA
2+TdYCT+PlV7v/Gg917UkWLDE1hzB08psXCPpcqYUMvC2PSv6MLDwglnxYpa3RZDv11pRgyxjBZF
MEyG8MC5nGraIfi3cRnyKsW3a2VT80ltDe4aAykCo3aw+aRDaToXMZsZwT1qpht/9HtgMrdty1IW
gbgxXQXbpmcZ2svv2vhj6Kq+WtsWlGZznHO+JFK4WbE0Ek9oMwcsA1tZLqg25InMvLAKTO8XPzvS
fH1h6OYP6HdAFSKb5KlNPhpscFwqtEVz05O6fTuxmhSz0ZAJUxsedp167G68jJPulqI+w/IoK98P
Sqi9Y0uW3Eey1pZW2q/MA1whfdc1fe1cwUMMtvoQ1B0chvHOcQd1gooA5q6CDfCiSzVVy75hACD7
KzfB2Smqhe25+0LNoXqaGkvAmfeLHkSogltiHYF5ZZFAhFpTCGeg6iM8qra2b84L4YwOHfFTC0UL
72YCf7M21O8DctpMWOl/SOg7Jvi84f4QxyO+qMd7affGKwbDmTigENr1t4n7iNz3kSawHa9/w8jQ
Ckc3S0jgAIzgdgJdKjBS5oIF17LJQmO6QJXdQluZsAsBsJfwUkQ7ZZa6ndxDHs/O70ZdktjZHbRC
HgBNVERWAeTH34XGXRz0+Zk7EDroC4z005hgYyTflUyIpqxx4/kZHuIVFX6Xjr94Rr8h3t6+MUGy
lJFaYfZWBPDVqtgK+Ed9fcW2n2jKWLkiKTsh9XBoXfkU2XHK86/KkF7u5gSxM2mgiKmuy6ebNhSb
xO1aUhqGlBy5j548kB5i6UPLG2j2/8JfRLOgLqZmnV5kv6a5kD33GKyHD93oEptL2svFI7IECJO4
c9koRxjToCb5qOEUx9k17oFwGh0V5JiigZBdXeYPszq93kKwWDX3e5H4FpfwG/4YTl/oWpC18qFl
WS8CZjlti2x/m6c663h89DQg/cynuthDZLXUHTOl8BOoABRTmIYHywX/pu1RtEq094npI1WXZeFR
1/Li8lP7p01uXK4xPwMXbkMh1+yiknKpS1dAGeyon89vCMmgi3jMBxbia0UOJ7RhBHLeX/mqLTr5
h7iGzelYawjpKuobz4O0Qct50fe3X1pmE6NS9XDkSM/QHMqz7Ar1biDvCqqOQgimGGSv4ELNbvHt
jfK2X9DKzyqOmpM/VT7AV+Ioqb9YubqCK43FYvmPTvNvOSzzvgWHiNlmIFwSI8pJySkbicxVGxZq
pcDXqQPGWJOfHUCEUZ0r4owR0ZyBRsAe8CiA1tqz4EBgqVdXV5uKLezdncvXP5VdwUQyvJc+WlGz
87d+7K0Iqai46TLUVdPDOu9eHPGg/4VvkIipAZ77ExUlerhY+0o9J/5egQsnkjkN9Eb2VAF7eip3
oYEP4miw4GZjuZtNy0TRJTAnNZ96EoyJ6dWBls/TxVlKzub7Kf13Ash39rbWVb4r958ZmWMSUsLJ
fHriBZB2tXMsBoE8EW+ohcxd8UjUJqtxrDwATSDfSBc0aeeF1mBQiXjQ0h0KJAtb1JucVsO3zeE2
qnLcdIyPC1iuTEbcaoCwq2mvvietUSRtWr0FzXzK1yOWd+y+KbuG8w6tqOsPH04rJP+90BW5tX2K
Za2bOMEAW+o9yNhMixaXUOY9/EzyHobzIjvqkqGRXmuY2wFclaxBlbmgxFVIS6PxNxEXo3twEcd0
gq/BbvaHDmEIMMKLVN/e0vXx844n0Ns+f8jozuWdan3qN40Y7mI1y4ICANzM6CTPKlXQVYAgj0M1
JhK7K69l5mGXIsTNxf4s5PG61y9YwNP2fwaINwwMvg1Fzka2aPncph1Jr5MmfcGe8XDEJCwghPfX
VpB3XvjtjsD1foXpsZziB2SnX1eQ+IEbHCZZCIN+FBsSPVacpZKXSGvXvMJvexfHJ7ejlzP/DXf1
QTPpNWFvsUsCjpWl9siinN0tvqBC33Fc93YF2kZT0bZqEv9Yu08QDrCmOz4+YrAubzZDjGWKokIW
BXFL00jn/5O2uqT93PGjrwiVow36IKtGJtrUJwzRtZ24y9GFgboq29D/U7WNqOmSomGB8Ub8XVqX
+BfHUEgKXCqvgPKpivOCrSlnC+J5m0yWc6dJUCRqw/4nrzUtEeaiRPbqHzjK1yNkTo03teHQjNrk
zYUrhyUmrztIjoyiqBCFQjT/gdvLdMIa1cGoSx0+mVtuX43xaTQmH9OmWHRpg6S4CMt/jYtkDBoQ
XFdrCe/WYhx8FXfgf0mJ25bA85DFNiu5e4BMn3o/UXtOo08e5ie3keJB5pAd3l3Z2Wz/yyEQy5no
WMpGqTRrCf6WUVnmX1r7YwpMkfv7EwHxq8EdTecYcSPQ7V2T54W4dAmuCT1bAjKBV6LgvmWYVHeE
NeILPmCNq2ZtcGgr8Pat+7E9h0xJaAYOqt6s2CM1qLMkwR5smRUNu/UTVoQOTSRwOrz4Dm1kvArG
08Zx9ebYU4aqmKIQ9oknfnxNTKGAO0s59ac8vQVNU7Fi0P0XFvZAstekT9yXYP3ADujnBnfaXup6
b2DXy47LRp8ICgfmmZDPL8pxDMbqFGZBq7eoe69OuIEhD5N0wtSJlSZVIvg9iaakRLI95fIBoIma
l9garWP8oOrCmLccF4YTSIee2naASJtRYyXH0RcWDNPka7NY0iveyKLZavMHXX+eFNLorsM42ff0
T2CcyAU3C3Gfn5OBIHjObemgraSrch+GSWcnwDEc8yykuzeA95ecSIXHuQiqikHShikk8uVQjY0i
Z5RPMrlqPZOZnWsW9a9aXTYVUHG2WjRmaR+md8aBrXeo4LPF9VwgLqdl+cAL6SOzIHwyLTcUSf1b
lFHtq9bMlie6ESuU8uszXQaPIdU+apPt0PKS1AcuyLvCiNpcDWUIqDoeMYmoPCyiogs+RozciMKx
SOr8HaT4H/Evr7OWnCDyU0jtmDSW3AjdGP61JcPQf2pv8j5yt8yYmmHssj1mOOKqz+H1SErDCyRZ
AoDuO7DxZTq8uGwqJOwDbBiJVH1b5mmxXSZidsN/ZZYyiiJxGe72fkLOipTdUISgPfzfAlTw9UFU
W7cV6QC1mPw/9qtFybdfk2SABOjz6Bsx6CjsyCTbwZUqC+dk8d3h6UmhDpZJEtMNkLt1l/1eE7I0
MLSkk2GS+TW7FROOnJtRo7aH+ZYYUja2gO0e/YPYJ/JkVpjDwXELPPijLDuL8IJbSHM/dR/lcPgH
h8rqGyAUQZGK4NLvDywGKRlk+Qmt0sT1hh8wbZlMwvXgIm4JbSfdg63LsbAUsczt8erY0MSVY1ah
XFTs5QA/RDa0UtIf/CQcw3t6No/qKklw9R6LJiBVI0kpcY4JQvXdiCcbuVVZIr/WIZyWBayldgXo
AG2QgYkVmbCTDe5T+ugtOp1/oPnbcQQrNDE30S3eFoS9xoV+P8cZHKY4NB9/kp8AP3efm6BPsMV9
Wj8ED4SYdGGKojPKD9DG1KVRX2eHGm8htSaJttSFpxsQO93oywMYvSsrsondrVfpemW0rYu4c9Le
G9luo1WRby49xZlAupYHp8fTEZXdJFI/qppdUqXWvMIiohXswkU8y0j835bsTXhJo9bRSr+kLqd+
9CNDk7UGq0RR4YcQN3xBkTKPspYegUm98MFOIrY7l+DcwkqBMtrSY1Z6hdR1AwlK41/cKcxhDaiE
JfB3V+E4/3LJbasq1yMHVRMosUC0w9Y1q5wtIdjyAEX7yAUpgKTPlg1Sit6o4PMPjAz1gfWbe7HU
vYRWyb3dZ/+y21V9K4Bl25nQaeR/VYpRJy2j7Hn3ThBcQd3R6gGTRYqWL5IfeCeEAM9Uc0GILu1M
Rxwa2RZw+if/ZqY8G6GAHK9OFVo5avVZ8tFyTy/f1nyFNnoxw0DTy7eOlEbXA2xSgnI2G+jD2/xN
Z7dyI4itccCte6DGU+TlGLMgdThKesLq5vkZ51it1xTvXlzS6Z+URGtDpWs2QKtGDTcad8yIn2Lo
n9X4YiOcbQieLFcOp+5V/iwTEmb4NK/9xJlsB3ev+FzHgkg4TXJPTgMn36Q+WBNSVMB6yFlrTCU1
HexjMlbdvZbtEI3WY2De1A2kVj5PHIADyNEo0eXkws1b2oNZcudzKRO7BsSZ1klNuEblQyH9MX0P
7ga067sapcmRMq7k6DKpJvKoo51Itg0xTqvRHPYUK2OMCbv41BRZykgp/3vOu2hp8wt8wnIoje4N
3WSGE1XHeqr2uMISP19E67cV5iYo6jBlD+Y+8PYLIrkCI7i8bEHVployZhiDdtInVrwPcwOi2WKX
PEJ4p0c8H7rjeWcfS+BHcDaAolFtqRvij4yRPd4VsyIle7kJmNrPC4g2Su/ZWNvTenU4FlVJ9kdY
T3/mKNHAKLB+eEWW/xEQa5nMqtFejRLnRVbrM2isw4cL9jmLJSWIJMzuPoLmUG2pBH+krv/mkJ+9
eJw2DeOK6ponNk7HZvfoTaYtju6IngbnwxFWv0JAnrWHI8x2GCBtINAV3FKXInTHK8L4FgGMsJjf
R782yjLncBCFEbJOJ9jsoH1F8vcnYgP8jzBGgQtyZm3WNAuyG/ToA+UeWo750D4FNISTeaN/eBJR
FiR5ZZdp7ysDbuhTLPLB8qS1k4YKDZBg5LtqZofzhd195yqY7p8lCGCIgkFKutogKQNaimMoeOlG
7jX+6mB1wTwsG2njqfSpgNnF3KE5PwwlMi9KiE8AfQLcOkIV05npKwrVBQHSZpQoLsvf9BBbV3gx
tcMzZegrbbhBB4H2xzVGSereXKjO4uitzjxPeMrU0jU/ZI6buUSNeRrZpXJ5AgfNwZcEWRLf28Dj
8IGrA3UrszeGurhbK33qxVB9FUTPfUTci66PEplPKwVsPQPSQ7bTRBCIHwjyzXFgqZ3paSl+teRt
VJosEC0QT4qdZ+Jx+dp9vzqA0i1gqoZy5x0MB+HHWsJHnUk2P4kCghXTLGrxroIx2u9J5IYhAAjv
TlfQw/m79Y2ZJ1a+B9+iUuz0SaTwoqWK1z/TGZv6HDt1Q0zZzJSZ4rSvllu0ev6v4gsgAClYkXLq
/C+OrHbeqkKZGoJIsL8jOsTX0qJ9NhjVWAk4R/vrh/4xEwbQaL8PEenn1ocnMAarUTFE2B5hvgMD
eSsnHNsE6W+G7OMAy7ohiqukH8i1ZzOCL/omk3WUs41AA7BERRKKjAky9Jz0bfSAxRGrrSg0qFe6
F06Q/FwSQDaww8nfztN08Y//e/cdU9HtEDnPfNJ+emE1yg8WNCQe/Hdf0BUza7PFKJM2zUC054dP
McktsWrF1XEFnKacUOea0/HFuUGww4nJ1qC55sPCo6vX0wQ7IlpIJg0SAJihspydY+TKZeInM+oW
pevPrtcQ05/5LwJ5gPNvLDHfBZ+FLa/usr2s3sCLpVBgKnAXiFbMDS3/0nk/XeGRS5QSmOKDxPTc
rFQPhnoFjBgbfUW07aIU2q/dssnk3jaIJeO/yU4C9jxqIIac55c10h46fRtMkSO/v4yqPG8u+6Ol
hDyhguqclxlO0Rr/pB2yzu8q5ep1pU/bz0n7K8n4R9x4oqCBdLNS15OBdphGkCqMptoCVqxSCw2l
HWAsFKqZ001ba61tIS3Md7eN3HukFKvKVYgKQ5M++F78oVtWAv/kHNsENNVkkByNlL6fTu4XufeD
7NjZQs/FXFLxg83kJ6GAeP5EYcey1NiwhqBLJSNY/bqXj6iXOLnkRAELg3Z1VQbV6l5iCHyrNFbi
PU88WSvK3WsK9WuUmjvJ0LNCe4Kv+BzkBYY+w0G8s3koTuHPoJ2d+NvPzHMWm5MvzT+BqJ1EOdqU
jJrd39U9HguWv7ZwRdQYBm1v7j9+Y3hcUwOvsNJt3QqobYw34aJZimN9es+RvFxxGvTFKd5sGwhA
BMuvhTrnZ63Vklo9wWdi8C99jRG8Jm8w4y6PY5aE7ZzrbX8o6mJspl0kLQHJ8Fe0msrqAwGpIkNm
XmhiF5wwM3slvCY73NY92A/yJBk02V2LcZyy2XMJdh77BSSpagdaitWOtlHO7hmpjRoevyUkBnKu
GcdU/UGzhCS/Q/k5xBhUzQcahRB0EwSpVdf3FkVjUqkMdaaD9hohuLFG/XVB/aHQglLzK0dAcHTY
CY12Isou0eZfFDPpKYRzDLTnspHaIokcqQzzt3+92DLuMjBm1Xs71PoPUr3Ip+oNddMcL5YaJHhC
T3k75mVWJ0fDyRTbdBnx7FdLyosOlx2Pv157nfn10KX2PhH4a5vYmqpPEzKKZgfkpBvHEjt8+KA8
hA3osdymVtb3tiRFF4ohNgw3+/kCveAybt7WGpWVLnX+7+Lq/FIFSp3e55DbhjyvVzvOovk8Io3K
+38mlX/dQ0BFLL4XqjPkk5Z2B12xYcwrlh1+XhPhQp4S+BRBes4cf3i7eURzwPki5OAJzFzGeltg
Wk2YBBCYDhhGa0K27GunHFoh+5OFcgubbB8nRRoGsHcRf993LL9rtUFIXgNYTW/ehuangCuf35mW
HCSeKnhZw30ZkS1F2mq0PIHitEAJVsHe+FsXeBG4RAuxcHK4iit5mR3ZLrVftCRVTN5XfgP8gwTm
2ihlxNHHXnul9B+35dcqVzIrYis+7yavUWD5LfMTOZIeujaoPr5WTi02KGjQrWTF7I5Tg1cGMUSb
+SFlsgmmYKREgS8NsUMfC+99dCmr7XF27Z5bCuswIHPT3USvmCSKFYyEMgo6mjBUvPpykQ2sSoCF
TqKzZAZflpiRaFoHwQZAmmrbWSSLsCEHXtn58Yb6OeIXkguWvYksoqv1f+x1ritv72Lff3ljizWe
jdS+RxyxnL9ouPVIzwESATLXoBCKXsblRrdiYe6t7Ioia8grvfA67Ixg0toEoJ1FfQxSRqYjG2jM
SjAWejF5W2U3jjavKsV49Fljxq9Mz/g4MOmjTbEwLlEy6U8QdkIjoesKd2gPGMTAjAawC6XZfxcd
v9NXmwD5BiFCA2KRKkUndMH6MZ8rj5rsyHGSiL4D37sS50Wy/QK/b+/DXsBTH3q6+ydWq2JEmh2S
I052Mi5tcN3sdC+mRKbxo7hMSj05UarAbfHLh+VlPK7u2hdzIeDRhsrSXUuGH8U/XZluHQI4Zgpu
Y3Ww2O7/AbX2yJvAUXcXY9h4IOeBYyokXnMmGlY3Yx0WXwZmypozMBWicIVSO80drsChljXpCvZr
v5uyjfo4jJxgLaEbZknshOGHS7nxQV24vIeZWV9td8Wo5vI8S4Pu9Wcwprf0WEh3/4SuPWKxDrc/
6G2/fckS4yWO6+WFo5Q+mRWS0ZwkcHmYL1F7ZZzZQvKfFmKsSB4ZJv/Qlj5UN4c1C8niP6xUdBSE
/oiOKl85E+hiaifkInTIv+gLgcD96LDVqBMjgA6ySyb6AfwkXvSBVgTOOfFLJWue0p8yglStx/fP
e7TOOriAf403ZC80iT0T/C2URP7PPpcSES1nb9JVR0/p67vcuA/aB2uWi2ui+ETg5pcosp54FCql
8EqlWLglQGd6mBy8/2ghGnd5SCK++/LjjiNFPUTx5GnmJDLK6JRKFOS/vENPA2liP6f973WAJipN
JihsZzKy1sU8F6F/nobPYslYXDPqEUcUERZUswon3PDlQZrTAcqJFNh8eaIciF2mtlM0rzZRZqeo
A3gHK13zh0c2GpznnzVzj3LYZE+WWxb9Vsnhc/ua9Atn1QcDLZY1D2lW1rnHy32iqfYynI0bhXkN
/AMXgVKJanjg2QMJ+8KuYB/3i0J9dYi2TFyJqURbv8VIhe8CvVr+YMrOY9J02XhGry0IK24qipsk
SdMB4NSxwhExmauPFofe+QnBEznVNAL6osxj/0mi4HBHY1x/mNAALCLgMm5iJyx9NzQRsm84HYzt
i/a15M6wqmxASvmlE2vl+qxsFURAn+er7wSaDXMe1VL7n98FC4M5MytMUx4zh8ldbMa958vby/nW
iukSaz0LYz7VAtJZ23GSec/WLvo5wm7tVeyRSWg6Dasuba/7gLHOihRwiU5vY1cVanqlYvwnwZMC
Cz+MVIkLuf28qBtlAvehfu5KOCIcxKrJgwkyBuPog1BrjKcZdd+xgFv8wHxLeAwocPzg+n8h8RoD
IoKHztE+DWZffdU0jdxNME7RyzRrizGCh7NmxTOuKcxoa6sPohDOvubjJzJgllHPQ2jjsNjTJAVy
LmTTvHIBLjqvbMl+Obo7gQMX3t7oG8VL2OUOUweixkilAdKqXC3i2GSx7sEcYuvflVcUElFLH7XW
keLcc5KuXhziPBOCRxAC/PGuDav9nfFGK3qtS+6kP/ZRo+G98Iv5s5R2Xt/xcXCJBLZ9mswp5eff
h1UfDF2S09vFzFMuvng974ljqG87ZuekZ5qkeVzJRWksTvPkY46i7XnlN1IHM/T5vI5JnBKx+h4h
WPtB5e1tbyFQGR3rxAeHaZAwR5HWCpyx8YoNEQDrjMHSrG5M47RUxaLZ8XA4tbNTPxrKBFGdNCvY
4Fp3QGIcro02vjwGRIWuNS22Z1VTNrPSh+pnAQKrQFJKnmAdZOqfrhak6Pl4Q+HxmY/Aa1dNlfPW
zt/jYXBhIGVRcN691Z7WC0/Yq4WlrI5QAlkYGCATZaMgO3Nk8jiGdlCWTamTYd6xthKUL5z69ijS
Oa3gN/atNwk7RO1AtuRyoqKMLbTiF9lDXVnGfZKH/DjWpiVakRpm71b0B0N/m7fs/STuh51nQv2N
NoA1fWaDdB6/sHH6OhQzWZeR1I3NBFHgVdBdBdi2jfd1WjHl+k1QmIxx2Y9dP4PTCJzl4rz6AxoJ
3ynEI7+s4hA7AbaUweHTI0vsEOytDphO7tm6G1GAs8F9Hojuqq0ocyUJ8M00xNPQavu+tB95BQj2
SM6pIev1dOAphL5fLE9faUgSLBV8PONpi+1vU+FFtcR3Pe//FBx4soE4yyZ13jj0VJyQGgnXwfxc
9lKavtzQu2NqyoV5/+hSY4tTE0sCC6gX20XUnKcqdSkmeKQPptTcpTjSfzYSY0LJ3zXNGpOa6j4O
6jXDzGzTVAHBMkacIdmNad5XodoRIY6Z8rUD0kYXHGM6a0FRBRvQnzPbamG+R3U9df/C3b9+sPOg
BWkLl0g/gBgokyvZby6Mm8i4ywX+YakvEQv4Fd0MYatDHPNozOd/rpnG7cdoaKdeAgH1CZL50vpe
J+lvhXzYeNVNZROU+v8GV3COUs1oE2X1SmwoYNPDjqWsNp4wEottt9bGnK/IYR8rKv/gVgmJxelY
MyF1siBDz4Yiegm5Qp/Pk8HkmyvLJWahVTHoaIelvPKkWgPe8MaptnbIjdNKOl2Kd0hesT9aBVyK
TrqzBclYRP36FWrbry9iroLVOrNpmZ5vFgZp6hXaWGtspX+7HHzVemRqk/hJm/PzpGgFwcqEVU0S
VEr4zZBlHF7XoF9JjojcCG1+cjKmI8LgsEuwI14BzeDEru4X7bhwfMGVuAKd6xPHajjasKkwcJi9
svOlkU+nM6h68rESmNoQ+5x7Orcmji1m8xECn6mowOIKJSezR5yzFi0fOrkaVJj8cflQqLp4nXNb
9Kf55gm8S7v3PgOv/bUBneZuo8RQd+Q1LUKt/GxwLDo5lCUkmgn3512eE/4Nm2D0EpIJuEExbCAG
JbsZOzjChwJY1b19DHRuqOvj62x9LArUORWNYyfHhTcnfA9OcotKmOstZdSGowbsFuhH7ZY/CicH
0R65BakscuwJULDgqgwS6BhMIbsVgOw9K2B+BNXw+87zRYJAMUbFzKpHB30DzVzYpozThE4llOds
xMm+k/UFmuNjiOtquvO1LNbBBFY+4tMd0BbXwPOVoaRhEC66o7TL3C5+Yo3t4Fa1GcLze5lsyNJE
9RHAqR2iYFkTM93y10wFa8pyeB0D3xWqWYotgYDJY3geQULBKskyr3K8+V3I2EE7aZtIHPGPT7g/
Eugd6YhLiWjvrmqWwB4CBJv0xW5XtV7cGEiZQhHD9SnYZTziNj0zFQte+GG7ZHM6g4XcvYHe15Is
8BEJijaeYS6uTYh4v+CyGPwyHagfUqy4UVjtKzCLAjY+KgB4Qh2tg5iffgD3NY/sXYeA3+7hCEAM
lK9Vd33Rmp6IOwvnQWTFErmEhA8rF9QrxCy9qeUX6OC2ImfYsldp5JhhPrE2Q2f19lSynSqbFSLp
OLXzltT2nrLFXJTy9fu7RGIUTN1bgeUlnSNjJOVBXTsRceLwr7v0KMeyaQnYqFT2SLySuKLsvBaF
EtGsNqziyeN7wlKg/GqHvgd0RcJuJTBIyhxATq4cspZn5LS1Jd/irgHQtXaJ5TqM7gEiiet0P/wA
9Slb+eAD0HEzz76WqTHWPf1K+EVW3RhmyOHjErc4csnDdvkd0wJofk6J6N20RB5RoAoItQ/gFTdc
jOOp4GxpwuO4KrUYl41dHWeFrszPmsTE/ZIqXs6HWR+vcadUu2ceKzBUDNGnpedCzQCQEXqh6YDC
j1m1PfA9FIb5D5pZ7Lv8uI4RVxYZlk3yVAAQZmuZzkwFzfv9K2igPLEjqs/C5DjE487oh4Q+Qd1E
Ym0RsfNR129jToPC60U2vJU8LtZkiLKJY33fcC/EgbQbykVA6LgEZFU+td4vVphyR4xzY9stRFrO
pTnTB5Hdeeje37Q0Bg2ItZGpxo1YpsyvPwM9LnQDNWOEGXmb+R2jlZ5cZCJB3f8+tb3MYYWEms85
tXm15LA0Mm0e8uZSZFmxou2xpL3wvm1g8Vsg4Gz0oRSTTNhd+MVf+FbaxqsTQp6Yy4hublCEU3qe
csTc/zWoCNA1U0knTDH6USZGweJH9o9VY+l/DyE4ZpV1jBcbH9//nTjUJu0MuzlT7jyuXVHDwXzF
mJnirE5XuwYELpBqL/HMiqnpV55O8O6GQaEe8vrx7fQKFo/r8lxomKjGEuZqB2/tdEYYdLhR2ecB
8oo6wwTzQvOtUV2nN0f7X74mqe2NP9x0nSpxdPKHFXc6+DIqDCQt/J79JGLjX21C4LFr1X/j9cpl
qkmiZaGel9Anl8SeYG3Y29WSWiJDDqo+FSoDX7djlmrwtRk2mDoS7V02n1L5wZwYrPXchepvJQmL
U+27ammzJONOgjNZNaeBn9PtJLcSIF/B2uPh0UDSTbuMGzH1shf09BssIXoVoRCOdyM5lLJLFUaa
Dgl7ElCxvljjTW+vvwyhPEfF6jBzkIaGflXdMhP87b8DKFWhbs7YmIIHa9wggl0mtkLU3KbH3zAg
BFVvcL9/PFQR4i1q/4P/r2sNTLQ1bIGExKK/JtEPK/vyELy4fG7wcS11VtfdGtOsX13DqucqyNvR
VGtZQP5tm2etrfT64K7ECVT2r1CkFoXLSJ0BvpZVoDfoRwvsccmXW6zqNvvO+TFEpRBabpE5ShQq
GD87RPTfAKWzBS2f1DJCEF8hKfNS7QQSUS3cC225vIrf/0vb2+SPPzN6eJrEqe9vp7Ewt/jiG9Cz
kl80smeQfo02gZ5DjQ/Yi79HhKyje0tnD1gQupMJw1NHOKTx+rVNcNQxG4PZnz7mcjuZs1MMlbvZ
NTpS7US10CsKti7d5GL4bYQ/3k0iFhmRbfIQiLLB6aXzga6A5Q8peB/lRWZCpvOJF+DDDmUJVxh0
mvBMgyj9TeFLV9ypUrxzRFtp3x7GGf16vRsojVi167Rf9DvM54eb1i7kF7D04hZ9HsdtYb6vWTHX
087qJNRxSVQU0tOt70LOmmaQo+8XhujHsqE58rLhtBP+2SUv6hMIPuRMIPYsou21S9o8NzxgxzjS
7Ye/++Czs3fLdQZ1T+xCjUBP27IhjgICfTVX8O/Y0UcQEH2ZhjKmMPBSyEB6/O31kKLawRUDFbyJ
SIRnsdNl3rtT0MsrNRvKk9rA2+Qk+C/sGBjVqrNUwPuzwFsT94OsTRDzQOqSynKIo92tsIcijnak
J0RG4ySX0jf8jU9mGjAdfMICAGpu+LmQNjtv94ZmFGOd7dRTxU0ftKFt73+yi9sObva+XE6SaSYW
nlJWBU5z1eslZGDSSAVunxgZ28+Qc50ggEGaBaDpKhbcEbUqPk/ix8qS+7558WUPI+6wKBqkxVp/
ANEZ/k55VzDwMNw9tbIeTOZ8T0dnbpC/U30atza9VX5LKhOrCZDh7VnuU8cogj3JTEmamdsJo9f+
uM9T8LtMY08Pge9iMW3V4eNj6Im0SM+ElQtWx56k93fQXV/77swQGd00bvYXlSXSMHGYTPOTs8xe
I9BsYo909WRz+n11Vb99xoKSDA01VWfHuF3jYMfTFYNf6TMEXkg5ch0PgrCCgoyGAn+BdB4fE9MD
jVXsBqogJHWdEguq8I6dFhUfrCCE0s0O4o2l3yJ23yotA/ZgAKbXRf87ac9+rCbz+0W3FoK6A2v8
M+rhrJsuoWuiy5y/qVjhrPWxGzUWp/v4WrC8FlZLGjirXJEKyoxyKsFyytfdf4KOC95/b+PKPGyM
bFqPFjl+JElGCe2r+uami4d3EXGivq836kxBV3UZsCpLZkGDBgIPW7H4CjOCa1VDtSxNLgbOndyH
NW/tt1M9XpJLjb899HL68xaC+I2Ui2wOiX5btPeSUhPY91w1YUyeB7YkIWFpt/HacAiZSNoh96Yt
DsZauQ3pHM37JwfKWTFOy0G9LXxqqW59gA5cYIJGFYKiBlFPhOhFXIRc6TPVLhd7kuMia841Y5jz
pLKRqvMpLOb/lsO2BAtUkSniJAJIWTEOWHJ9NPE6Q3gWwjkUz//HktLI/XEqagemjFr62/zzGYu8
y4NeIytFFnEWjZdzM9fvO/BPvfcL1ySya4QOVrUbqnpZHHDuLcaTdegFhPcPn1d1/ZzHQOX3Zt1L
gYEXNVLonkcNCDVH7Snf2sLz8QUhcvJyyYx06eC8u6YHf3k7TghUOZA0DAoTXGVMGB/iPE2E2HTQ
7KprAMtiRCrMp+9SMzYkdTK8Sx2owXYDYW9s3swyVEcSyARw4YnEEF8CYU+eQZVjnKJHeudEKToG
vamgiIbwn5yxLu6UpanVflei9tlLFEB66BY54UsLkOw9HfuHOz2BIkc5znHyA9RlkHPTYepYYwm9
RMqkdeoHfj9Q2p3eXF9Mr4FU3Hac7NL6DELj1AYWVPZgnLBxHHAodDoM7/GYB0VvVT/2nRptd/i1
x7u4402C0ZVq90ZKp60piW2RCCl/f3UKgH39jiHj7CSf1o7cToiq1Qyt6Ap9LFG/4tK0UrZ2yn9C
K8K1J7GSnmaOQY4TtaOUu2kAikuDoe3ymCQ00oukhsc638o1HVv4+j+yRTaNiLn4+yk89v1gJ5we
/opY0p5Yah9R6xGKeMBkO0bk9KRtwWvtnAh8PYNkA0l/EN703HGuzzJNctYcsGd+GuXJahqgatGZ
TJgvLqb7jQcKoKPET8UoJaFArfrpXdumrHE9TTHbfLzFUiMOR1JzBP9svCPqhUpNhQnY2upzxEVn
ohstfsW9sA5I78gjOU/kVwQHjNizVc45waWFH5ayN9yXjwh/jHKg/gXV58aQgG8ogytj95+K/8l/
62oYUQ5qA1DeFlkPlu59uH7+DbYG8xLfNwT4vMs8ipo522Ltr6js/DsfG7Kv06eRkkCArW0zfaZ8
QHub0oxtG7PpEtz9xJhb4lLtc6akbi9LDpWSt7m6Oe12Q0a9caB442jYtDVMMANTEFHmQimgLhV+
hW6TXltjMRy80/ivVGYHBzUL53S5w7e2EzNYZjUO3yPAQMW3FbVJoHV6IAOnkI3LzJGrpHs6/Va2
eql23cAdDWlj0vg/ZiLOPd3hMPwv6t4vRv4LLeprrzOli3Lv2ztNJDFpDf7G1rT27VZchTITc0pt
7aF+gM1CoH22r9elYGY05TJYOrXQpiyIDMlSQ/p0h2OUbvt0TrEuX1kaB3/+Hi9P9/1JFwvtRDlQ
JZCbwF2VyHwPNXHFEP3C6UI8Rifn0tlKCNL18pUb2vJvv6YVy48AJ6yraV2dfMiouR54gwAILhcF
MB1aD7+LhOkTiAQ/O0QVqhQyFqLIOkqmvkKJYOtLJcRJXacCA2XSdilBETAO0D6fI/w13+2Qbvq0
3CgoqLAOHmxTtejmL0ehgP+TSVPt8nEm9M4LXITrdiUn0T1XNMN9fVFBy8fJ3o4NfGJBgxUcAqPk
dq53EgPxmllOpHt8dXLx6cb2SJakOUbSNT17CqGZdV/khmqlIJrNpOe4uCe5rSkl3yveojqgkbfT
K6PMRbpuAllWgyOOcBhw9LYJSHuQADBlOGvQCJHcgti/h7zP8569dtIKTV3SCeip8/nHq8/ZLa2m
nZ/pqbm2c8AHQyMS7V6+sCZYap1rcKZJDJXxJZrTEyxtzxpAK5qAbNQKpev1yCX+2auwuJOJ8Z2E
AjakUfdcHqxqVU90lyHsQC/mNEXa0knnmUsq/QmKpck9izo1ygNnsIl6PLy6jvEmlGSoOJTtU1Qs
f2QVcKm2loH20C4P02OqjWuy0J8r3K1jIi4/8MgnF1Ysc/HA8zsfhUSBL0YypmdpodE+jwSOYCsr
yg3MvSMnwAhfFJ3ru9Hy7/bZAGVaONyDMo+ohQ0cU17VdpA8vxjCRyX/tT+rNh4chI0JBumdL1SL
wgS53afcS/Y3fth6c+9GZrYrWeckx3bu29sG0wrcoY4bSZgaMmZHSPcxHeapcW1WGSFekd69eX4g
qfEyidJ2madRJhSZ32YiEviX1RlbK/Z3feMr6X9MnGpxyv3mgODFWiDuYud3mgg52/4r19bKYbj/
9ejD8+mIV9fYeLFvfaTVug0ybVlFJMpB/wefNrCwh9UXzwAGY5iUC2+wi0alF13PhviyVLdo/ikH
CyL0UBB1ieqZ+qwhjEgZ/ZVNhSDwUY/6DEdjPMNTpv7vRhfPImeAqxgQc+snyCK4KpcBE1cm9Mzm
+CHBnrUkCj6iYnL/kD1sK97Nh/7I1pJ/MqfqGAXqUKFwJeR1BNu3YGAhrEMOkidixrtf89jdJ3KQ
eOvuVxEJZKAJgjANyjXhgxzuFIjyYuOiIdDlN4C6hxZsz0NR4dcrSAD6M3Vr71oX2yB+qSCLi5HG
K1XF/yNsOQADh4eXDdEDvpvhk7UhnvVKXo14YRPmvi9T+nhPHaJgsMeGcbddslkDbRVI1fJrzol1
osyCw0Z0Ua+LU3cBYLsXYfaC7/t6mjoaSHUOZXgtNECiRd+hZa5zMNd456pF0lW9D7DS5AKiUXUY
jrNuARXcDqWQ5G4utxjwDWp60qVcFOfKaaWd3KHVBltoKQPMQFE3i7k7TAVaNKowPiKpcD2MQU0l
/3RY7vX3LoHjR1iXlOrH6U+WCX7la0NOk2MKCkHmS0DD6Mzbx3/lzb6vVhp6UUM3T/2BWoqZx/IL
FvR24wNVBOJviKe7m4xqrGUVsSVM1HY1rxyMRCmu+QwPo2JfmVPAc3uoHAkp09zwOxDuMM92zqYp
8Pa5sNRQJdNmlxZPeuz4/I4s03CN2PvYOMAQHP0LGlsy4KhCRJUVIjdzzDm7OBj0KeKVKV8GKMlO
8x5QwIiyScgCRNfyh2wVWku6Yyu/RpGedmgSHJngaIzOAqkPDM4syqcHxQzhhA2Mf2bSEvDCwA3Q
F9BgVkeUy7VfosfMxXc3gbD9eHjqLcH9fdmXf/U4xMdO8Qho1CP08+JXD7wAmGpdlRQCFw7ojJWr
74FiiamRvrveeVqt9yf9PCcQcyiUWdYiNimF72vML7EIprPbvCseZgYWz873MC1QfyI6mko80eix
p0i5OxxjlpOvx0+pyzJT8TntCCu8CMA+mSMx9qr/wiISZEERIA6DVgiUhxK0Znoy5Bi4TqqZYH40
zX1Z3UfXVr2RPk8hA3vpojQScYFUs5eheeqozRNwD/q9W1t/hfitXLJYGTRxea085xasz3grXAeI
zypbTkiDBb/+Po1k6WWqKCxACE4gJ4FfEMcNQBjkSMKfZ8LKIT0PxVALmhJXds/0slXKtB9fL8hC
xVdmotKOa1Vh1myUOI+zfvn3Qjm1/M6HHAYD8il4DEVzTCs1ee+edWdWT7Av93Jx6ryt8NrGk+5P
LE4IZmr4ZKnWROs2uAQBrFZoslgH+OEzw5NvD6UedsE0mf93cSRIlyoPNNkJDMzuMeHSmJLNc4Oz
uzD9NZQ3+Jw1njjb8L48hx/3zohIzIuoWd6AQIPOAf8fnnCiMPNp6LP0G3fW3JTCQImWtAHgVIWH
zhl7/4Phhrp2ah+BwxBABeviD144Vkag9I96AIdiSZfxrQQJWExqLo7gaI5BAP63Z/Sznb1IHioK
6lvjqC2BD80qbHLN4TXII9glkJsSxRGUtpNIRI9Nn8xCLy06lZzQXZU9TkoOGS3MCXgMAvBVLh4k
RH8ik/gkybGb8tW5UyKgqDN5oVqaVr39Y5FqiclRTOIrWVwtFECejpCE7+KjAMT/sCtPk00o1+pm
LTvcCxlYpKsEpHicG5Csg+kSFxzNFiZoyydfi1LHZg/tV/tc80p9zfa9d8c+8p31+DdoU43uA+w9
K/hGspHUwihWU2N4APfQpYAhlFYmnIeXfeLuLUieb2OvOHKzpPTLWV5XLbpxzDgV15aXBt05dMiF
kgrOHjmsSC+CviBZLJQdGg7r8Gcq2vEpEEEWGXCq9LnqUhaU9R3WtMy+q0HjN6V0yArcsPjnuxii
9E8p2E4gRuUs2ePYjsW6Q5+PlxEn9VoKe6iA2x5cfTs/8rSwDnKnHHKQW6WVCgse9BC5roh4m6M5
713L3AhC0PusQH6P4G8Y+7Ya4msG+aCeZ54pzwzoT+XVztIAKJBVYdJlmb86jV2UNP4lSBwv1rL/
ZNW0eKpksBOwQJsoUzsvnzR5o3QJ86ImOoaxa6PZLekOlrXSGTccVnyD2yGUuYjoGO6oY+MwsjkK
El7cgRWIeQPtpVJ5zZ3/Ui3vx+unZaLLfXnWYtICUrzO4nUyaOfS6ZxVMoQyZuzZqgn7t/kf1TiF
JL+peDH0yNDTOL85/SvGrqi/nfDTqDSSxACi0Y+2Ctg2E/oqMWRS2e7Wm+ft1DthGK2UrUulkzdp
/5R5xQYzuWvbtqrLbbHzof+uMN9bleTzkZplq+yJ1D3HGzgCzMswN+67wCua9EFSAkjBDcm92LSu
UW1g3ukyQWCWeMNlhUd2hHMuWMxzkdBYBVMmeWiVrmKA/N+jF5GxeLdz/DUB7sllbTYHzmHom4aZ
vCEzcDuTj+VDdJWCXQe1TvroN19AsRNzifnQaNEB8LC0yFSpYcdhLnFeL5BpsCUufQ9PlAQ7KR8Q
rKIpf1oJw+aDnVj4STFLgH2sl2OGKzkaKQbjadRwjl5/xQddvJx1wC1oWmL4m8OQU1E0PTMFPEy6
iJPkdqhevF46gBdk5wTD7ovqd0b5P+/km0/9Fm/ylhqhp6CYABXw59kxugLOnEcO6peQQ6tvlF1N
y0AJJoQMuCkQXbNuiMjEwijd9Q0ICEYfwkX5xNog9TvKNbDCgCTrfGJKAMSMFEQOBUBycLKzWrKG
pmxnM7AfFWQDXIk9pGgwv1SGgNGzJkkof3THe8/012zKVXOdrVzU8Rlq8dKU7R7htWJcKzveXFZn
tJ4dwPu5UzFvgWGM45jqM8d/TE6x54kpTuY58kCB+GMdeVdnPrDWq/FvC/6Q2Fi2tKr7A5u3Rnqe
NzCyYf5A/DO85UEKjpnlC+eX3cvlaBi6itEEgnPEKEfTGY8UPZL/Ff8Blkz3b9P9VgjK4cNyWA08
ok0K88yh7QFxMp2R8iImLughViMmroUkyM4ryUBa0v6jTNjC8/Eu4pql94GKiL/nq/lTUA5Ec0Kd
c1f4fD5BBpMtViLUpmFhh+LRYUiexdKuS9hHYiPNUbfUlEzd8S9tgJ1cLgsxtywteclwgoTkuc/f
XQnr45DKFfUPEQlLayRXzBn/b4g/ok4TDz4rLwgj2/0oNfiVxz7pbvEOrcNo99cGe4gBiXmG39jG
LrYMtf6pIHcGpRYxQZM/mFEPjZVvlwlF7dZBONBlfFvVeZEe92BhAPClkLAF3+mwQ38ezmXUhZwj
zgsF7MGmNy3Lki4N4qKeShHj3boedueZVH7L/OGl8UnjQYXg/Eh7hC31qg5j9YVF5eyfe1/aoWYn
Fpv98IleGO6uxfZCW9YzLY8LLU/1RGxGnTL+MrYYWeXvoSt3Y5pxmLXSF/VpogajEYI5sYw5wK7W
KIBZexJlaaz2dJw/qsxX3xJgaxNGKpy5mAMcO3eKoVNFpkAnar4zjXKdqSXE8SLVBbBjmgkJ9Mjf
NHN756mD5KHQBc4B4RIXI+0SP+B+jlS6W0Y7XLW/91UbleIbFAH6Qi0t75DBXr2Iwee6h81kXLd4
2UCOMLz24dLu9ID8ah55F38xlhM0tx/t1rJWSxsjI0ckE9NmQU55+0dlE6p76asa1Nhq/fHGGP0W
HgGHCY3LJD4cgjpOsg3rIP7qhTmKHHSWPxjaEOE30eGGxMOy9KGjAmPNzZ0/oJ4Ia4dCWNErAdv5
z0dgt6wzN4Q2DTXWlIUpKWeb2HSbleTJIml89DmxL0aaImLtkZnaU78z5d0U7j+2B7FMajuMkrwO
zRGDgACRvb70DW8JTyMKNHWSlsS0xoigbj9dF8reVhLSwZaacA29Wxk+yxXwXQqdWdjOBMKGE4Wk
oExMmqeEeHvim3DwkTkaIv5BCvSrfGSGIz2q0vd86ZbfZPjuCbeRNBw5VbPF1XJghqdsSTj+p0jQ
hWbwhzMK28VTCrnvSa9rpdDMw201ZRcdQ/zSYdXhDllEyh/3ax9BlOo6/M9q9q90ce0V/vD7twHZ
SHhsxT2AoyLFBUs9XUb2A+ts2CdpEM5oufm0PIKCaOtgxh0XN9VLIH2G7zUmMxWumnAvfK7t12yE
u9yZujtO6zblTx9bCbp9pd9YnHVowbKz8FtQ+aiO6v0i0/CdVy8hJZ783Q+ncbTrEnf8rabgJign
xF+8SZuxZaeC9qv6++ejYdp6tgvg01hgv5CpjNEgrJ7eyb+um9Jv5yxcHJ6dDUIEfdkqaaiMLIpE
M51mV54uv7ElpoW4RjwMZ6itFayzECTZiOZZTD40NefyRqDdp1IBINvOV/MH26ZEsRmv7ockTho5
R4erTokXm38YZqfoidslCyO5fHrEnHtU/Xp0Z0JY7oBMmqbtJavkARXRDamGl7pp2AcZ2oQfOalj
WO3N+wVPJJUzJueRj3JnsfD8vVNL6zqrFMjO3KPGtC5KvZuVQd0wT9bsnLEZ3yO+57pYFs8dWK68
CCLB5w5HYe3piV88HM3o20OIBD+/DO3Di+4C9zDKbY59PN8+BZgNZkP40b6tWpNILVM0+km66cnh
EVFPw1UR6IxkLsorWK1h/lGNyHrBzjKYcAuVIYBiNIBj/VFJo4+Qy1wG6s76rrpUQFIpp1NMo8RG
HSGYDWsGZ2ICr/cX8uNz6qwrAa7ZWoZ7vufvwZuKcMgcPriKWM9aRuuEQ5l6TzSkfbCXWjsV/t01
0IcswQLNU75a3zvcS2cNyWp3jzF90fEgnTrHw2eSwMDR7uyvCJ6r4Zdp0dTl/4AiFK9c/F2cz6cz
3HCSajbZiUXGZFiNa05w9Xxn4wyv1resxkhSGoCjVRQCVQ60Tfrqf6WEfsdxUEsTEhIUaQDiCfrn
YLOKDQog7Bweby3Z4B+7MoiaSuk/iP/MHZTmbGhN23Tx19A4JNgK9zcOynCBn4QVWaDCVL+yjQJP
8K0thrzllLaqmXUdCi51BUM8E3FFpaSEyQdYzb9/7HQeJrU7HLaZx+4UGyHNPZa4P2mnQxudsTqn
bAWEuc8YZlQ6AF1sMsOwrghRQfZmbIfZIBFXpFxSzO/HrOrPIIPVcBzSTsLitW+brfmbwokf+HLW
8r0thPsi7cQ9efKOaZxH3JDpGQW2wISuMarFYjiT3r0YNxdbRvM8xuemwIHSE9wDi7AsvfMclAWY
h1q1oFGdL61ERYsbJa+hTfQXzUOhkDepNmfdA5feZ3uaaBWdt4wCj6Wno2R7a5Aluu2xe1G5HoZw
RUHmsqWd5Y4tHSToJSUMPvnb9Pq0gK05sFDhRUxhl13EoWK8gChj+b9NcD7mk51Rrsf2aN71KprQ
OIBwVwKfPpKSCJcJlczmvo55dU+6bv8vAAMhoe9Bu3ZBnbQuqUh6qV2XZrP1OensveWpJoCGwXmJ
BBVr68nKdUhDwujhqOmcFeyUhGyz0kFoRUm9g1UY4ZoMOkZgT/z5LrtHXgDZA7BdSKFTCJg6bZxB
EB4UOw+xL33J/bKRPibtSIw7Ib6pJmGGGHuezPafyW/hUgu8/4EM72Q3LmC9BDIt5tClRhn9kY3U
kaO0Qp0ER+EDN4ZqMNHrlKcHLAfZyMu9D2XX0PCiPQ2cpzdruhjkxaYg0qPDJMI9e4GYrmb10WG5
E0gN8XZhQvdst/ziaT5DaQgu6fhsrBJvTigucFUMGtw9A8Bmpys+hg1ICnTzawz2WSRHE9ka7pOj
DjkISXewC6nIEWz9pUhtTSCwo5pxOx9vXb2X7hoNbjrlR27maVXTQQyvjG1jGQoQe0dONyaNDhFi
Wl4wv4kR5ZAAUo1jH9msGJs1jWU5xGGqLX820uadEa2/cpT/j/rOXhdPKZA4CqxtfoSyEyYRHqrb
IkTkT2OCrXYK8R76UGdu3GnlOk3TxhQtlMg/KPQT2U1FDz1MwqRZCuMq+9gLcX51zg+LmsHFXJR/
KTtL2oo7jUgx42gFwSb5fCLDCQKM6hBtRDztw5c0E3xG61PTCQ4SCdGH9jKRENmovFTxHR8jOtn/
GpxG9hgrR6lFs0SQ5DgACRS6VTYMuYi7eV/RZ7x3LxCT83hxsaVeOmd0KZXdUKPJao4rhhzdZVnN
DTI+aCYci+E7FnGG5pMaicRhkQEKemsKsfncOuoZoMp1pJChbBpVd00ssgyf67t5sssM+bzoKV3u
3eVehNbTd3tmkPdOqOag6E9t1a9ykb86O7EKKPXf3TXlZ3C1Z3dOUXvm1xtA07nVXsyZzUUqg6QB
KHBIVk/rWDdV5B/GKu35qDu13b88uFOiyjtLIEfZ9K2ROPT/zogMaarOcEGI2g4CtJA4rV4GYoSH
zEG5EKZ0qV7kOXy0MlEfW9bpVPTm/DOgiWF88FSy2VqC5Ltyv6jYmKNIGQ4Oy5filwFZgJDU7dEI
+KxXGDBI4zkV4giQuslA9H2Ri1y8S09eoe7H1CYNTkfa3//D6j81uvr7NN630VJERldMyVmIj9tZ
OBj+iT6Z2XBPC6w9E/3ii7UkA7nBfeiffyWePyj2fFhcmzF3jf3QhgNknujbT7eZ5ZsQiu1RBkZl
gzUT5GekqTVatI4eVH9lZ4I6gupNCoBbapSorcxpbhnPkKa82WHtj9SSJSNqEqswNr+y0PEbtWIl
5rjxlKC/gsB+o8C8ej+lxPY9FxXNC7MFMsb+Bc67rYgNuQ9aU/C+wZNbfiZ75/qDuZ6XR93fQiOy
u8Z2NJHfF61y7BT6wbXpd8sY/uO3UOtkgNqovMi2dsKXzzbMdPS9Kjd3nIoM7j8HAwzmjriEJZq0
bkgFysGD885SbKVETA/H2uOvXRQskOeLgT8w7vC7PK6rY/fIzLogEhX26ZMSrwxLAdFsrrnEHShc
rAOA4MZXggxZ77I+g2hoXiyn4JxxAXuDjg3e/SfpECvSFXTqHgsnnZ+lOMZ8x5ApDx5+/Kbpfwa9
PHZ2i3tc38csopksbCc4ooxtwIa5bGJ1x05Y/LYmNKuOOh33rWGjHqSsT1QIr+0XVyvxt0K/wyyo
Givyq5ATOXy4o1YZZ424vpxpRa04lblWm/j+hnTo0evVIV97AD0ziWXmgSSX05Tr7xjPnudzl2Am
ctrkyLMZSi7u88+Nr5IRhSWHx+FfbtQsqVDXna5vUZZroFqVLBz8IoirBFtAaaSYq5dqv55k8g+t
xEey+gSAxK1gZDuXhc/NkkC70sxv0AntDrHLzFDwrHa4mVEXmhxSq22owJYINCWT+oLlJPPzjYSq
4gAyYAACNYAZdSOBF8ywI5509F7kMGpiXMkyBL+STzITpjriLENNxi3E5cRdLwPGGtMjOhafj59C
qDx6prd16iUANrTTHee0cTikDIs/46wuLrVgPlaam1VUuQXO6p+HDwPC5/6Bal5y8OPMJSHW7gkm
o8/DcLYr6pzmq7axYZjoILO2nycCVGjTC6cchyXuIFVe5vuc+4lxm0Y3B/85Wwfr3QRmzWv2gyqU
PnCZ8jkZZo0Q8xfEZotULmjK7vsOjYkSti+SETKr+oQW6/Bkl2wlh6YUfRo6bcLz7CDIWSvNuNfk
tMLKbFW4IzbdY44+NlVE4N9PRzvPpES8GgrcdIO4EBYmm8wqhgqftoUq87pr4n3tCYf7cf5e5GQW
Dyf/usBpMqN/px4e+ONE3S+KzZZQMvD2hEfeXKPgMNjydkD9Rk/KZf7Ym5lodW4gjeouqYx7FjAp
shKL8JCBff55FrV2LwYa10e/I3BdAylHf6lTdImhg1DkaVCq41v4d9gykcaFc7EjS7QvL6trwsiv
wVLLJwen68eqUdfatX+NAAYGXh9VvWsO04CvLWJ32dLn+p51hHUffY/M7pECkQR/5y/W5TU3QTWp
p82g3TO67uNyEXTPNMPS1YKreXzQd8Ck9f1Su3l261LuKCcaFAs67PxdjsmhowHT+soEroSm2ulw
nzkdchr5xnDoeho4wx5nmuzLTJCCTvexYas7H475Xxr+fGc9ppSbNk7uBiwHiHbC24bGYhoB/AWM
IKhQ7M6izvjHtRP3eHZ+eop3KZvo9PMYJAz/WAK2j5vsPZYA4C/y5PDK+z55GcmJ9dClm1lDmfO/
MF/hID85yveJNcWBMSTb/MBeZSvHe3lLrPvtIUJ0pUooP4oukAfRZYjEaLchOzsnUJQAc7o+HjfE
gasxsJ/0Mrtmy3t6DoO11OCec6cj0EtEoo+hwgc1H0ijbbZNw5DP5he/N2CW6XjuGhx/nN+gozkr
7bIs3KFrept+Yt+dNwc5vP2duDAgih4ILeXXT/jWPDQZ+O+qiuEdBzl+Hr5+7tT3isaZCfPX8Ebh
yG7qpO5NGyDuyUMWCtZBmIcRFREz44VViirLeggjswzCjp6DECiCNewytEESo18HlW+MXozrkBSg
BJRNsu8vrBizjnZ01FsOzq2b6HQOlO2EWBEt0/+s/hEAZXExzfHr6RavnOGgbUzC4r4IDldrYTaS
OCtRO+dsuWGwnDGOJo/gscLGQCZkjd4NQZGc39tzPw6TgftMzPz/mMcu31pjT++1HwT7zevm0LD9
L3kOnlOWMBiIAC08JwPfffsaCy9VjsJukuAu1QemY8Jn/AS/28UiuhxY5CZW/MCVGqWhCKvP9kQg
qbpE1NcAo1/QQkE8W5RwPk69YyBcbnc/ycNww+f1PsBCvRAszoDgmShRamW2fASiUL7b3g0uPqWR
FplNZ7DUvPwFu3jh6rb3xTNs42PNRRUO9sSFvaqC8Q3xhOpiNSlxpA2RwD9nCqveWHV29SA8VOK1
850mW7PkhvHeDP8z05OAEVhjhpOxwOFAo1tIERzPJgrdIEq+vkC7XvXwPLPx6p/FsX+TYrne50KK
jT3rwqJZIwG+ogiVnOZBQFQlVUoMTWj6RpohVGHl1fj0HsSC764W5A9EjcjXGutGQaSfbXaypEyC
jsLQkZx0ZC3U11yx5dqQsB+zn1iD1naXGryMaaGk7eI88mkensI7X8qVvhOKMTsFpD3neWywGsBr
63labvsv3XUvMEdZcOr5engasqZ76pC9kK0YKsh4qTiodv+TkeU+UF11Dnri1LB4/nsNVkLHV0Xa
5JI58jYlaXSJRLe1xZ6BUJ3y0O5SvqbKE37PoQyQftJGMjXVm+8vQDkHUxjSgbIYx5ogYDvmBgCq
txcUsYYLSgbcqJEbW5CP4QQojEdGADX/MpnNkTKgNzYkIab7t7DbzYFNPfBZHu3gnMmZjUHi1BiF
27Mf904YEQJm07zFiqj2sy6ShQADfgGlzGhn6VV82i4QNTooU1oSVagKHdhBrWQM+jVe1QSNNS4S
d7njIfP4gMPVDnlMqXRIKsmYM4v8kV2QQbOq99t9iMN+8ZT1R1xo748Xz/J080ifPFG+EWw0KKd4
AlwpZErpCi2QS6BHPp9tVDi/KP0VKXyGWY91fsfYB0t9X8C64F0+zgYEaSiHyy61Cbb8Q35LiLbv
/JN8tbvMGmeHoF+y4dUqTczt0J/YxXfJ9FqqHytBcE7mUIL8iy3lC8Iaglp4AgWB4TdZGR07nNKz
b72HEFRwusXJZZi+t2zkr+mFj1LP+hsf5rF9y3d4aFWoHmHmS6fcbkrJ+B3JYW5rdS4PkX123Vi9
O9X3SPwoD8M1zjqdVu4GslVOn31gJTSJ4Ajhogk9B/78APFXuMEiE0fTWiNZD+GpEiMo38YSxF/o
9sWJwTj9cgrVkwzNIIhQl9WG2GEohdb8XYIyP8EP7QFRyIqM9gmytcKEEN+lN/Ra5OupT23nfgyL
hGxzyn1oKRb81hhRdYH8gtRME+c6SrkrPXyyaCaEdFLuTdmSLx3T+sC+LDtooR5+lMTIZjYlbpnl
6oDx35vsnLW7sCksE5yByKGmDIU4EYWUCxLazVOoK2I9AXFCGSHAi/C1LGbJEdzKh4Acz8UoA8gn
Hz67UqowmJZcAtAuqsPm+GnL709+pvIOiJ2YaqYXi20OOzOt/4Z1yY3lNykoY3wr6B9in9bjWiDy
/9AO5IqW4zDw4WVftERtfGD0/cwqUiCfAIfic7k1CTq6mFE2FACZ0Ijgp1uGzGU2XD7l+qqPqQDU
U68pv6w0yPBwPEoNU53LfLMalDMD02xmkGtBcgFJLpnaZLLveBv/ED52O2cWkL3dVhaJ8uLi+hZG
Z4D/pAy1DzsJ52dK7uT3TXx9Okxnqj5VcUpr1u9e59cB9c/wsVzaxaFhltpzJPKqlVzMx82ccs7M
QjulAMqszPgyBDkDs2IzmmjzpQw78lANKzldpwhfv8M6jrnsGeBV6lwsAXMMXsxOEHon8V/g8IJa
7pS3Gp2OADhbQL7/cky5r1viPGxEoXIOmj9ieFv6hj4wld5zKopSqhMFog1UXLFtiYaZzsJbwmSc
m5whzDF91fyznCZ7u2iPCHuQxcvjKZMOTDvLq5lktDG0qoH3kbZwlQcXo5fEqk+VYcxBeeiaP1YV
hl4tJhOVAuhLySF9RVhO6/mvWeSEMvUXvPjzJChxEcbY1Xp1DriEw9lDoKVdHd0aRmxGS0j9vIVg
CACGfBbKPWG9JSlPYGsZ7DeFslWp+W1cC/toLaFDarJSqDHdcohv8PTlSvFiJrVuKreU+heZlUVo
A0iFPqcIS7UylluVIa1XabIwhLnTXQ/gKJDro2auhWtaxULQ1sTbI9Lmtmygtw+2K4sRwhcOQTsu
q1PZPfur6TM1ANdJ5AEJwOJ2hK+VD/JLvBaRWE+EtlxmK5Vt8uXY8G6aD3z9g7hFG7cXVIvk0hFT
W+fB4/ZoJFnl9gzJ+SFO9hBGIK+yCoU1T3qX4PQu7K2jlT5C/Ob/fu0KS9qee03itWmYfSRiv3Sb
4CN/YRIYWC1S2MSoNTruU9ljokalVXTjASLP9M0GQRtb5Z+xjwH5Qzl46iE18nZrjPLiGXt1mXYj
2AwqZt7kxV2YVqXhoRexk5vMhD3XPVT8rw53SiGVDhFe9CQWJr60xtD0FNTSHxc4VX/cDwdv9Yqv
zIeS49H+E7gdZMizLVd91fnPCMxZT7KW1vOldxe70KAIJq+8vi/VIajXGCb/kMUHYht7971qDO6R
4oLQofWIOZpYcKvzC/SW+hie99+8kbEoHN/lwmSeNFIpOdWtT1zBsib/GA7fUoIBti1ZJFC7dclR
lENfbKQK9Fp3t2BfstkT3s41IjoyaMTn8Nf8gm5HsrsKtg29sHWFQsdGh/h2UeKoO5l81bUoJnMg
yzKZ7/6Ye2L/HjRF+RUGNIltQueVlhheHd6DH9xxbcWiDFXTY7GvxNjgF1Zr6ez5XvhgZfC79qdj
C4RHWqcwFuaPJnvzQsVStmHHKDcA09Pwm4r25jbUkaFhL2xQ61/Jlf/i7QTe1MgX+ie1i4dnh1r0
5v7s1NNsOdZxWCgcPW5P/D6e8EBW8xkZndn8tOuFqCv518DacGPy7LMJWDLxVU1+VY0AlFo9zXm1
JMm7YNkmiIN0+oFZwxCmcxgVOx/rwuD7u4pqQDCqzb5D0I37ydAuoSg8qTX34lPE6UqXeUw/dRH1
F4wpr8I2RAbPUQYMgnNQ1M4lrGr4IyANAW6LDmYqYv94duHYt31RYeMxO1+Sai8hMDeWyeaWJzmE
mf6XDcdoMmBUee4iLr51+L8Bg+43/ejxxNCr/kQPUzM8CkhwXxcS/KnYQB7vN6mQsJjNBdDYHdzu
3zkzm/wXHtyIq3PMsrO8B5sIdQhMedh6b8GtY64cxA2a+8ZrlhL2/j1NrSCRB1Y9GZejClJfbXXD
npBz9Ip2l4zh9tBRP+dGhQnfzkDXw3xay3pSH2HnfikBs/ysKFcs7FH5s3fKqgvgcEfjzacQ1naH
cTEYGA1+YRJCMEvR+hoZ1pQ6dD+HEDTJv0s+c/jpmmY5l8E74h11vOM1JzFrjRksUuTsFKaKpjZX
/3Q3/Hjvt6EPSglmP7MpKF075xmyryL4MFm2rf0O6R/i2/s3sjhqsS00ALcB8BwRaJ8cx9MQiQQL
LtVE30vxWeaul+T2+tfQyf4Q8y+L7A5lYv7K99Dx+F/nparUETV0ULz75Co4uslncwcUOKa1Ie3A
il2a7nTkS4zixx5iVer3TP22KsgwoYe8D+hfzRPcc5iXfLoartOw2K6E4c7QuoBAaD/DHRE9qo4Q
aJIRVe2Q82UGsys8k9n9MNJfY8Nf6o604zx5K7q0DN5A9cxPnjNQq1y83jUS8xaZrYuEvM3RbNke
ykbMwRH/08SlvZ+MnfE7LNXzaTfY3UNigDsKTusNNkq6k9wLMdNvStyMUcOz5skR4Mz1t30Pl6Tk
4aa6rInLmWDv0WZqU7JkKqyUarwwyXTTD2F11MCOFKhL1vPN2x10yczZyWnLv65/+V65QMX1U1gx
Z7trbTKBIkJXqXyIKtD81aB9cnUiH+G0bWGpKxVYhwA4buC4GyWImwVmrfn1UDHEcpVHDAu1FLqP
Al8Ugxl7Mg0WsMvKBrc+/lbSW3WH1haZgx8XH8NplCydyX8dtFLEBdTI85vzZTnjnl6o+S3exsQr
5qLZESzlyt7C3Nmh6gJD223Fgp5iD0TYgj/CUMtxskAJVOl/isrF9uFAUi1PkKbxZoLwhLegrNnr
vzqQFL/71wK2WrcMjDgJAjsuBvGFx7N8Ag5TGaECaN/PxByGPCzmWw95+PH4fbRtPqqyMputks7d
ekyaw9P3mWROAMba0rqYcH6ct7Otk+ADtDlCcEXdXxRhVbVs0iF5MIZDVFNV45LW2BCouH6nZ7be
6pgfo3oqakUrx0FYElITl+A6FKXSoRFbCvFs2GVIWyaPCO/BFUWc4ZkDZA+NiL8deMURdOR5p/Mb
BrASzzaG8mBlFGHJ1BQWExR5xu7zP3CUyFsZKafYbtgNaNWfv8S6ORnUssPgdVL396nLcxK/iNuE
X0Wfs2upCPQ7agD0XnEPBC2ZGdV8ERHVv10dIAb2W04JtgcYmWDraQCJWFTG7b8qO07Z2WHsjifk
i4FflhJd9P28O+bAI67qTcruJdw0gjzXq5lKlHjXBPDfxZXvixPHQlzRcYTw+EAXrpvjCQG3Ymlx
rTOWHCsGzrd9p/q+uSYRyYCiRAX8JXFYFh+2GLohfL97YeocYRK/eYGGBdX0BiL3XW5RjGc54qad
+cdMFVzpxjeyUPiJGzdSm4GAZYO81vl0ZqlYdkACkcIwHYxm+WpKrFapHHugPKOMO3p4+dSpaMOC
xKoITrDHbUjxKmtLqNGxIYNnPkyAF0O0u19x8tsOmXGsBhSP0UiUse9psJioNKmol8DlBhDnRHBZ
DhIAzx6o2C6TRka13O43mm7V7GjDr5xQu9x3Q+ufrimRy/VKmebEhfPfbMIUe2yOXp3jXfdSACkd
c1I0okYFgnnBQap28hELgCvK3DMLcE/jtZTc6uRK6TBED/e1Ke8EiBHAOhqMo3WlFcb5cu/CSBZT
Z9a9Yha+I/T1D5de+gSp7j1W0gw6SX58uVCfSWDaw32ojmsMDTVBKbh4lfvr4U3ZdpdWZkEwt0C7
uAocZlyTK5vE6wWNV2F3ikSkG3+p25+xzstUeE7DoiYIRGwV8Kh/29EoXxAG2dikmlvJi0uiVAZO
qqDEwThRDbij+65Ann4yP6dkbwze9Du10XbDDIQeGI6c1hSFbnh/OGy0uzQGrHNO2LicQ+b3A9hq
HtekGNZ5iQehqHqjNwLdtb0zzXqBUC6akLbs7p4qELiOB5trKkvEY4un626yVd9u3CcEB/OUIzlR
OdrFjp/Hv6fuAXZO1VszZsSeZff2rK4VjUQcnVGdfTzxYyYKUVdFnQ5YDcQQILqQmO/0bI8oiZyG
i9KLurUM8Avz3dYQA+LBYQpgRidc+B3n2uIuMiYCtZDwBHhtSi1CWRUo6m4bIDHnsg42rRyDysww
boj/PIcEiEVriz2EkeSuiRqQHweFVpSgvUSlB+u33Hmu7s48ZAISVVcHfEWK+mIaG0ma7T+Zve8E
YSqmeHHAALz3X+FV9XK84p/iSBQ3Hx+KEQAvNmKq5YfhorYzp9zPkmlOXhRbmnan0jAzTYBL9Rua
u0ZTlRUWtXbiZ4Xs8B38gJZqCEKChFLuXR191bf1ZTX/TrbuCAlY1ktNhVPJTO6TPDZH3FfMI54t
kgTMS/A5LyczhdBLmtS8FRAUyr3CkAu0vjgSNlevaTz4PhPljWc/YRgAoDWxZ5h7TKAj7umGe+r9
uGc5ArsQU8+ThrsR2zBJDw6G1CG5cwo8OkNBOSEGezB58/lBJ0hhnsMdgUxZFgfOAfE4HC4x9b0y
PM0vFpv5+5PfGVV2ihTTnGAAWl4n1+w4G9hLSaOrUlroKFGas2WkZNv0w1Jfwcb5biddOyGvFTOE
ESoZeYCzqSrxYhjoIl9ZZvRrjFHgx1HgL5kADovDo2qqSoe22mazLrEC3p3JANle98qh3sWR5qzb
jHev4BVry6cqpQ1jo44BmkksqjXNYAYNPcIo1GtnI1GVFDS6bez7b6idSUvWTzkeEYmxv4Zd18RH
bW2AG42eivdDN/0HZxBRwUXGNoOdKxJY+VMxQOKiICwqf6I3RjSxiRspic6IFEnnRXJticT267My
pR5FWD9EH8BgB+BLrPHOj39giE1kA9QO/RBMQVdDTM042905JvJwpV9J49ZjOEEqa9IgOOhWF/ot
BcnRWFxMWR4pHjorqiMFCGKZxkJRT8dvytZU5bNsy9Bq2gT0FkMPF1C2XaPysTM1G5VxPzoAJNf7
0EoqEscMfSez49MoJF3qmZLJ0fMGaPHWkljYJ9Wwle7jTTXYvpaDMPT8gnnCRsrAmhkwkxlVhQFl
qWjkX4cOoch29vI4vI5eRUWFD+rAf0DbY8bPp7QWnHBAzVT8GJiUH3dyU7v0QkM0Yf+TSgmSvLfq
XxsbNLHvVP1QQkRwAVLpcTxqjXaWisqFLLiSYrAdsOOGyHdMVhOiBzqYb89Ki6FcCwDP6+bImRBZ
VP909CBYZdzaGVw1MmlSUw4DwOc5ufu9JH5ck35VJapPSUsmy4Dg+ZQ3WMHujEcnb2GhOEYorjAa
2e5C0Dy2djb+I0JEPQNK/u5c+ZlwNJGsV9E6M7OXPbYuBHMbo+v6Zapxpkjht0cveaZ9hO5nazxM
aeieULR4Q9JzBhW4WFk2djyTHQFihG4gKLUDb469DkF7QAEqsVEm0/RYuKXdqYwuxRudsgq/K3kW
BE0WP+LFN/nbeoyMfAuN/PaEQwy+84SzWAchshbYR+vAefLfUljDzgs2rb4KEje02nTd61L16PmR
NObwuhbmow9UYtA+/CeLbVDoDwIsMMp6m6TG7eCjX9yEUy6/eMpUZNu01DxEGdLiqMojrBLx6CpY
1JhYW4KImfuOaNh+Ga0jeLSs65Sfjnw5Kts6xvJpnhs4WMy7bH9O6dXhKepXHQiS//K6Fa6AWttn
0UA/O+f5+HPpq4wEC8FfQxatmkqQJ1WnUIZw8bihMPLYRgeDnAGNnFON9eBg/NXHHa6SZDbmAlh7
HxUMDA68G9dlxmXdzHQg3tL3jXBKZQUgZwgB1ol7xW5qU/mMyKywcCpHQdLCTaqjzYT8mmHD7Kbu
DqoorWvGuOYOXnlk/TMu3L/6cw2jt3GXIgNpvsgCfRq20Deva6Bpv3edyoA7w0FBfDDkD8EDP0sn
gwpbIAnB7odYP/m6vZ/RYMCnA48eMyEaQQp1JLCeMEVRJoNwVZLdl8knLE4+h6DxnMyby3d0XZ/X
BBupnoX+3yZ5XqE8jdACGVuZBR9odtqqK9ETDuNyvJFP9hiOt5SCqWarB8R8dDF+zgHrgRTZ9ccS
BC0gmdcgGuvWcz2Lc/S81QMEVEbjGDigZz2I3DDhv4XhckvaUlXKUDQV4PLJhqO3QvXNJFSjEGwY
Zo4bfhT6AVMGuc2eaDmyIZTc+jg5bAFs+Jh734ZXrqJIw8eb01hzIoOzcQ1ZB/yNyMFeNR5JVTtD
8/IGK5Df7caLzRv5Xz0tPdU7Zo3FUpbH/T/6mwQwOB6FZNemP2FgDVSnjRMzSMN0uKR+3plzhXWI
moN6bsdt13PzowmMUQUUHZcGJW7RnSOUtnA58JNaxjSloRo5M5lyHBEhFuP/q1GjemgMdeOvyJLf
bH77Mn14FDs6Jsz1OVlky7olsIt424iY18MZgqfDmKxCjh+TsYGDBW+3szXBK+TNodppjNEznAvE
7DkCTuh8TffNrEF8vOgnH4qzRvrAS/e4/vKBlWfEWwVmqNcWYbFTQzRMO7FOFp4BeOt5O9iET7Px
t1FwutC0aPec7Dl5yUWS9goAg/Wvse7k6SmOnx2QvXn+T0cfTIL7JZThf8iXzfnaRDZKm3qZi3uM
Woo/SI8aGdaWCbiNPxzELI19HxEd7XLJsQPymxXWXl2fb9/cwvko6NpkLTVbP2wAlQPSfQWbUAx3
rQx3JZjk/yZ2qNtrbQsGFPB8iy1mrg0vXrN9n1NfdNPNmL0mSbKj0nvqThR695N+LK1YHJtU7e7M
oQ3mvEFavMNFI3oMgfeHVqf+drywSJpeT4Vfwjm8ynVdmyEBMxVdrPo/lQdq5UsCJi9IQPlub9Rs
en6dIeUbLZHzz676PkqbNshhZyWkEJ4W2HfAkN6oqvEPdMhUCJpujTYjvfAXWKfXqQoea6BIFXMt
XKorHwsbXefCN3382yoRxunkCfJT4SeRjvJVOIpJLRJ1KRS5byKUFjOcgEyfPIopEp7lDYbxAjMZ
sKqKoA33T0ZR6hiZEBVUfA7QElguYuwhMEAOJfv38IbrSNHR/gfBzZN0EL1MM8L5qzuo0whwA0R1
ryQzBnDyF8oihbmIrWhqUyiRYknRLwYK0J1/JH+YzDQ95L4nXtBCp/QnIECBxoABqqKL7zYwiR4L
2gcjHLXhMSF99418JN9Fyo1h4Z1pPXF4Vb3d1QEsh1XMNx7XOu/LGrTrUHG3ZgFEIyHkgZYKPDk0
22dRzlT9XDtg1KJIDL2Y+vtbCKNrNcu034WMp+KceEzBsz1g/9Z++Xvt+FykpmAn/zhkn+gXyane
OOPS4UcbddgEBWo4YEuy89NYQjLHuuF4nvACxKZAS1WAW+1mbwz9gDJc0jKum02J36rgv3H5jdPI
qai0S877EXlZ4CT4LhKIENPZxFV283QxY9I5OKKJysVKo8CmSPFSrKNRlo9n/DtRBr2Z88mIgNPm
ZE7P0JeDagV6Zfd6UlNIiHxc2GpaVw+WPCHA/8NZvew+fJN+NTYv7Yt7eSGhHNiddncirNUOYLcS
KiqW/RuOtK/wsDS7f9MBfkdwk0/GpyBInlDqvNWdsf+/3OEBGXc6qS9fa6TLk7nkBiDi0HX8mSfm
ec8tHGdIfLC5+IhW8qn67wXDBLEnOSvTsw8OYJtVFp6CKs2l+pXF6gssgoRPvS6mmNOIlwgO+uZn
p6vSLpUiE+5TJa+XDFeu+eLkHaV91rMESqcQldDfgfZLcOjyipS8hbkZkL5E7yfUDb0OSfC2FN0m
DHHZ9BShLmUJnCiY6YnKH+Tur2NCVJbqHac9rQSlkv84eNMxeNKtNK8J+3rZIJJoxHd6YbPGFs7I
jUunb33wNS5tlh8/TnjCWxAV7u9RuRfB8dkVTZPmTFfwGmyXyRzuNIYE91XK8IDMvyKxawlcq7Fm
AIF8iVJd5YDAK+MXL6oDZpKLO3e/xDFs/YfRkopV4mTsaVDi5N++I+vOC3SsEn7qCh5cmpMKrxrh
+1+N2NF04mvd/jvC+PwdQo0OqIrFwCkNmg1uMBntpxdqLFDyRjx1WKxI8ZeBtsb105diffab+Znl
QBO8kSjnhs1xFvguWDMFRJ5+xQeFqm50L34LwH4W74nOHcOD5CIbFqMRtKAALWxFasxwY6yPSSj7
PSxhhXHJlOJzaQ3r4WI/NDeRFF7rlf2PxLNfEUXVrtzpna1c/IQQIrZw5VAis2HzycG0VHlh8HYK
qD5Ok76FXPav60/voifhLvkooOneUvGY1YXF5GrgFXKP72kajpvk8NQAFiDSfh5b/ouBjGrozrbg
D57UyGHoeUElzVZZ+SvTvS095XbFEjBXTuDzse6AGUsCHo0hUQ62UWvhkGUizIAmy2xROSNi/9ds
YA3YxX2IZQ7iz4nUCXzXuPhToEI6K8/biwPRKRYh0vBeCtyO1CWpQcBqjMA97FalTeaMBOOkYfnR
GgpkcN4tyYhrW8Jutb8tLTzQ7gk/9dMyqEVegLDL7zVnzYTxP3UMx9YL+t5AaoAsTtAtQzNYjlEM
/qqnx+B5LOeRNnNOP/lP9yqA595pR3Any4L9ZNE1V9/xFu647eo8H70R1YhGXD7d07KmO3kblD3R
JxoPHsG9IEIAAzEjSqfRcM7Br+5Ncl3FHSdeuhAw84O+OSBLJN261OMiz8ThBm52nSkgTiqfp39g
LOs/dW1bGx4UctxM+fT3RSG0RsRhqTEpIYyOPDwqRfIAa8ZG7QlGGIye8rfX3ib8aOdbQn+I4TrC
6Cz5qXWzIJnE0NdQ3g0ebQKc692S0v9aiwVCM7uO0c5WzyLku73KX4qUIudGkibFYztCKHWpMfTu
slfDi/eNG7ZO6pR5w2Kgy932hMKWH8cf4Y0sx+WoIkMJxWJBwX5RBKJredKCeRN696B9apSqjSEF
VWfliPfMnv3gNx8sCwPsbo+XgI5ZBfGRMHwM2fq7LFYVOMKOnL2RL8pDFCDQl8+BJW7fiFwCa478
nFiZyhbUsbc83ZQ5g+ksgcLWCpzK7yiEziTexq07WqJUgig0vceVgTLE2EiyWq28Yv8vLn3/WzW9
jcLDRjYWijPPWEJIOkfCGKNQXSPVldaziKjuf0o6VBxugO53AY9ednH7Zvua13mau+Br30hsXTc/
g7eL8H6PDcZ8uZHpcRvunAnhAnRojEouS3VjzabkZJfuO4QjCpCKFiJVqWoXqKnKJf+psUBsfZiv
eLC5833qC0+7Lz/PVX0q7BKPVdXhEZidXdyFJEuuhpUVUM3V1OVgSR7yhU7yUWiMPbuKKIrD0+Di
yC/Hsyw9jmkn6hmjeb2ZDmZBwDOpnibGyPc9p5Oo5zkXHKAHYl+XgPWb9+dp4yVcZyW8XR5S/FlH
+6HdemvCS4D/xp6QgIfooQFJo+1Fhni45FxYJHs4Ce6T/zMj6oACj5oA1IueJApk5W3ko5+yqkvm
iBoo2qTqfnm08bIIlPTykYpAV5i2ozsHYOvabyvHDW7AyhKMstQPHcyADzW2rZQJwFsP3HeCRFak
VqFNHXskItpVnwrA5nHwvJ7uQUUZq8ZAQBVyUeoDQUj2m/NRdONyuf5AbCupxyj+FuO/3AJLf3Wo
qNCRqjg7Ag14JKRl0UGS5uNmQVSiRUW3AvYeuIngVUmbwRjip8kCot/3BmSaFEyinp1yWjuplVNy
ALcu3SUMTVTME6Ozk1fNNtruQfB/gMHR/c7Z5Zf0n65GxXmSe2GquAr9IQViHAdee5Hz6EfBbL1i
Yj4+FWffQpEPs7ueNEiRoAEu1we5Q7CZycDWEhMe1NZJT/+UVWgp0XG8vo+CrC6RmgU3UjVoyEij
6FNtnjMwGn+kcoN3MN1tQcqnydqM9Th5h3k99VocFphN+XxK7N4OEWkUR0glRwcS/qYlp5DBXFdu
Oy9s5Lm1S4pyoVOyURRvih2oCO76aKStiMNUcz1LyijcyORk56L4gWrkegZAyvgq9Syos4kLTFZI
ZNez7+I929WsMOUmjK9Xe6HKgiSIDuwSsiTLSpLuUYqHyLunrSCILjXoyybr4jHns/3kEj8Mnk4K
Ue7g9o/QSFlaHTT2YxP7bvR6BNLQAZm0zS3zCWEYfgdFsTwYx6EK326aKuMRWyWFNjj0b0QyEIjq
fCc4UJasY3HDzbvurylyWVf3XkqyrPTb/3XyQtyTh3UUJCCFd+MY56MIM3fQH6TE+LKQxzPsiQSz
AffM2dEk0sN0cA0T+LpQUYVAfeUscAw2snOLtL1vyogUsETyQAkgPnMMamVY4p1M5XIgkifywH5X
qe8rlsgwjsqJjek7P8jqFX/9xjma8JikIi4fwOwThxZTELjbaj2iuDUevq/3yNNXyBT4/niJoB3t
aZc6knf6cLTvymhL8x0+LFfKboNdgCil3doXWD2yzzjqL3lED38OriNoXBL4aQWMga+NfGQg69n7
QAGWc2lnK5+1jV8trrW4M2r04N632/saF/xySBkMeTGqqnh4Yhz6Y8m5EEdn/B1esFY9FGhFG7ts
OhcYwy4ei6dJ7MjDyvYCFb3RsQcu+ztC5bNVENOnhqX6xZlVIb1m2Gp6KNFacuPkYrq7Kf2i8MAk
EiDvnV2tMneWiARFrV6nzicOQvAWI2283rPoCoM8TEI/soMDruD+YbvyJ40Ja97SqkPHmjMIV6am
/oqPgokKn8GVDJ2k0O1ho5YeZrcqOQc3H+m6zm1PAjAFXTPl5l8RyPEfE1fOUMOHnit5M5s0+kU8
flEPXBomwLshqE2CuwHhKV1xJ5I3Ld/tOFgjO8wUTCuXdUVseocnfPAE3pHkGchWWJ1doy+KXgWz
aczXSxD1CTStokafdo7YvvMXv9G7SsAFLdUbk0a/GPFK1fgG0Hn4EatyKdWytnNzdn551KUc8fUZ
5B5bInKL7KKN6+pzyNJ9ZowSqnyeE3pufDvf2R5mO2KqkGSWNrMDFRaE2slFWZMUgPMnSMT26U9e
bpxwKtTmVkPCZnZlPyN396mDbMnp4WRmBAcjsj2f/g7aIqdLQ/1sEpiMEpjGRAYXyunx6+dX0QBv
RyY3UCVMWLMxK0WgCrIGERrd0VUDgF4NJEzrDUhPUJhyFTVh+56VzEDhMFtx8w28uztiQxbWLX8V
NmWvGtHEMcsG8LSWwm/1wY1h4RTJRACXTJKuTkeLLr6d+9MNoPHDs2vAPqDnGP15im9e3x5o0iwJ
W5XUzzPVt1mVluJfD6VvYyCkyIRaRaenIq0Fpz+YyAiwyfu2cCiLhmVwqWlaHJ9wSPfpjS3JStwG
S81+0z0Uv9PlcIDr6AVFIP6U1KP4Z9HyRtul5EbYo+ePfaB3om/tLVFHipysglvJkPPQwhj+jR+t
0mR5UryxsLUYESmBMuKs0NNm+VY4TPLdwZznun8+43aQd16schJB67kkg7ZuiD5L/046zslFmFJ+
TQBjjX0kr1q9evzo50vutVp5TZkEE1CR8PVR19sn/1TrpbP5e6Q6DHvN/31sLfidHgonKlHrTe3b
inn0f00DA/IR3XhM0tRe/Jw4GIZEX88njWoJATi9uCnkaMUVUkiPKyILHlzkBqtoZ8OOyuvj38JF
MACTLsSzAiIwTTaOayEilaQbZvzhrROE5jp8tEyrwZgfBjS1udDxZsrxfXPvOeejQZFEdMRMdUXl
BS31ru+tR7d77Lpd9rh6lhKGCRx897x6QZyWpnwNn3q9iIs543fuftZsamEMT9ARd+xoHvrJACSc
n/TxDfdysG8SOlongyzGs0ij5FGdo2D6fW95ZOnjUOizCrdXJcEjM7KzDnBK/dst4p1TAPWhvbwI
uPyFMuK90A6N8y9wo3ph2cDH3uHtU+Fyh5OwX8/7US+7yaxkiXuim5Io+rnVOQSkaXPwKdYUlhwX
4bP757L/QBQwYSnvsEtLa9OmllXjjpDqSUGj3o6A0k349E+jhMs3/NadRLcTN6jTcKeL4cCdupGP
cnbN4gee182fiHf1EeT8WidlAHNNEm9TfPt3Ir5zQhy3+NeAKGV+Kknf1ZuGaQxp+LSTEad86V1Y
FjcYUwI9OCl+9azdcF/On2NtqmgsLQ+dBpwFWViOR4fNuIJ6ePktvrDuMXJDOqKvKBANu3z0fLxJ
VoNISyHUmorp2uPz8MQMAgZvLXditTxq2VLu5PGWvNp4nZhi+oV4u3mlLwlTA7hAbk439v1OkHMz
UvZhTAR4Uqk8o4NvtBOj6AxMPq7D1iqDT4qxSz8G50/w3MT1WUva2miVP+NwuuaMmCtkjPK0T3yB
mdakl0B2hMP/V+3cnoTKB6ivmgkt4+SAk8NIF+eC7eP9y7bGVnwkcNtuUFjqy1+D1NEr7JTjjdUa
vQlZOsBcwEL3U+XjrrTtUcMc5xedbaOr5a10BZDNXWdO3q4403Vkl+FM6I2xHfhYf1MVpSLoxDyh
5Uw+kaZ7kCQmexJNVUoYsbRmHqHN1ie8QK/jE9tM9CfTvaZFxnx+RPv0ep04BhrW4r2fHP2GS0eg
/JJHZZkSY5zbjvsOI42kPPtgTBNJqlL1CK8jRD0r9eGVrq6sUJ6A+rh7GAaiRa594dmtZNjXFkp0
aH05xjWRT6TAe8XCpXmwmnpN8KpsZmdaF19EiJ6Odedkmn4B+wL7XmpFN5TTkuOWG7ybJU6Tsz7S
Dx2Y6mY2NlXep5OsEfPZQas1uftEL/YU+pHRxgmkLN64zIrOvSbiejqSZx/z6lsZbdSYIIs/cQtQ
S8nbsMvCoNq6zTFniW4aJsBUOXluBAHEqRNrs7r6FBGTjJtCExYQG+2bLT2gOo6SR4cefMkq46Gj
0VGc1qC23pWendR72eD+ekp1MGrxQ45Gxyi5NOc9VNK5aycWnCnqdRad74eZJe/+mKiHnlSWTu9k
eIjq0S6uUqCKwpJfADAoqK9EUM/cvXdB4AvYDv7MCmeLEIjzi+fKHxIAa3n8oc/8PUucZrwBuvBQ
aj2xMM9wFM2mPrHBQuXCDxPhZYw36TKgtwMXM1oMBJA118gu0y6PwM/QLQ8llBZqMrDLL22lpi62
EsdZcQ+LKFZMcwAeLHaRkq3cY22DTn7uIlJ0R1LXP4JfI41i0xmg8o2uYF6oiPfjndAWXSYpIS4Y
egRB83lvq9OpBB1qi9IuFLC97Q/CKT6Z8JJQ9bfgtf3K2GFmLWH1j8pX/Duxb2Zwqx1SDgVMI+UR
P/fCKgAxMgcvA1EH1L7UKLWTY+67Hq7OprsxcD5zD3u2ynmhEeEHrB35LHTNTwadUNNqBEF5rA//
ukmeVPF8pAXOUXfTzX+t1kf24eqI7aR0h+UUED6OTfrvgHI708FqdYcMWGQDvwRzllMmCr5zQks/
QiibLbcajWXJ6QPSpfbpPaBnyZywr36RANCyClz4+s2gjKBNutiNhjzS1Dw5E2o+qxqnapbjGuJV
WQTi4Yea45KLU7kVxMsSY5IFIp4PyVeqKz2d2qlolb27I2whvHAMbliWzAn53JxDoUP2G3FVwGY5
dAIbYERlrRqVtQ4CnyuxLI17lFFq/E7RInHpNAPnQoj1qzIts3wwuMEsb4ByhrFQD7inN5kyHvT7
empRXu56YtRLHet491MAwfsSo2y0aYxA/wxH3AnOuIEEPNJBIyVu0xmUzzOYm90rwnX5yOV49PiM
rlBP3KgavuUVE5ibkjce5rjIWkjAbiy4RxNlibqmE4xerMfsuYW/wOwBhacnsCk6qnoUjijpoEUX
XUwSmg9oBiDjmn7+sOLYJOiVYvGxh00eAoGfFqbLV9Y1Co9yBIulJ7Lzwb6mGZkoNMM0aINk9Rof
7RWqCJcN9PySIxWlJaJZt3Kt12fjeQkVMUPFXU7GT5HcxOcrE7Rlw3RM3Q0DGj/yfdMKj9bs20+g
l5HqhM65TQSzOMtM3N7K1HxBwftd1ToZ6ka7RoZXNIARjwkpsAvHIBaAk7qsROS41ZsObHyow8Tp
a13+QweU2yk5g7ZbFFJqOn+4YwCqNTKWUR1nt3sbG1l6W/QiamVNQMUlJQ8HsFaoWN6azTKgcv5w
rymbbGBY99WJT+9OHq5x6hUt/vkAALn+6QuL8coRNn1/Y63hNDIZV2ZaUZHMYimkYv8lsmNUFmJc
T43XJLDbIBPpAbk5YeRC6m32MGcz6dHpbZzS+Ab1aGQaaBsPYFhDKhh/93i35mMPk0Q9c1NcRqA0
9XD/QsWYAtPMl21FFamgpCy4aEl7gfIFw7Ggnnve1sJR+8a63xR5A1ar1CG+57FJH4IjVMr+Mtbi
sqUuZj2Jy7haloi00Bkg3ZbCW9PgBhJ/aeLCPQwWjlBE/UXmhmOZkh8KXdUwjHCz33Qhwqgvbw9S
IavexEl1MJTEpkWC9mervSLQQibEG1MxyqLC2SQldcJG5eYDKMUV+cBiKJnggj9hmZac63OoUPe9
OhpBP0e/mdvWuKe2kvvi5AVRoBA3SE3WBYidUVIucxJvBwU9AKLnyeOB+T+Qhovy8CfveKuRtsza
zySty6iBTHcvDCTiuf1ARy31XMriJq9narn2t9YpOjFwL2QiqDQYEytulArmAsccfXaoOsXoC04F
ehERwSsIgjfnoSzmx2Sp3bVaH8OdXjqMgM2QiEcLumznzI6LlfjUwEEplqc/1oawBfHA9dP/i3ez
GG5wLcM+Cy0hOWOSf872F/3dZvAf/n5jd0TIweUp0Xhg2/aXgYpJW9QqhIP6KY5xMZBoGnFKzfm3
K240csorl2JdUnX/t0+JHfIrgrY5GGkT6RloQbfAPT8lmP23pSmrpfzuOLPPFO68asQXOc0v5t16
wj3hc++dNjKrTLrUsiZxk2G2BeeSDIr1tY9/d3OjtAH4KZ8St8rpKCctEFvdY903ThVPa6zcsmYC
Rp8A8WWEgAdXuRKKZwy+P31gFwqx2audg1QhXqHKL3h9u4fgabKumygsu6dsHvckgyX2HuukGOIr
2uwvyIV8YRtG9UEd1iWnl9RGN6OJuL5LCaDEBHaaWPLio+qUsD10orudp3LILVaQxZgf5L0Sk3RR
hJXo8482CjTxNqJ660MTrsgXOgvIHp6aqxEvmc+oa053g/ehqLQiT1pK/N6cJzQ05R/rKNEWgPPs
FE6BMpqckZF3oy3xxaa49ugHxfUtvxlFteeihe3Yqy/we+EE0Qov0j0U6GPu2XCS5yO50+vGQOxl
9i4kh+qK1DgGvTNNcY0LU+BQlFBZasCw+MTtfBm7/ZYUxEAb9yJLBFeMrFbeLYAa+0T20t9CJAYm
w4r7gS2tYA6sd1CtiyCWLqLJVFnecIYFR7TAaaaHmydvHyCWO5NgmBLyRiTBMKKet2dZ16XBmaYP
cu4D76dOuoYd+MmXrYpp2iNbFiI7SLZKBacJX+4poPNX2W08QEbfKLjCq1P5r1G+XolppAqenRLG
qladmoJ524IFt7yRTtdVVBD5YwjqF5aQ65le1SOsbId5AfUnTFM5wpS+H034SVZw2XGnuZSoEp3J
5KNxs8363VaNNzcIzASkKWcTQz9HUDoWq9J9AyGNhNC6MWHe0Ran4VJlilyfWeDKVdrkKM/iHShM
epPyN4/pBrPE6ihs6GDGUVGA7+3JNvKb4vOdS36qyhza2JWZ7kU9kGsKl2ljAZEk8bOAZw2+lOfx
Upbhs61DDmOVSDL7pnDLfvyYp5qxWMh8TiBwDa7pkFjkCn3YqxDf254cQwMJ9uK/IUXQxHhem4K4
8YLNbhtOpt6/0D61wNpvOxD/Bzg1kjd30U7Czj1iwaeS0T630jHzSpU5Kw/tDZ/j5iiwllAT1Dab
kYIinahuDUHViqKKU1VIMgpJWDN2TyGl/N2mz9tNuKqQSSD5zC6MGw7ltVByig0a3l6lAIYW9Uiv
Mme0jsxyL/DMFwTEDRIYEVzeJwdXLyZpNJr8Iq8jKRFV2UD8GGIj92H0/o9nPsu3rG547etPTH1C
ckssvbCr7op8Ouxwwtkq+GuqV9O2Lxy+zOF8lXCKIpaEvWl2HXN7MGD0c1YwuG9UqKNmROdE9sZZ
RIMXhSMT+gB3BFYrPK/cydFd1UDBMQ4MjW560fRav7A2CG84MXNwiclOrWxTb0tKfCYekriHzxXf
rDyx8EMHVepuSAgYcgFtjUM7C0lgljgeAUGHDrHppcuzJk4uPIa9pJzCjlr40cqOIlQJudbq3Cup
muZ5uLRiWYrhSqm/bWy3qedwjVmhOEJP5JVsRuruYmSZ5kE/C9zR5rW9eUCi9qvd0JIdR+uEhw4J
U2GZods2bAexBWowQkRNz36mE8oOo6qdp4Ho3k9aiDwwShTBEGdmT/bWPlQdMdOyLKVYKpsW9WZY
M2jkQQRvgj3npAzvx8tFD6kZY6VMEReFu5ZnKToG92+by5wmt6xSkgayxayWIClUKM1ujlfJpbAI
MBfWy01t0bCt2kfNWLY2GUyJaz/o/NZ5GuwDM9ZlfI422GN5XUHvD9gjq+Ow1NipKNjChhrnetil
nLyr97/BJ22ETFZHuN3Ti6XWYoSnrG3g87+ZXs0xsWFH7yl+kQMlkDEa1pbaptfWPJ3QIuIP/XTQ
2ZNaM+tMlVIE3MUgp1zqI5aFSFxi5aIv4nwDy8NmPVKllyQRt1WPe24SsKMWk4+OtvVb4yc4BcrV
83oA+nzhKuXMC1tg25ZX0fB+miErHa9dbazosrOdFEjvL8Is+pySITMmAgYabAv7Rr5GSZ6pTo4v
M0h67fXyuL/gEy11MpskVcmdRWM7Pseu+QDX5VR0fpdwkFNlf5SK4CRE1lY/2yHn74LJH/lPMowi
+UPYI3oIEk7/ZLi5+3MwjRhe04GZo/J5gH5GiqmR2tNWYNvBvwXhYubT+o88mTN6HjemrehHl6y3
KZj/SxoUJOrgIoZn3RyRh06LRheExUC0V/VBwjrJHrfmgKAD0NxOLxF+JioEKrTNkmbFzSfQbM9/
ryUIJUmrynV3QVL77/5fB9vTvjbVHl2YPnRdFBxpbDDVEvYwbvrmHEForBweJKwMl1bGbK9pcr3y
hlj8o6aB/aCPb1LKDckHGIi5zv6JTlJYmETnCDXKaHZq4nTm2O04OX0/RmVtIb48RcrIyBB6rb99
nm/Hpz7Nx0JzisBhRzV0s07IkipGhRDHVBNV76urCP6PS770h9LrxMPUYuTyt+KUb0ZcdGipfE7m
2OYJs9zFGl3TkVMgx3rvu/7I80qCv+6kS7wV25jyuE21BbucXLxU0n+fowQEwaKSe/KTQoBuAwSs
r/uWGWtVj7SLfVwAR9XcSAiZsHWveWik7wpc/WGRGuJjlerbBo+cWu1fsLk1ytu40nvsrjDKPSpr
JY5S4ybIFqpyd6Ntnd6BLDl3PdcVdiS4TCLp8N1UYJaWNAvU1L6XM6+1KyU7g701aSoL68otJJo4
KLeX/wNktGOc9cMHx+u0//QT+b1iaOpGq3M5Ng51C46gNe3MJk04qu/ApYc54kYLoZgkV3azswJz
15+2reSRAkP8Y3I7dVRFJ9oP4Qrnp9AgrucRJdpYrXxNUTs716t9mwOKPkzNCG6V/hD3gJeCWpU3
p9oED3v1DpKKrhsT072M0VlDr1WT3f1Z40JU9A+NKSZ/qPKCAw4Ca74gtcfYlZFjM9RWHl9pTIi+
dCZ4itGY2f9//0fYHcbq33rshgsyy8I8H7UTuJ/YuYT/jSnCmUOuVVPiHjbOnzVkbPA3+pCJweei
C2x8YG9/6dIkYU+dOHhH5kDBlABwEVlkyN/NYwjn9PaYOvcr3oeGe6Ujhx1i/RmJjWBbAHBgfSSX
ys/paTgoL/td/91r2ilnYgsGaZS2aS3w6NbhmjfEoYTYm5njyEamL7ZZoiC4u8tA0UYPNKPJ+J2i
dnE6qbBdMlfsZQpR4MNiqE4yfm0UNmn4Cs8Ym3TRr5eTlFfbWRptO4Cd55+jOrqFjLBGYSWcpjAk
QLiEGSNR3g7J7vFacCRE2JH7CaSkM3nMqzWfg7R7a+D8Yp60wfwiRxHzCIf8vs6W4UwLaGs01YtV
ItqCsWIADTke8ELYh4eeTex6bITzWctiWCQR6+yYmuxKObWZdKaPhOmqu6EdBTu7a7AZEZzjLJ1N
StMlDsA9PSre7M+aTybwgFSEPj3NOYVuu9m5YBFw+b4NPgm4wd7HKSz60dQlbVrixJN2seUvCm06
Kv+cdQV3OUKCtuBFz7MMrhL42GCt9LF7mhibr0oGrbD2BjqxRfaoBpQWyR6sPDVeggQXRvMsZ+N0
yPwNQAOwVbXpSvIyFBx10WME2n1Bwy8FCrgZOMp9o7Ug9lZjXcxY1zc/Ml/65QDyevGJZGm5B2m/
EeMaWIy88ub89NgR9eWmOq3/mpFjzCWMYgub8cBrJaSemKvKc90RMrtbId1dkdpg7WKPNN3ezL6C
apltRTNNj4UWXsKwXU92w/3FINvpNVN8fh1zRwuTpfwyi9pXt1LoWYJwFKVZe6VF5bYjQF3fY2Z5
vOS6diZbX4a+h6uvCwKwvl2D/GSzffv2ESqZCInr0kE9ZmWiTnLT/XspBwSmZQVCP8OAmDZNPUCb
m5iRMbszudmjrCfI62+MH7kRNdRWVquBABL8Q+PBobgQx2pxjY8do2mUogBtRL9zN3IYE50DpnUb
an6vojl23gzcCr6k1lgCkUUJnDU3DGKIzvX4+STwh33dTby5ocq+t8YUxONeB6AJvIYqkiqcwoIn
8+4w2NF/3bFAUM6FAmbvQj1yGYxsr8tBY7n9pdp+G7cp3zfVnLo07muoC1NlczLynt/yr4UUuk+Z
95lIydKnoqKGN9lBH/r78yKVAheehbCh02k1vmcNP8kK0H67vp79FJwj697/xYAYpv9kJLE7y5sh
xyJcXFITlbs0IXsDQohMfOgAKVj/mm7wIuJn0AMHn5pxGzJaHwTdVOvCwi2Ergitbf6Ry/id6c1N
6bjVzoO8t0DP+L7i9nnIYqbvv0sttf0GMRpiF5yG7BWmGsGhhwrR4QPWUuYLP0ZMAIZp3eBdYs7S
wDCCuHW+APtrnsWu+u/aK7A98nT7pyt44QqBtdwhaJthHP+JWazH2c1hwmLgoaqP2k8xvrWDAZ66
PvTx2W+fkkpT/+FYKL4Fo7Um4aLToSjVcMG+UFylFkEKmLt/4nJ5bQbu6r0CRaQjfajD08wiXMi/
pk2t6IrqubCCJ1StwezdPkHHPd2REFXpAG9DBA99OUvwM8UEqkuIGmXcFolciccMOruX9MfjwSJi
eMgqh1jIp8sorcyfjjSGJ74kx4idhjguri6kTeOFi/7afiqyTuoQkVQSfSLxTdz2bJLFnmbZpiEa
bD6Ms4d3/NeSAcL4AId8l2GcYBjebA08xt7lx5xY0VIwCrQGTr0D0PME+kpfEydQRsbJWnj0OwlZ
k53wTgnkhCxxEd54oKePWxIry+9i9MCh/hSOImOswnENpQcHGTZ/miOf0dtY8ZJFPsWwaF7F4fYw
fmv68Mq9fsbVeZxv9ntSeZ9kJtGVRJohrxwKZ3dZLz2FDLJXYFJ7PPg6J5v7uIKw1IyLLjz2Rfhl
UCTliLRyX3CL5yyejKvqqwRNMnJpLGo9ryUMM5O7nczzQsOC+V6wuLjTNWTaFXJRRFsDATmrgo5F
zD2bjSzTqGissAc/ChG6IyChrg+H9jug45CNWPuaAmEJBkuLsBz8PnFVRdmOt7txSKD+xATuQ63m
OlAukbQY7cSaY1UhKXSF6LyOy7EchSnaLXnuDXE82AwpVgoesPjU983/Fge73HocLws5Ms6qjnaE
zDz7pEny5aTL32F2bchOJW7sI7K0/HGQcL+YpEeV8HJkMHbVPhpO3x0GH4sG5wOxurNe58UXYHPL
BOEcBrv++jLCitlyZVHOEjLoYxiJpx23lVJAqeCfLOmax9DCVIvvMCGiGZTfjrnbZ3bYMHWRAFxy
NEGGri62NcYn9/6rvS+nelpYTj85ckNzpR7eStyYG0ZJgehNec0EBfzGKSrhRqkJxSPTLB8xy1MH
ZfzcdzNRJyX3Ztk8ym4bO6wjgfwgy3t+PNIzwEffRUZ1/iLMSF74XCXK2OTj5PJbbShOJ2krw3jU
QjuNU4/+xmAOgOO+Hj2GBBxqLXBxqXj6ldd2cZ2AZO2Xs2r4kOzhDviKO5Tt+s26yzLjBz38+heT
Vyy2Ux8ZJOKoJkUt/aK5H36slOshthNtLmwEaLm3e8W2T+RCZ8PTvPh+2kqJmQU9T9UVsZqV+V3C
juojpukEdd99mXIHn5K392LaXWjgYxyqgoKCaFllsk5//Nu4FNfHJha3eiSWblNvCxojge+h7qPx
zUTtj5Tlo+BOR8oNXZWOEmq4hkXrHjwQxtdxH4PRkm1Jt7zNWu/YNWEa02en8omlTk1zufMaDglA
KoV4rF2P1hRWwLnKFU+Cn+ETp+F4GC+U+84S4O0YZ3mZ7x30txHuBKCe91rj34NLjGF5HWFunWw0
0Ad7REWZyISz/LTApqz1D7RbO0RoQQKeasfgRBPaU2ECQ7y7OBnD0/sBIN4JF4AJGagkK/H9HXvE
Iq9aQvyHT9V6GziAXpeeIFwWbTW6l8m7ZnLL7X7KaxJyImG/JWAVm/id8f1Jtle5Y/og3FXqAaCB
/XWBnBXAlefCNoOc74mt779WnCVZDubLVsNquTB+Chkalt82S9LsZHa2wkA2srnkHVqol0b5pJYd
6MpKFbsDw/iH7VDfcVe1rPrH2S6eIDDkVJypkbYFK2rgvMpydae8wJKWox0vVgV1K/qOk3pr4mGY
5BGdHonQnhsMg00CahgB6rjEII3Qdw5wF2qCg4YSUM9Ih3SX8aw0u1f5OJODMDiX07sLw+/bKfV3
KOzIjcj3gwtOg8G3+50N0GkitxW7V09w6iGUUze7QXXyxg1Xu9qO49r0px+zlnKj5V/0/ugllqCo
yywGQZFEPHsDgy9kSS7+OyssphdYMDsxkVnbm1YQVf0hebK8K4qyTxNINkucHz7YYBbCD8YapMfU
DBXNDdwboW/RFbIwzQKOnXyk81q3cTi0HEbKwplspPQ//uuHDt6KDpbmdYI2btArEXgCU5JF4lEz
BrCoUUQv+0QM/G86GTSu/3RQ4lpciJsdTj8lXeTFkQZbGVgVTyj04Glc8kE9NPY94AdcIRTT8wlM
/H5VfV73qiKXzBNarW4oU7MKgxlKLWcqgnt0++nu9oljbVoh1LfY7ILYnuc7Nryc7C2r/PhslHEY
fE2OT3tJtKRS/+hADKqMxkwe4WqY000lDf8dGH+VyGVV9Q52QdBJGo7p0KW3TxPT0qYz9natljnm
fq0+xXsjf+n35wMItiKUpp81Yb8xEiUshDcokbBOL0OYpB6s7ui1kU09W+5yFPbBOs6BABL+eRek
1GdBaMrex+Z/1fln3u2+cHhSenVCvEt53eVR3aCDr8zmb6BPd8Z99BSAhBllc75fPAtFf2EFDM5B
8VVmn97kbaM+4qC6eZ1SJ5s6MJuMNioDrecoi0EJhbIEsQP1tZkPklpgBTZv/i0GgKnC/cGQZUN9
JvEvPmtva4i+cpLwv96gLasgNTG6INqIqdsbS7sOkxzNLImPSRMppKYJNK8OPylC8tmErKt5fvjh
oDcl7FrY4k/zBsOxE6xV9pob+VqbOg3w21SiE5U43SD9QKlxNip+Y0i8UUYku2w4i7gj3PD1Izj3
+NoY8bTyiTGKfuV5lXFNMtvU6+IgSfSmCoRsjywK/2V7A/tH4riI/LY3VZ3t/mLBNSbNEd6g6ATo
iBa/J0B7nF+D/w0cz3g/sq02fwlXCcQeYbygbmV5V5iypHv+7nGHGXEOePZCxCs2DsgUfs7F8fBp
+fHUfBv2SmpRmIQtqp+Tp7WEhJkzwh02EyhUUZlSU0LlHvTCpZq+UiLWxpXbous2mKzPDnHttf3r
nPiFlJUmFiiMzSdsoJ+jfwfhk1cULh21lrdCSDhE5IBpgIZdn9eF4dQhkAukKQoIa7GtLueZ4XFt
gKNGDCiNxxoS84tWsd+Z44LGqzCD+pkXpx2qQhlI4j/wDaYJr7QR0TGGY6jbQZ7pc/JJD7IJdjRw
SxEGocgXeuiyJKZLaFfmIzNSG8qj6n3C3iZYnelaoomInhY2eHnydTVdrIV7DK6eedRfzGHCO7iH
nC2YkZzwij4WPQXsG3nLhBnFywB0g9be8brKAa7weSsPaBp1IR9Q/ViUddNXr6bbKbEGYiYRv9C9
wwf4MAl3ORXBNTPGJIQKW+qW8VgTiC8g3508vGQVMSYTtPlxhHhqx5U6b0wcsHFApicxiYwHNPm0
OhLrzngMmz8F4/o1vZ53RVDD17wSZYazbeBJi4Y8aM2DwYMk2c2FahaY1jRmkETE4VSOj3VzTUk/
ayZMoFcakfyaMoLR4JPe+Fmen+4+s7BbwvJLTBS6HZEilQFxUAPH6XdVgA1pJO5zG4ZtNvgk7QHN
n8jn3vnLgOyN85XoDYNnrPBurxRdm0dBPm+CW4CJUiV5znPkkm5d9JNQ5NcaLmmTZ1/Giug2fowC
ELwsy9tFtDBOLrRBBezUH8GAEzBfwFlivHisK1e32Wt+kIw57cQ1jEVD4rUABbaZLUBTCs0IjmiL
lS/pcZeDA9fo00wCSpWGBWwsrX6QCpnJF6I/SgPaUopw2ciFnCzmrU+XsT1bVV0hoIsjB0thw+Yi
RyjVSiwM5tTSgCUpBjNI3ja0PL/+tQeL64meIfZJEOGbgqymAefIvJWbSq47m5PoRZumkYhTgk/P
6SHubse6MAGIyZNo2h1NshTh5yy0R6AKa6WYBhEcQaYo0cC5OpkLWoMHOuEtJ7PiDfWKUdO5Lr4n
g/HtAsUPUtx6Gni8zfXjR3HI88rpXVpYzsx9ZulNWUHvgBZzEu9rxPeypvW94YRVE1WUGZYiiIbX
1xQySqPKQ6Q3b3Amwpxa/2lLfmioewAHR4qU1EGO1ibrUYILQZt/S+PReP/mDptOGBuncVl4fwGO
bZp2V4vimUy28W/cNCSR52lbJi7i+jwq35SRBRvslLnRiQxU4MfdPzsIEEMnCMTJWLiNETU7E/+g
mYP+RE2HGLFuA6YAs1UCvRXJv01ceu3ctnp1eVEVv0oxPsgvgGu7Df5W/gn1Hy12sqfe0VhBQp6S
wkVRekoE4xd1IFfspWtrCe+bO7B3rmJRFr1GvySAM8et84mzLJ/wFqQ0OUuSANl0hB3gjpxj5CJd
Qw7TbYKK8UsGX3saeBzVjFkwWGUfbuNayszYrew3YP1sdhjsBc6LjQxKbb7z5aICdehJlSdD2fQL
X7plUy9yY5G3whAuibIBgc/htgCHS+YzS/3d2yHbM3E86a0b7uqpnF9vErEFnk19/AygzJBk3aj+
p5WsaWaMo5Myn2j2vRIqelnPgOdT5ZizKSkqrARod4+2squQwckH7BvSQ9ITV1kjH77xPiyiF6fw
V1kReMfTVr4Dfg5JreRA9+F9wHdG
`pragma protect end_protected
