`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3152)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpIYXv3IgOlkpdqxtXZtNfdu7BxMAIHPBQnwK4Qf3rMs+ej13W7HpIHk1a
nobmPKBv27xnDBfx6tR+BLO9eWr4d5yFAZLdvziWyuq9lQP/JEJgLZtwmpaeEJmiyTSwhBjJ1IBz
y3BtZayzFWUmSkWng01uM1+dANNU1liO3yKm8y10MraUKAstawAZue13x+YmrLaLF5GWhNzak0Z7
2o8YbGgYDZQVIJ/5hwR5zRo2mABLicp+3SeTfYpcuhh/41ObXVFbtM3yhvrjPABUPUpOgF4/IR4w
W/6MjoNQUqpMsEM0SoC05w9YmrJlpOPb1a4Xdy/jp2qx6sKKUKCYvR9+3HtUMErMf9qNFc6oSk+7
t+HDv77rFU84GudNoJ179/5iK9JheMlHYAB2n+TxAw+hSczXeO6dGz/A4pfFasMtT+TAFrBtcfoO
DUyRjGh7WMc3n6oGdH4bIA7yYnSToht0oWu7qHCkocEF59/Js/s9Jj4vqeqCIQZv2COUac1ad1Fu
rzOCgDHO+HNmUyt4UbUZphMQZsUhzCTFkNEz3fA0T1JMlqLUUitJ7bpGuGGcWNyanDbsi5HjzEuj
bZviAUiYVfxkFm8cWiMiB3+RhTmAeRsuAOK46D7gYdA9oYzqIwD6oNq3a7YgmS9gjqus5lV7qFya
0bsoeO20FFM9q0+So9RdSH2y5QucAboNwmR7qLEVPhzmGvx+D/YcTG7hDBSRCPMUhHO49I0QEEdw
IMVPF+Qj9NS1wT9dftO0kdOmyxucnWaj45I67kn7MB4pg/iKvImVaK7nANpQjc4nnJQ7+kTLE0EB
daAjlaZkt86EptWklmFAUEIqVceReKFZYnPYMPnzunyMdRtReniZvCeW1pOLqKpasGQOd4b2ZUyf
0045KPIlAnKMUxSaUb3cZSAiInQ8l+oks8o7JhcLBQs9WXsnMnWUKJewMbc6zn6sd3DIQ7EXO7XK
AbLdP9/M8cYc9vPbzpOcorGYk49NBc4url7Ooodb5OfIYnjXoyQcBcpGKalzSiBD09Csr2djHE8A
I0rtsWchTAXwMsUeB8BlhWGgENnfmvgPUCaYYCajsDUMolbG8WNx1i9jr36Q9JfaHtH/m5lvxoIF
4bs/esHx6+1I81nb5+tRXDGCUh9nz2E73mc+ptKRucqKlpYNCBbAsN6aRnkMU4uoh38Sap2ONZw3
YAFoV+VwvhS1gsyNEgT13UKwCMfJEyuyrPxq+CvL7VIqnHU3XqhgtTq6BHGcy3esEnkBtPKsMey9
g4KRPl3Zsui6BpnsA5BoIF+mE5hJRo0AMuW/WYstTHtDGuDCNG3z78eI3aq7ZFMkqIuALJNpo3wm
iQds+9HQRhcOrxKAQKjv0oRmGu0rvMcX0ux6yWJmAG4PpMEdt/BdA8EhDn0Fd5bwnI13yXFcwYUx
lwzE6EPFOeMYz3Auif6iJT1nHUf7dc+9T286nBnwegm0abvSxRBE2HhInb/awX8nHXWW7P4vwCkD
G+v3GpbEA+rfSG4Vo40edyukHcjTIolO4tRM1HxIZrN1wlfb4fdcalA0ON5Zvcu746DLwdK2c0zK
lO9028IJHjudhWz7Ssytt395DpBDVVOj2omicwQPyeOIRsmT7nrIEDwIEzlQjoLie6PRxFC6TMWA
naS86mP34tH+5+O4wr+6mNugZB86tS3ASBi+9klAxqCe9+FejjqV7jNQQZxKIC6SbOGY+x+ggEpi
H2i+nneZdKcQmE+j073sFTGjzTwVsa8v2Jfmcmx7F3ievb9T7wvdhk2IWcr6aXpJZZ3Io26GQ8Lp
LSzmBl2uoX4blSeW1Gp6ko0tjW4xqq87o82HgSyFXOdb4y8oYY/aMtG0IuMo8l8IO6PwY0w+sO46
gLi0vNklLGpYRYIXmH15mxk6P1PMY0BkRTXPTF79zhrF0Fx67PADOjObj4Y2mHn0MJvnwgxU1Gxv
snX1IvQdFImH3bEwJaS0MqW9I5Z/MVppDnJgJFzgnVkK5HYNUaTytB+llIUDImn62ENVZFhA0De4
IliBf7ETK/yp51whefYa3/bNencm7Q3Ovgajqr3sunsDlh0jxBKRZtIA4Mfxoch1sZqKU/u6q1Ct
1DEilfA2dgaJIGnUcDVSQsu+c0JK1vD5W5vTXTKvVug9uBowpX5ns55L2ywiDqzrelW0sgvfPySV
A/M6JqUMidi5R8XoWVOcBfj4hWQFUHkaaMShj8BeSg0J6pfGci6RNS6h18RUE68JjlNKnaxytbPw
E7W7mW2lxbYOaE9J9Xjk1xTykg20xz0ZspLn/I/ovNU1hDEHKqJ3DTFRvTQVgHeJy902rn5iLDxY
dNvBTuZZElfzkEDXaJ6pjk2dUg/0s6MOCZK+rFVYgL+udBw1A7oXrWQyRTE3JwXZaiPT9YzpYEHO
MiOtZArGdjMGYMgWOa0BIhTCG+BpXpEFEI3MiChoU4knUlDN+vqn0SIu4ACYxw2zhnZWIcmTN+8E
DobOyg3fMSScrQFrrwkNZSvA5WVI92mEoUZqxYYvdO7PvNJP4chmzDCQf+5sVcg7MMnE/preC/hs
FUtkszE64y73zCW1vxgcKQbeD0O6gE3YD1geMBeyCsONZI7Ka70qoS/0ef2zEbtPrGLlyM/npnow
PaKk5joiKVZz4Yybh5TZsucvsvAl2KH8UWeXfdaIA17m2kkQndenGTwTDeo41SMxRCrbVrbxfReP
xwd99y5MkkvUBCvLS4scQbifIMvH+5oEawsawzzAHgIu5NAvItIK9FBOyd9OQWmJpvSg00R/4FXq
8/DiKNxfpO9rHFZLd+GxN61GmV4RX0VH5cS8lo7nWIA4KvC20XoXkF3HNMh96WNR+ndHOzd8jcj5
V7dJ+5afx9cHk8zgpkriMZoXNjmTQgOf2DawNNjIEPsX/BIqY59+ItT0Q3BI89FbnU34NNiviRt+
ASdHLXG2xBsJhWrpX4OHcrAYPYDFCVr3htmpzGw6Vgf69CQWmaCUSvQZmj3Sn6UAwvJ7J2lnn5YG
OpPLzLhVtdtGrjAOyJQkPdX+Qg87EXKihgpNX433ub9nYmt36dE/P2W9mnOFC5vKaLWIIxkzP8Bb
02aTmY/N+kxM4I491BcSE0w4XuvaodE0NUc6IdM321QKh5F8YRC9/qw465X5R0pGqiU9dcBPSr/p
+AvVTQcgIOP95Ihdsa3ybnlV9/MvYpEtRRtn6X0rZVbnhC6pS3TCXIgXHG1M5k5wFcmcf2aHWWNg
ByW1jhONhs7RwN+PQ+LSGPpTj+ctUZtImRt7vuzvi9hiYvkXy6UqzmLud/vSkJyUAEjcmqiYpQJx
PRXDj8ex9WejF6YWtTj5a6KF0+cGSmleqWIEu0kwOH8yOGZh9Yik29JELe0cNvgMzsW3vrJF6Xkk
ztDaEzQvT31iu1VkBx0nTGPm9GY94SCTlHqAh5/eMc4YW8XxoFB2mCm2UXY4uW9MyKjVDG0k5qOm
Ni8oxu8OLnS/LeSoi6A+eh28+ohyu4+cW11YCUgVi8WyS5g7tYAaBnLxb4eOImsagocwHeJEGwp7
U8UENd3VEV7CLrdSyjgn7kcvEwH3d2MHvj0iyrr/8tjOj0gMp3NJHWcXxS9Askz34gY+p5K3zk7d
/8n2GfeW5h1Lz690HTie1mY5nF9cxxpGPo1/yOgCg75uUBJsyp/jge5zjgkDI8b6wQuMrxe6A2lF
14MlcyCYvAqSMzOlXhAuqLl6Jr71Dcm5Pbfkb60SoRvgIX2vgAYfm2rtZkQt2XLR/FN7XWD30+/w
/F49sl1JWkVZ1uHnhliSSn97n2CJTyiGZyJqv8q8LqWIWi1e/9fgjhZ1KZFHIjrN5NS0M4ZNKBEg
o/a3ws9ik+d7ilHhkdh8pWd7KFGH5r7ZCU0Dpr3Fs2/rHq8ZH4zHjqCOJY/ZUDnNFCJKCibi7J6+
ZoLqcIijaM3ooDj4FBwhfJ0a0UaQ126UqrH/J6f/88eCD3nY/oP74vv9w/zEt3gxkNpYcY5OlsZP
8QfQ5QHN1dYeMWYN3Cv9EVReSSZI3ObiYDU2lP7aiO7PKnPNX4FIJhII/rvzR0JPC32lT9PfksfV
R2FJm94yXhQtWuQYd9fl90BVyrGaimdxnf4UVIpI86wLh27TzgVPHmFz7wtHppo2FA6ifrGqbRgC
vPT157WRkAgIGi30/6UMUAo=
`pragma protect end_protected
