`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 236256)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpIWLdwh1N741cYz0y65ovQWOvQS+HQxb+48fKT+jdFrMW6TJVez9S+loA
XfaAcxQ1NIOUrANwc4BJr6ZN6v7LcwxYnA7R7cBY3z1HUplqfBBoYSnIwtIvTfT90LkK9u1cmZ0O
LMAo4ApYNNdPj4YflVewbsleJ5BTx+hQaxchHvJPbbXihByyP3+l8GfhFfqagh5d7WRnOT1LO/pL
z/rqWxXsa0MrtvYV61tT/Oq5NFpEX9wXeqN9T/PYy+ml3oyQQuWdxBd/oWkK2YBUf07AVkxIbVZc
ISkyOj0+gTkxRZnJpkd+uRxFC/XKsW1sufPv+1QLSw6y34bMLYMIqEAhD9XRbz45iHQVsdoW4xU8
yF3H5Q6sHYJdwOC84AC518muMJvonfgJEmR9wXY+ebHH2PzY7Rc5BUnMH6RRlXE2tNyDBlgT6Gs+
PawHS7PVxykA84n4hoisNxvGrEsfO2KxN+s34r1eMd+PKm5zJ8sL6aPgENwI1Z43eafgI5+qIWb1
YvccwXoM6+FiuiI6UP1DW1YVykOnl0fccpPOi6rUYMxJcr6VdSMPnpxyMYEq3OvG9NOPHD13Ke/g
jS/p4GxNlS425RgCZ4aaJnRCxxbLh+1hJ/Mkqi1gwxxYlR5TszL56erB5hp7GH7ar7lUE4vLn+mj
iUXrEPef55FSxu/eJW8JRymaAZUGAYVecvUnSOsSz3isDIasPstZfoJRKtICiUM7VabzWL7a7LGW
+2B5aeXW+UXexLvg71OsKhfXkKcwhqdeCjbG4iRCB0U3rP0InLkaCjCWnHudntTySjheiZ7vTqz4
XuC7OKVHRf9L3pojaPvORqq3Paph/1CbUiPl5Nc3KHkYvQ/C6fWoAoX6wpiDxGV6WoX9KRO6De4/
j1vUONpkH2hOhuh44Jnd0R1GYTq7huafWpJzeu8TP9Z0pdhinTjpBY5HB4uKNrBBCMAKaErMMV4J
PI2w3rxa87+9PjOWi1nEKgG+Y0kn3AemmrfyYde44grsW4pnNPG3+ooV0vZquikGB64yF3WqdUhK
x5FX5OJUGveZ3bFVxIsgSxtnXQaq3pCuHhect+RKF1gpHpm7bWXiiv3q03fGsOuQNyGLJWPYpTok
sfcDc7Ndge526F6ZuiFB1vF//DbRoVYtj4HMMRia60iqgKuy5Z85hZ/am1g8ktAGJ4Kuh9AAa03V
tGYWvSbg+6Jc0It/VE0yGiZfDJ27ff+/YCLlTf/thVqIWgUamhIV+521pi8BcYxwY+FTBAtRTiF8
4HlmPL9o44Pq99EkoGJVjyW8+sHoQmexFKlcjZB4fHqpe4QMufBsupZJok9sWE4qqrAw9gpndzP4
RcyYDvpSrc3EzZhV7U+jEmjqoW2Le1a65oskT9Koj1Lj2LDlF39NmMoQpKPmJFOfysQ6hnXA40e9
aw8an+PnSBX7OPUnBRySgrIQlI2r/ZIi1PiQRj5lht9kPm3NQkc/EBn6FI9E14/kWKV6t/u4RxdR
rWDslBbBiMb2tsQefsO4DVmP6Mxd2FUdi2+tIyHbL1wsX/2mmLb/+wwT/lg1tns5huuB3l4B9coE
IWV83UiPCfw4abj7oAOPbj/qlG8lsOaI9DCzUgCiSXum1rkbWQbUYW7thvsQ/sBxe1OeCYXqjIXG
mDpLcxfI50gVgCw5CNrTZWN8IgcFbeSfZP5WG6rVMKMMzHnLCSiVJQ9MUowJIRgXQrxPtPsb7CNT
3ySpCI+dyXWs3XnLeU/EZXTnLJDKqZxhSs0x1tOV2/Rpn33dKnorjYdAdVHitzTSgRqayieWMxqB
QiZzxPtYaHqbec6zGF1cMviRrycAMhwT5K3adCJGWBqReq1H12gsk+JqnVhrnGK3G6VLReg5m0Zi
cvCsZlMqcVacCMZo5dHYdK5Y1vRRiVEJlCOxx8lsIAVr+W070X0iplGDAP/vuSraYWw5Q/n0QJZC
eancXTbhlPUsWU2wa6t5gn2E4HGZIetRGTlmaZ2UFBLcbcDGOrKO4vRE5JVCxeD1rQUCfIvX/oIi
ruq48z6S/Ux5CjoBlItf6Wt6hPK87+ibBbqipRUNI81gL184pnDvwuPlsjEAiWlhwFTriwsGlfJn
fJGxu6XwRK5mL7tu4DWgyf0aDt9htXMIAHKcLI1xWKqt1Tg/Do2/BglWG8mChFbMkylksfKc3TVF
OaMP9uQVc2IXXYD72LcyXDgvpRnboo4+7zcMMMf1BcUJgV+MIFblCMahe+JCKygbuDo/3ZMuLJxw
OOZxYd9NLfSU+v5KRh3C1462O0oaJFaNhZ+si55Gn/6r9q9H0yuuMk5Ph/n/TitemvhZdID00RRQ
RjS4b3+1PjJGTrF0XcmzfPsNItuK5DSzCXU3ecS8lV8FKggV4BP7MCrz0dv99Gv+GdDZeYhz1Xxb
HyUoMKFBp4qjugHUbAUUIQttl9LV9XLp8T3fx/SHlzjD+utcjVn+16T8vMwMzfgkwtlZsbWOCw+s
4Zb541sm0rX1v55vna/1tenL8jQBlPnxXCzNPf30X3HoCn0rvRIfsQjl6iQmPljAsJ09AFcVZmtx
a6vZJ0YKCil0cBcrYp/CbdrEFPxnr5P02ZTxgSyWq729jMQsGdWPMsn3B9OsDL8W4cuQD4ETOKQL
MZKCOPDnaxbtkkDkjZ6Ngs2Z52N74EDexqYc3EpM/SHHyWUJ+/uCt8OrDJpVf2zSXcDLUvkmTvLQ
xKQNcsjjPn6lC1KwKVB3/ncEJ0ovHHG65UvB/WNzSJR5MJcEYq7r0scUer9uQzsqgWFqH/WalqKM
tk1YHmWu8u+LcGO07Rg4MImot/np3rbncI66c4OIfPwvpYxWs6uh0q1nm9A3SUx4zNjlLNlLGGab
PcitqEH4BJ37mciFaWCqWaSjobD6dR0mMovj8tI8A/A1/1WSXMsjN90K6M9w8AUwKXq0OM9G3NnA
qt+QOO5gXkH8qtKmflQBMSIZhHH04ytq0B/8CH0g595J31fR406MZU8G3IuRkUSloggx9qBztBkf
5lb8rPBVr5BanIRgwmWD1avcsmszFrB9l4oJSBBcYroPw8OO8Tfx9UM8fC1htabqmDcXE1hOeYml
hJP6ykvxPlNvqiIYi0jEZXI8dQseiILSluEkhEXWPhXSliyf5apOtmLGo/DxrA3I3N94eDBV4FAr
+XhVZMJ/hnLH/QKpc2LmiICntquRA2EoKuT2fGWrNBG46hvsWSNM1cTPFXj9zApHZ48xQHM3MG6e
q40zvFeHsEtAdnuecfOlpTDUBV37dI06Q28iMP9YBUFIb2wHRRAj9mAKbbbNncQ41TET3uG27593
jdgqcH/v9RsZtI7fKlZdShMOXDpMhT0a8oMc2IJyfLkbbbHDH1NqXW703ZDXAn6ukdHAaIs+P0Xl
0J96VbTzlNGrcjp2HBufh9AU9BIMjMSQyQGvKfX7ggI1SKu8Xkkcgu8Ln0JVQsqidHt89ptqy2vK
RBCf93DPFXwAeGDw0tnaMj7CPIggJVZ0qrcrptnVlE6/+s38E3SdJLIqkp8IKxsvKcPLA5jDiBrQ
VcLxAYGLSSMPMqlFIIZKNyRPdXXrWxavQjqMwm/Tn4/KrGymKG6EL2wgociQmtZwrNExyVJipVJp
m4qKIP/VdV3VJup6RPF51g/wp1b1VKUfcZznfPZwBHE6paE2prFwXXl66ExS47ZG5raIdtE6d1Xa
Si8HmTvSC9qKqJ0R7imUOwz/XStfzThJdJhBUifEeZxmWlY7vnepM2dMZSKIM9I6jGfchErI+hKn
FUHtUkog0fkeQaKIT6JbJEWTQwjiyqlUMSvz+Fgx2rrHhiclLqlrs7GQkZk7iNDt9t+BU+ukILw8
EzkD55BuPEm9OTCXCMJQ5YEap0U4vxBDhR7EgOtsPsh08zZlgOX9D6vNb93ewZyfNEc8r2lf3hJg
JFw80qYd2OutICNPXrYRwlTWbn6cLHW36hXWcWfz9Iy2vGSEaLa+wYkGRCPJ0jWVKJr1JckRM4YZ
8sl0GZViEIFDr/CIafrQLG7v5mLhk5Vebj68sSZvnhZcn3zhVnlmR+Rdf3beJ09iIVG6ibY7vw+q
NPQqBadATUVRhU0pFU1M4RzJXWmrtUxJvs2R6sfZg4MTdVza1thirhe4yJprZ0ISY7ars8PsVQ0y
KpjZr0DHzspfx/p8rznnQP2q8CiNMuJyBd4rVOYmAU5KN0b+zKgKqHjIWsvip2QLV/jEavAifkBU
KBn1YohxCQVTRijqPCYWLxygi+iTxpSsOeVHOVgW42tA0ipxppAdv3m3WTFws4wmhMH1DIveKa4U
1CatwC5SdBXI2ULFgM7dkRlmLBcCZTcai3siUgTquoZ1pYeUotnIMoIEPR8fbmO+6VMUPGpyLzvK
WEcXHapyZ50R/e4ACIIfiPFeiD6SnCb7m8NcpvfSyD3A2XWPpVcXXP7hVHfKu79ag3BIJbgxRL57
TgASe0UYic23fq1ymzF0An4PkCeUq5XjAH47DmG094CwOD4LwY9O3fu8FKx4jPccqqCQrtnm2G0p
s5yA3xcT7WYfPaCE8AIcnQ0JRbB1O8t5e8Cy38xopj04F4Li0HdRs7JzRPIHttZz515grfODzGSX
WI7j1tHqP+aTPNnMT7yZNZsrfTm+BwMoUuLCub2k0nCWGVChCksfNFR52BrjEUAx+wYfGD4necyu
W4DCjByRtBRwQFsxl1pkYFCCAYex9Nh9GytMY3YW3MoRfiY7WFfEqA/qfrHL0bBoL/Knnjj9hf+h
mkEgAS506e6dIo39hTCx1JIkjMiVqepAiokJIuY0agAcuHqyjNw4kEr49sqnFsfDQ5YPXqHuzvIY
c6p408D7mujvSaGWDha5gF+JdNKj+aps4DW6UudiSPwq4K0L7DYGhiQoJJJMYrH/tqaa6BrLPDj8
DsF4w5MppSByKrnifERyShurl9hUG3fgUplqXcCcZVv0GLp2/Ze1Q1qaq9Y3P1XhJXyaDuEjgFUk
yEVQN2dfMUjiXdpc+qVfeazroe/7V/dswIIiTOhK4cB82bMXo7A6sP6Yl5dF/5kiODdDLVig2HnG
o0InLkzl+bT7DvRupS3ObxWfPGCzAQ+b3cdHse+xx8XHQe+z3Ed9wjbCPCo1pQyNWXdHAPwCLKi2
St7TGExxV2oLzZE3g8h7meTP2LLd9ORl9hf9S8f7DoTxzy0O3egxfyMLpW9l4420U2E3VWsNl/Wc
lEhtk3G1/SWeZMeO8bGrKb76vCB/eBGpeYOVKYyaZB/9Gv3+uwSif6Yy4oFYlfoU/783B24UVKnd
Xow3uok/BcjwN1apZk9VkdMV3gLh3Shy1LWswB1t0YQPFIcqJ9tjBXyfjd9nO6HGwWGhQP9VGK8M
ARKBDX1X0A2guvRr7H/c05VKeFYjK91kXjkMnNYqc4kFcj4kLPvOBODYvVWN5rW1AFAlCwZax1cR
Jb5mTTh3rExBIlrowlOn9E7eDfYVchOWh/AZ04JW/FElzgpBo2VHYTSIIAQeIMyT5xiFxpNqUgvd
W7fU39+Xhfgg2so2dHIm/nmiZfZCDpiuGj0Q2+vu6l8+FHkIPcNBx2n9DHFYPd5RhaMhtJwA4B6q
93xwfQZEyU8nZJT3PAkY8snSK28QMmEY4wMAOblg1OnHdEweCvFHC4kbL5EXo1cnje4vNHn0ylp+
nP2Hglef0FUUF3JEaisw8zKPQ/zrmabGV9Dq/H2vHxjr7kcS3Qw/gS2nxJ1UlcLvun2nv6XQOjtb
z13ZurZFzEJPfviHbSxqwwxllLNLO8AKGP6Cz35q/3rOpCrjE0NRSRmAh8IQ5SA7/mL9kThrrTKi
6MJ1DZLk0Cl4bgxOtH/hx4xKRyd7HTHBM6S6qv8sGUjpRzgcvWSgFIKAQ9kQTarq+U+R5QDIyiBv
P1inF671OooVTIam8FcVr3to18epKCaiO/lAMiXq9ydCzDSmr3y4gP4QUsS4bHesQgC535zl0IQX
BVc/kRIS7dI2NHnPdIxlNGPCjf7qKiDISmwEQJBpIjoBAbU9W+Tx5QZculhzQzIBSla1KYGljjBS
jfFzYrXlS143a/gbXuXmKx/Ce/zEZmJ3movPkNsn9ZdBfFcoviUwAkiPxsO+jp2/0A6J7JvXSjs3
p+TMFjKqjXiKy+Juqpje+skBPpkwGt0P1gDUN4YcykBeNb7MRhaAoiyjK6gEa2XSDf+m77ppm9I5
Y1lg9S2xLrCk8hlVtZ01CKo5G78Xam7LVE0p0eiu5vCJuDsjQukm/UkI09ZEAF0Nyo/S1t8aI1b4
2OVsHCVWYOCY7PoOhyIn1I0ocFDPeljqTB0q3LdYBbqSag9EzEBbQWVAIifde9p2kVDBnat2ZGJp
fkNfSCYBvIztZ2hU9e5T61PTKE6QIVCYirCNl37jAQmmaBP23VTDPFhH3Iax/23czsOdNgXEeFk2
eFivFRiOwE1lVTKdLTiuVyQpYVoZ1N/ehxJMpjvb5NSzrtAa/8IONlYXguExNXajq3jTs7PpsklU
75+6cMSHQ2UGMrb/9QXd5sVn4FpxPh6qnyTT2XkLhU6MHAoWkQCMmNjoA3DBpPoa1Bl0Vp4x4iHk
1Wg4XfCB6rVsXOCsVx5LAL9do7bQ9KYoA5P6IpiCvAWSZjdFet1ZiaRzNi7Y6tDtrfqPzRgqem/E
30JMJhPqkGj1sqA+Z9kZU/VZnZhTn6sPmvT2TBFUUOIxgdm9jjvpZ4yhNuz5PkLKhXf2jGcQIXuf
+ai0zVtX5a4VRIvtryiJoV77d3I9t9QrYuuvkU3bjDnhGu9DEDEMFRnnXQ9uRo78WSrijgLLruLw
ZnfP8ElGxqKqsYhtt3cfzbe7KPcQc7G5fUWB5Gb+KYiafZzupVgiLZKX5PtWcVNgyNDemO81Zc4t
4kb206jpD1DOW3tfy1maodqZRbLZvaSiwo754bZv9/QvalB8WVmI5FBKLUf54aRFmNwn9ltUavuX
XUsRaEWritMsOvHm2VxuNE1Ge9M/E5z9O5HNCc8UZSW1JOKzNy0TXwa1p9YHmH789zZlTRqCVxvO
DAEmlnDZOY1TBH00kqD57EkrvcOzxzSU/Pce0egvbGYDA2IOhveeO0lP4ly8RwRenCjjiNaPRnT9
FYUWpaDWq9hY3kCn+1jfveAEchdSmNo1q+pTlu25452JYAgK66c4Arc961MH78l7Z7RuW5ehSOgm
FQ3aOarHovJLOJigjRu7JVk2u2vW5uq4iZDEHxcnT+wCbutIqC8nxw1e3c1RUJSyfnvwf2+kW1s5
evxRV16cIDdmCBLGFbU/C4ZlopnHvT9zLJFPOxJY3Ps6DEySENGPFTI633X46ymJwX55uNrRXEVa
eAUE4cHcZFbWj4Ao3y8EGoE3AkEmkfXhTkacmQBBgIf7cvO/nIGDVsa3tmcYLtgYRRFyEnl0eBLe
l/NsQbuIha2nCJWuh8dgv4QH926UgPAn0C0P8ymCJ/2SLWeLDDVv9Jj488YPC9Oej0Oaoab1uU44
LW7IiiOgSOWO/TAZVh2Vx8uUifDhTd5EJDCJJtWL+lvan9TI20vF8oOqvaLe+gmucFzX9wheVoyl
KJSDPUO1vrBDQASOciXtlVEPtdeO74dK30Dq51onRzmeRGGbTGd79ARDUT5WLPieOVQ8IT8veloN
uw/Bd0Jh8EaSbIBXYtu9kdNKXrD7RUbY2Y4Z3U+iAmZBraoxf7tRVNIjp3LPMGRkPHEIbm66ubGp
63kNDZV4D42kL2DperOMLHBy37zFMBp8jnlO5uR1FujfUFXMjZyqEaXDIdk3A4jW84m22fnRNmFJ
f3Px0JOd8qmmD9MPPkkudQ/Q76jXe3erCd8eX8PJ2X5YeFqpLMHVKSOad6VHIN0t7Lt6xMpx3hPY
zzmaOJZ5P7S355O/tZ6lkFZ72qH68sjaNYnfgerObBHdz796RItnjIFBcOiQdegUSKNf5qrTI9ov
Myv6YJXwQyg9SpzMCG9lhmzcpXF7gYfAJdEKgyfP8v8HsZ51J46wWy3zX+NwnbqZBmaS3nEgAAAa
c+vrXpErTdSMaEXWZLcWXux1odxd80mCJLC6GJ4c35z1QViJFZF0GS9EFZWg0Ok66YqOht7aKquN
jeNK3Kah9KltUmiVVZ5cteDdp/d6D78l9mouTZ4kAgrCymQ7NR2plGNVCaIezLaclR5tUEZZEDTq
xpniAQ1JBMFX/vB7gxrIV2wjOW6HnHKLuSo2Widu2v2gQ42zojSlxqGQDNYBQTXBHdyfUcOlvbGs
jrS1qY6cK5J59Wvs67xfhBnRuSav81rr9vC4Yvhdj7g0Ln14TOvUdL/iPdYYHEia1bqpcER7Hyns
/hRYfSmhoddfWhCCwloTjEF4gRLlnIWHdal04YKkWWuFFvrCznD531URpOEZrU0RrSN1RC1y+80G
Vkkeggt9teEjHAU9BLU8t6rIeJPiH9Dkqm562qUcGCTQi+K8gphq5oJs+MjnWVY/kjq4oE8kT6za
GgkLAkMBYthPwxrTxwjkdjxIeRmovN3J1ndCHXxD8+HbwMckCKmtlRyYXnAu4dXuCc3mPXj9pY83
EZi4N4bz9SKpVgM0+MPslbetuJEf9CjV7PyRzCY0UZm4+0YnoNnooVPoTnH/ALRA7oOWVJjJnHtI
/pYHKzRiA30dNeOoZy+0qTp5STZpCp8gaYfpmknHbjtI6uE68XZMGpl+Yw3We12mnFcPv6TvooBt
QFn2tipVOH3D5BHMbK0tySj2XLY6wq3SCahakb2SGXz4oS/6+EbtU3GKfjv39Fd53JOWsn7b0rH3
J5JgZrlsSwWo0d/IT2pysTyDI72SYl6EXyyosCM8siJZGfa4SSjGrGO+RpHsmmO/ntgN0pMInEhC
AdM47dz/XN9Cd1M1o3AxEBxO61I4Il0NdhUKg8fsEesrCQV+wbkUC9MSkWCkZ6PlWMvihx/nLcUZ
iFO9pnDbnW1KrWcvuwf0S0Z965lvfTxG2u3yidGG5YneBr+/3nULouMj2EkjgoIfDLXDKUTis+q+
aDy4qkNhy3Dijpa2Jffl8pmKh3cZBYV/0Lof+5Um7iltIMZbMb9yUgYfGxsnsvzo0rXfiZrj2uEG
LWHPyUcqLMx54hEiVhns9JU3QLvNjQBlC47Qbn5/ft5OMsKHuERl3i45Is40lRBNi/O3cP4HhcYI
D084zFLOOjaL6sxNtpZXQJbWcqKK4KgFlEkvyFSIKaEd4sUwiSeReK3h3ceJb3snPivEVsAZAr1S
Kv6ykq063jsD15j8GwunPWDsu9LpBnXDzBR23dx2n0vIPe4hPEHOLVPDheQztbBOWbfABTjd8jz6
XoM8oXamAe4alHFUylKpnwiR1MiR5UnHT6N5/5CRmWtAtXCr2v2+GeQUy6V8Hg1+v9awGjWoNa+5
f6zPHVT5P79Mc2fiphuiyWTUeK38jNNTIjVqqaN3TYZE1XANZf0G17HjjTdgN+fHRcfMaKehzkGe
H0nb9qTq/5AHgFI8lF44RAmER1tm9NOSORngjb94rcmCmJrwkpHpLt3LR0ZyGygR2m7V27hutcjP
FoUxJ+Z6KJcRskQ31NCezOMO/ntqvk6MVkvySXvUA3mwQ02tcfZmI0JMCra0aJ5huGNDlpjPo1QP
i24CjutVTOnhFhmUwJbCpvvcWPYp90cBR+0yaXIc4txAtyPBHBmJ3Y+PLPlhQX42eG6Lq+R8C/RS
WhMC81C5SrbpalrK8AOQSaIj7S8GSapu9n0RpywfflDss467ReEjTLHx9kVB9SSMfVO1yukkrgnp
IfOmbaiH/Qegv4jxbO+QEmAf/bcu9V0zZfM9Nvodl1VxbeQEu78ynKfHNVTL2gtOn01ra0x8BkeW
9aOyaFXoWTOyO4PiZwHj7qY2M8LT1cuSOIrM0MTFrvSCasdH4LXmftHgXnoh0IZodJJRGWPC+dHy
vbheeAya1Q/6EARTXHDwuUyK8phLpb1TL15qjluiYmVS5IGEmE1MD+TrHzoflSRpJ20cGOkDvSnf
FxkmPMhgvDKEXcCEBuvKE3uwum9YoSghc+F8kFYXSuyELYzmpfeA0/07FmZ5Fsy7meofJnLhcbLn
f/U2aZ7Z160IKVwmsvlV5Ghe2lwAsTc5FwkqPkAf+wm/p63gJlCqqv1I36clZS2eKsNr0dQfQhoo
erxZbsf2xDkPCB88+GJT0ED72v4a1AgIBluXSvljshasvxXZIOqJqQyHcA7XwnHfda8snMnA0NBC
FSAMQ6P+d1RjAp18qXJJY7pcQjWETXDS3XM5KSbDDS7Wv8WRCw44hTF+LYTbmkRj36OnrYr1IlzO
WHc8l2t+IsOP9dNsGdfBWVIuVXty443Eb7VEILnuIX7wqDXDV2cc0bAmXvej2535G3mAtLhRu8Cu
fGi5RwpQxcjdfRf8Z5tglZ9MVCgeGKeJuwHk0McBoiFSOljUY33P/zhc6rne3k1AFzhg6Z34xVTZ
VXPaVGntn9XdiK3VtcWQM8byjtc6BVABey1hyXFOwQ/vidhv4qdGsdJ/VORqto5kz/lizBl77FKa
492Tblj+vSwFNi8+9RhZf4wZeXrTrmoVayFYqiGugF4BUFnxJKX//lrxno/sPfp/GrIyXqp0SOIR
JNaPkQMuXNhYN6gX1MXqfx+D+BB4EI/5UGEmdkwnwib7R0oaKZ4wCSYtq3U6E/cVQ/ciZacXPC87
WzHGiBzGwaECOdrSRI5kSmsRWIGivixtNSfBlrqIpp+jyx/jJ7Qh/vMj+CocjJUbkvehj4Y6R7HO
Qp/ex1n/OnN90VSG2Sqr2T2MTYvPCAMSRAYhY9QDwL29YsDqNrWSVGgHdHg8U/h7s+MJ8HRNgFFS
RCim8/hRWq1R0+TjUksyfx8nFgri0rmB/5MkXEjZ8r4xYGZ3u+W6HljArm3y8lb+P/JXlAUF3fNB
5aZShDZU78uUONi+iLCeMhcbK3FfSLXhI0PWJCy4tDpPyhEMblLbBxjir4urfLNOMaaWbu4u2tCH
WZXYbqc4cq+hNtp11ylMGn9zsrgQHbFv6j99yfmAvNO55elJ4OftZfmxi5uvZkftpMzqyssb78AE
z+Z/XM+L+Iy/UGMhLj7ACNVYXodldKFI+dn9+ifrjQJXQtPnNZJGL2sIGvXl+ud8DBs6oZHcpgM9
uJAM1FEAg6LwQ/kIpLkMIlMufLrq7gDFMPFjmikz4t6dsaztzVDCMsc3jN6QbNlWo/OqfskHNgNi
NxY8Vnjvt9czqgOwAudYlTQtJs0bhB3NwWgYieIGOLwo8dFrxTn4houtdK3qjK2qc/bdat9vwcbt
aQDSa1m576F1dDURGFrjBsEtRqYpauV4mG63PVwgGYuBfl7ouXr4QsZ1/DSo6foL40Kr//ilQDVN
vvbNXWKN8mfH1eRp2hHKhl9GdFsJUJsf+0FV2JIcjl53td33ymhrvbPsNgEgVF4suFuw8nFFSdat
AmIUMbtv6NU5HhxsXcdp/FTJmuz4gOWsZzId/yN8ii9eIAfE1b/GpR2cWdmBmVq+CcdpUqls1DUA
WZaUpMTVox1Dep9Z5G9lnLCU3FJ7BXK4Nw00dI3bv1CSBZt+4KuBzp6N/mNZHcg5/ha7TmC21Ndg
cEqvs94s3yjyZDQ3d6E2ROhnA/2zC/PKPM7SBXISh4UdHaoEO3YqYGd8zD/szRwPlAG/MKLLjB9R
6evb3/HvKEWPgVtusAE1h0MHQlz3kxIknJ6bgnrtskS4rUuK5anjqm9Fh5cOZicYVxpzT8tWe40J
7oc0VluAW1nL8FjtiTSzSKsj0PXYV1zq9t5TZqo7He2A2kFpKiyz+q10x18TJbX53TUDXwQ7DLOf
jqYbKBrJ9k01d8p0dneXvZ5x/uALGdCZHPFor5i/nTgniEq3czNY5wz9xYglZ+uJnRA896wOHWVy
FQ7CzMmWOIMYy+jJMJhcadUoL6edVYhrKZI1HM9/C0yD5KIHoXfmbvbITPKINvYd+ECPfEagx6TP
AJmDcNEv/HWzZ6kss0D24Uc6qqFrcGSO6suiQPR9QGZo9VkBdHv89fH47LAKlyD8pMDge42kmHnY
ysINlww4PaSP/O/MT8iCBgpp/2endyCEwTsfKWKmpzWL29jKmEJOdBSJMw+0MC+gdF3+aSvewVYD
pNTFBq7EdiplMyP1WF1UC6f1J1ouiDrCzP1ffHRRtiIqT4ApdpWKAF7fgUqgmbemHxpbLLqJKZy2
p8hSYAVcp50wym/GyOjzW3pv+iePLf7G4asZ7G/CgmluEqpS/v6jB/7rkt1e3RfYZkkJ7JHjxF+Y
TadfYxB1BQdZooVPrd720W0WI+HqXvqW3TaeUaJSAmXjWB30U4XQzeARHN0PYxJLFszxgoyjkbQu
AHVaEtupsi24VT5SZv3Hj5XWRdDHI3MCMWEPai0fD15gBsT2P1oVwUwSPVTmrlX8KyVggnH8jT48
BmEijFEoRgE4Z/LQkp/keMnIY627fDDbT/Wp0sqjrs7O9dgNh69qJy6Nsb3SPxAWMoBHhfBMzUEU
Dptp6ScqFFCrAyOPZnBagy8G3LIj80a6VxRZ4rE2jhkbCh+vx7lD30NM8lr9X6VfKQe1QehhvKfR
KIrzuA9MyTOJi7Xaz65BLJCz4wNnpiSsjrxb6Ewcm1ohUlXrihHp63Yg9+tKlmw4w3qOdj7bjQ2T
q3x+CiWdRXXx203cp+HXiUuR2QDTmLE0ePJoTpPKTF3wXaoPQAQfkx66pj6pw/Z00UnMJ+6cqTW1
+02jgZ+7MIHGFcXFd11xDvfjJpEeBtIp1uobFkIbbxM9SwmaDoB27OZpAkxPvrZmb9SFPrfBLkzC
r90RG0VuG8pdZ3gogE/dbbP3Ht0nrP9SjJyjGtgoQOjfxn66j3Q7ouVhXJ09vUevUDepOvQq/Uux
XK2o6kzndoZ7VkDPZ/r/J3Zsgc63Y3gk9Z3qOYUI9aqnlq4RBh+Gy1O9Mri+w9wMrKcc7PiuY9Vd
cXzm0oT6re8VGazNxSO0BN71qX3v+smOy13IaxCkR0sPTFkXPY2bonpziCT49aHK/yHAiOxywDEx
DUPtnPjVEUDX7wc6z8FpNPMqg/l2kUZm3gJxee6PVRFv0dLP5DwFplHLwEh4aPnfn2EpquI1F6C7
ICd3J6HkqwiRZfzjqR+ddnfM2gvL1V1jT7prZk7zfVLX62vQ14Vi7R/7yeMfOZDMQFY/XFfLVcpb
sktLRGaRXV/gz1y66d5hgz2kCqDm0Pkw50V4cz9mv/bABMwTgtN45pORm3jQ72vLUR9PP6MxK9zi
Sn6rBeoUU52aA5a8JIQe87RkFkuxT2O81VpS/SZz9ePIjgMqS91DYg5Ewm5ChpTTPboJeibR5NSG
rtsTEmVfUiCC04VowpYDAtUWCzjVPUjRZZwFe0dJ3nDjVopbfk4KGC2UnQOtdBMNEzbSnHXG2StE
otRh+MUii4EswOdrpFHE7o641fT/Q4XUS5laXDn04EQxYTyJVz51ociNYaVsboqM5P24yLgpP8+I
u/kTRkteFfkOWBRUn9tU3RNAcRxVeCLbRPhBBWReA92qPQF9U/YEvOFeawG/see7EPYz+bak0XkS
H3uIv/52ZM41YL1cWKY4V9c8UjPZXD6ILfcv/S9Mx6lp9cVkUG4KydODzwMBts21VhLjKaPmkAvS
dbkDuoJqETLQJIKHZteZT+7QP2qfdN2viGo7QZWRib7Zv8YFnMIrqoEnUrU6v1MRQvv8LOyrJ1Wu
qdAYygWc5A2rEZoIYoVjarQWLZaipNu8rIor2NT38DEFXQh0zuAa8xet5+Sj6HfpGuzhSsc/LeHj
at+ZUYPMj6OXx0Mi+WegFvwnnrtYbikvW9QkEO/l2SA52YR82jMsqaGub1cwZDTpvgGNXiHpz9cC
1+Zy5WJYkBgPGex5SDGl+tY3UMCISw4z3J/Asj7aJGp1glEtygDTw+ztKBBFGPo6mYUBHlnbb56t
ogw24wP29D5xH5cf+YuDc2754eH/UIwdtjPpQfDzSfVPGo5/t16U/8Bdo5y1gaC13GMR/eJFLElp
1g6rJgKyL8tqdgtgRnZ4flP3e3cJYeJ61zsUu8AXaqeRR9Pk9TMfeUNbCwb6vrLwcWQ/yu9rlBx5
KV4HB3GPm5thruxg8ZGkpwrNsY70UPiiXqS9x7bc1DkExdQUaumXbWaN5z3xMHH1S4hvx/00XGKu
HI8+3PGnSojM7x7BJWC1jqyNBr5E9rKW4Na9C+D54BgI7z/4pHMxVtuKxa7ARB3FmaVWHVP/4bsP
3KsDoCrAD/1+01cER04FlgJoMv7eY8yMo2ERWgpuVqthYW+si7ArCcRQaBwIZNm3umDZ3YkIR7mC
jtXnd7QxIh6Cof59+V1OMk/qEdcfYi1PrLQsk0bD/FQ2e0Bn7pbTZfKugANljPzUn5DOZ7KAgrIT
1Oe7IRVBGbTJvBa0T2JBctsS4LQQHIDKeJ+EfTcOMXpdk9DGceaw+YMSnJKAzvNOrycWYRDfsSgy
XsFy2IMj3dL0vcQKCspqsIwsETbF/ZY6WlT7fAbL8t+CiaZOdD4rPHiOD/kKcOh70hE+MLCYDDqy
4znS7yHm4ysikssTYJD/oMFzh283nPIbR2wMc/Lgm6kACwqdZAo2XDNYdP0BZgk94rn7xXmwzWIh
bB3CbCV5oU6Q97SD9N/bqaYFV4TcY01RWyfw0b/BNSEQZXCHwRbAv8fAurjAQbrwBOnUQPxomBnv
RcJ4dfRuxTjg8d2sCooiFXLr6Mv+4QOW0+04cM59c+4O/qEuIDGeg+lXVv2q6T/7femqj7HisbuD
XIwI/K7zL9HvBYL/0ltYAUmAGxZI3rx0KdDr/VNuQjPxMtc2X/Ljc2evt6qWneu96gv9ixdQp529
y6WXOFEOYjtiE5ANXitoAOPcYvjiFAumebCqQEi1fwcTo0bT1SMajSmYNOUTPUY2bWgpQsaoacJg
ac/KDVQqIpIF2ZaK29o8WznNk3LkxEncdHnoKyMotqHJTMdG1NCHksnuCUgOiSt3/5oACTDm2OCF
971bpdv7NvlsMDtKmspYqtqo5Ok2cQUf5ScVhLyFtL9TLQXCDpaS17hkGuQ9K8tLvWV0ZqMu5Ba7
v8j7xCgL4/vgx6VnkWaiwD7SRuczijowk/qGGaOWTwLJaVOLRSa5Yueqr/clnhvKxl1X4Pjv6Ght
+jgJhT+QcuXzZKPNkRcwWj0UlDFfdmhyziGLsGo65Qvc+U6r+Rn0+chMZWBiCrEsLVBsFhQu2LCD
GnQmS6tD/WZ+4XkmPxVEw4bMgj+njjq//9lcuZ/Q2Am/kZVeh+TA0Dmwze0vtEdKfDijShh0mqXs
nbC+TmKFfIlwZKpVOVMgGcoHz1L8IEut08pugVr0zjhVmP1n8l6/iMr01LdFfGSyjPrM/uaJXSUB
H7KOE+K1ie4iBEh6sGSNJwMdOl9tcVeaGW5tjRJ9Mp02EcOYnBdMQmIkQTdbLpyWVELM/R+/x/JC
m1wff9+ZAgJ6nRoJar/5IQhgmhaPG7psUHjONp9MUNyQHVGIgd+DVCvSFbwOHxxQ52N6WP3tBNIe
0L+3j20dfoO0ID91F8ncRJUfq7vmqV92L/hz6in7G+FI6c80RMYzamDy53MwdgCZWC2AbiyCqjiA
cCLZxLjG8DEr/9+Dy99GVqRbvHKoe8EMp+xzC6RYWo0exvMp01dcFK1nzwU0PJmuNKzd1f1ivMQA
G9LxVTGZLiF8W8cPoYYQnLGcNsnoxzfGecGQMH0FvqTY7b/AIlf1BCwKTl9JfT0PyQOt75SX1WgG
KaZsKS0hbUIL1VMw8f9IBegdN/5QiLEyrK8gjoLxGTerGkwPBPnbOFEjzTEnuchiAHBJJ0fAK3ho
cyNgy5Gv3N8QeQHGDMk+XmB7AMUDVmyho+MTfJbjAzk/5+GUqsHMgrgPdwy7xtwtr9t1Dv5bNlsg
jOPBnx61cBMuUpL2xLCX1IorzMOXHytTpf8ucA79Vab5oKIJkavlhGOq6KoJmVs3b7szgVuO3J7q
vGA2iU/kxDTMgr3fVWycTOiwXRvtatXRdV5eS6y+l7Ft+7iHisWvSNmg+pLEDdboSgeuVggQqpNX
XyOV34EWzc49L/HNGDd6BNVsIYY0MC3dqHp91QJNDvAexGESMks/J5KEDP3Wc8SbiTi70Mxp3He7
Db/7Gh0Th0gmoJYnSt323/bi53yxl4ZSVrxejWls3GfL1PlxnuQiu6FM1j9eh8zjzOxGSTxnJrwp
rTFIN5pOtRNpIXzRCwQ2Laaep5NbWW9heLBggpoAzURpsIrnftlpklw0eQzeC5oWWtM7FmnAec03
om9xud0B7CMnYzD1lh08cz4j8WZanFbKVeuMdM8YS7m2hqqkCg4+cLJwQ+xzeAPs1uO/KS8s4pqH
VaJbOvpRKJ5A+59HWgh2FNJcoELreGoQitgSOjCGFJxmZKTeZdzXUYqAh0bTmgl/47mg9vkGzyQL
goXJmyqIdD6aD88Behh4MKA36fNneVw6EbreH9PnVzlSXlVd+qXW5uAkA63c+/k+bhrdLhcVHY8z
TtP6lBOGO9mQ2AjTlOJ/lxPFDgd4qw2qM7E6bOkIFop7KnRpUgTbtKTSC+/kgR0zEKBOUUyO39Yh
vCwD/xxd2PfF4EpUD8dhLsHngdksSN/qLqsilZHqAcpSi1biygpqlyE5JxaSJlK1SDoUxAo+IVcZ
fTY7jCZ05rRpnm9ajk5tVZR40qzqcWe4r4FBoehz9VBZUDgKbtJGBjPg+0HSLd12F9vPG0wqU4dS
v41dUGAJJWWFB0MDtb7JcuBotyqrKhUoP+985MwvO2c/FL/3jWBIwgomGwsQEwTXwlHy8/MlilCF
/THZhb2RCNoYMrITKOrsda0f1NUvnPWh9zzxoJcWaqUyD2U5N3oF2uA9yIvrBak+nTQbXtjUGZM2
8VvQIoqC0m++1ddyP0ZXaclELTNw6lL6mlRuZn5XdQIK7lvKoD3EdvK7ADJn5/eCFQNOhiRAl4hE
xlYxzAWtA2/L5eKgDEZQeHg7Jlh6EyU5jvRR16MBPQfPFMny2/ItAKuij6yRGB5cnhCLGk4cBQdw
Lr+MnslezJbHh/7eo19zd1ErpCll05avx4qZw5j1I3BjXVNxjbMHy75i5NV3++Z15eWL7JvWD7RT
o9w275bDXesU8RyZcRogY3+PX90IxHA+vtfsnW9f0b4pC90ivMG5NcfAgdK47qui5te5UWToBW2H
eeF2EIwo9gQT9Tv7yKueCGpTOb6GzDui5mOkcGdpNRP1+1DEzvg0d6qQ55kBIOzYC6WXg2UlDCTb
Xf5cnknpaPymH+cd4JtpIg3sMvUmo1NL1aflEGlBJwtAbgrF5vJcJQ4kJIqF1kiCpjViD1Y7vYMT
qWRqRlZsQgXM30abUoKVHBXzpPqAEaoepDyu04JYFl41jhS7T4Ry0BZ0hUAIwY2WmW5dDuF9Tha4
P/kkrAAl2tuOjHVziQww1l8x7Ruh8DSXM/ipptay36QiBQ4K3I8/vci/w5QWd3NelOHyOI1IwrOE
lbUTr+K0Fw6eutKdIpVBgfDivg6mmsxqKAzW2hB6rTncVkZX+4j5zQAbpiu7i0NOYb6GUyt08BzX
V/A1/3LCkEZzib82yYC2vJ/NRL2Q+mluHvvzDDMqgpFHbCQQLsfU+9qoJ55h+Ebs9inWMGlqFwQ5
FCUvt1CYTo2MdeGzvWXoGvkTmFF8EPZA31aS9wE9Qli/AH10yejXoeWz5MD04b1nKd3kz7Xq+XDj
Jnlzb9ulHdAYQ3c7Sgbtfm2izxGR7vTE8R0epJ6FDr7kNkSL04Ed5X/J6+OVLiuxnF/tpyDVAgSk
bERgbPqR4fv0LQBquWVJNaZmaiRwFT1DlR13jEJ1I6oVYFtuhdCQlDBcAcyTI5h/idlvXeEuxZFn
y2Dh/+ioOc/0h6ZZsB1gsmeTj5GErwovpxorDfxHhOoq7i7iJMOzcAA4giKJsd3AFx+RsoVxFxbk
yfrYw592FrlkovHl2uoFZnAm/XLXO3zo6CcCaBy+kDMQkigGsPNl9DRBwBUYtQBd+gPY/MRoXp2u
zJj3EP+WH/R0OQ0/XLLHhWr4iDx6lYxgcbwg1YVUN/72BpZJKxE2ClpENtZtOmbANnKgwf8MnKhx
XlXQxM+T70gL5Cy4lmyENv0kHBjPpOixcIu3FJxb+HZHZT2ya35AJxJOonR4sOMrbibUXJK54s68
GPVR/evm/vdhewqCpCiDUbCppwninWDxg7u+dxZJ9rR63QMYH3fdqTQxwBswePNJEa6GVUmhxcZM
ngGAucpvB2DClf0yJxcMVy74uSFoo2ipCg41T6YReyUwamsf1eUuGek42bwrg7HU8X2FnLEGC5jn
qjEs3aGaUeolxAw0QBGZKfli1gSPbmAIfsF5Pd4W7YD0Fu/TYAWqzZ22rRr57CCVM9MTpFnzvhHg
2apvbyNet8RNAN82cgqwvk7zpDzN4HAp2tQfdfVqupxCkAEA0OqoreMToWOLEjWMss3O6yWkSgjV
xdh/SHZURy9MvXEg1LHAoVPZdD3xdw3VpsAm/Y2tVcgUMk4Hk8X9KRF61eOAN9/huq4MkoKMKZik
1s7LoCF7Dn9gukKEQfDu5mQouwizfdkex3kcxmYgNLS4L7cbixNqPCgXrbQyy1P/CJBP4m9F/VKf
rtna7NhE4uN7H5igd4XQOAyBKXqBPYtC3owPJpVG5OygRlhc7BmndKMZj0sVXC8BllhFBBL4u7aR
tg4NvBGo1V2Hs58JE93JKcbuXm3TIVsmk80yicp5yeBi4hgvy8k41trFpkvIsbOp78P9nA9zCQTQ
Mb/uNirFI6LX0AifK7LRKpbTiBy3cV61wRJ3A/PGLBZOo1yWc3a7oE3Y6fkrP3pYLVw84St3EOBC
uSYev4Rd45Qzzq4oFh+qJzyKNM8DLhJLKfeGzxWP7okW0/CasaxstJF1ZRVzdaj7GJHvsx2nPAnZ
HGfkTiEF0TsUE+47QdXh7CjDvdi5nO88ZuayjBOLEoV4FEchMlJHXTiXZk8e7Oc4AX1YLsWnwnWo
IX5FCE0Q2OfGRmcN3RX8AOqtsdFrhVf2uf6McEJF6jzzpjZknXY9Ry9/P82FHm95T0C0yG4j2Td2
tcwlDnzeWPKIA5RpBSM8KnuA7HsyAxIxgBLlLIt7FpKHDAn8tW/RW5rd9HATZ4+zmFE4u+4DBf0w
8wPxCbdYoRAOJ2PznYiBEYP+J1fSMKLME2exQnfdg3TlEXIlT2YZOQGfGZw6idEehhdhmeaFiwh4
v/xnprDVcD4UT6n3JD5+8fzn2qSjUVNyd8OE6gdqxWwKbuCu6hrO0Wf0gEprTea/CJqQ4egIPJb+
HMjp8HRYaRUS9UglUjQ7CZMOWifGjAHxhaPB0SUgq1vbv36TAw5X9yimVwA/c7yinpa+429/MZ2Y
8AFMn/R6JVVEfE1S+HbGECDgFEoLz7mcGbWgbA4oTsNGDTX9oXW0y9FnXb7S3ckqNhOJG/TEDHCm
UwFjjqTe7IM1j3PjGijlYi5WY/4A0rg4kb/ejVsKiX7thUxIJWwjAXUYWf40RCMz++giw7yK0CXY
rY/lYK0e67EZotqUj15AmOzl9jQnmr/IWItQz78pRQEXZQCRVDW/X6+i1cs1y+OBxGMhuwYRz1xt
Ik85OEmERRhp7RzIeBIIDio30uuY28agW2lYj9QlEBcHRooQ2Micr5GLMEYGNtT977/GMHPBv5hI
aG8LwaKvkMRd1Ex5KLV460Taj9YKMJm6LQjKgzJN4vth48EhYCjHLlF5q4vnFeHhjDULoM1SGApO
fS2BSsKC9weJY8IqVm0/bQjBMKPN6MKCUAVEL1OukbGH/7uGnsig+0RZ1p+98mq6bTrFXcM3rfkB
d+wSR4stGScpubRfHdEhwQ+esGzfUO8dNY8+ep3Yxy+R5YEUmZ6W8dzk8Jiknzo9NToNRh+hRVFd
LJewMakfEb9cLQe6QIkQC3JCrfD1Uu2ft+BU5chbH9/Tk/tc8DFh8r8kRLnxLZ6GWWOw9hAVGhgc
bzXzJy3/awFv2GwacJLaqMsoXHBTz4pSFuLae6Fez3CWptYdc7kofo+qKyiSVCFu76E0mXuhZRvf
5LJqf4VNznE01YgIfFvKrM6gKztj9dJ9pdKxnmrW69c4xUYS3pyTkPSYCpjIcvmolHr7C8mBO7ni
Ro1YQMnteP3tToYn/dSaJrO2HszgAORDbgUVB4RykSrT7hmrmpcbLClHdRuKdwnnInE1XXw2e0+p
tDoPXKoWKOgAnrtQohQC4S85914+v6ks72dTneb9hCSIeFqgaiACiP7HXDyESqYI6Gq87IJ2ZX0H
iMKAzSkLvNqK8U6qm2Wu/CGoo/XqBQcF4mjSQKioCwb0p5VKy12TV1iWjEVAeDyl+vBDfosM7eib
QdbX6vbGklzJf1hr/s+P36IrB3rk7mCx3VEmzMvJjMhzslhOkBNBNvU5uYz+goWeeQ0Ye1PT60eV
kutCTgL8QXOYg710JDonvVzNIFZni/YWv9ZH7fSLLryASfIYVMfkvwMubXQ5EMYnKTyXu1cJaoss
g3V55+ZORjuXxMrPr6Irub5xlPRGlblq2MJTaTcZM0/w67Os2DacKAs1HYbUI7aHI9aP3DCqz2RP
5RxfExee+6o6WLgM/pPF17QtXXRRFb4pxoNVMGG+ZNVa8VhShFbhINMIM2fMZPXqPNeCewnkktzE
LjDDJq7XfNGJnrcl8rsLThiE0HMB2JgT3Z/TcxqWnTMkMxm9DmGjxlxSMcqwmHJeiryHyVxOjmsw
luo0mUcewez490Z2+0OoOfbPWmIQ3WaI2MviN/NUM7g5iSWwBHEQgIfEYP2hxXb1c7KYG3BFhru0
WyfKCamNSQIThDqwlnm8z/6hNVNMuyU4Vdd/Q75ilUkMDgiavIg8BWYbRQi8N4cIxnZ9eTMA6X9s
QaRg3QaP6hXHkxGtdzK1cHXg3bJpeBStGHoCf87Un8LEfpJxxyJvamNpMxWYlwyUht0mqo/HZQvj
J8To0Xf2FsrHDP3LsRUpzHUPuQkSb6lH/Zci9rMrmDRBD06TVgB0DqgmsUuD0a3oapDWujhxozJ0
F96ZbbYqYVwHzymcsC9iffProalXkUcZ8evWjF6ZG/CIaCbN4lzJbpprCtkwwqVBWRRfZITonj5q
V86mklKFwenour6oG5mdBPg33KNHvYkHlA5CoG4TVW7kJDQOJNebkiRunYdYaJAA1av8WURN7xVq
gdwfv3843kw2ZFnBDfhOpcXZ4hM2ds1pI2jzKkTQM0X4vbg3aweQZOdfHgzyVJzpekyJJ1mueffL
qDE3UTolGts+FyVy3yg+trWNrorngD+CacpefokWz7JUCv1yCOiheuvNIA/iU8V/y0MP7S/cEG+h
KYXyTL0AYUu59+7yO/a9cb9xMh+LSYbxvOXXgnttuKFPKLon2hYV0BrnqgisicrP9xI0PRnNfwNJ
bo678deKztl6ABNURVKbd1xo9zf12/8DGmvIMUN06bgFcDufrru7WYT9HGpciEPLj53va0Ot805C
fqwFDw4PcexXtGDQL43mUEHHPf6SrLwP3hMkzaCAq0buv0Oz6qkPLBsYWQexyQIzsMJdGF0lQQTN
9twjAV8X/k34/Ubn711zJ4KOTuXsUAA4n1WxM1brOsUNHlX51qO/qpKDMfc8JByu83omYTxjFhnm
d8xfFgJ4hhSHtylf/QNWlsIhI6K3b4c+CfGMt2YTOJVGkV0aEMPREyYoFnltQKOCp0nhtQkgaxMq
eYO+gOJBhkedEVg5GHF56nyBdrb5yLDhw2Jwe2l8kDO8IaLWfN6bwQzCAJfIxmj/3lto+Bqp5h2d
vDvJ4SdiPk/Sqk3AK2GKkt8Du+av1kPckhy0RpaOvPbK2TfIU0uVeAKXXzPTC8/lhVBSz7xJKCrx
LGd2aNqgGJxxFwQ/CqyWWJmo9yWR1yykokN//fQE2l5p/EdMUcItZ2sDkZkPWKF3ndP5uF6Lk9ia
81amwayl+svx6xlkTdbzEdka5JLUUhWhCV7+8YAlWm+LX4T5riKrC0hNcv8zPcVRKIlfGv9qrQrh
AraadsLlb2/vAxaCcWVBdpS6zPYTbuEZHazFjx89Nyviis6Q60t/pk98ewssMmyfhwi0o2sjewM+
Nxxxq3aXBX2QgDDl3fQA8tUIf781ijK7ii/ipiHUcW620c1A5YPoobevc+em2kvGNqNhwOydmXaa
ApjPHvpKyoQajTI+/+ykbspbZP6gBmaImnzqxbKaXGz8xxf8NKNTMq2AwourTUA6Wc2VyePYFgbh
NrjGGsZ8umAlfMzSviECcFRrBEH+8taHh7464vgudu2xVZqgjjaCI1+xko9lp45g8BSrV4j2LfJM
oPjQbdiye4f070IXlgPHgZOw986YW2YEkqfeM/7Rt5y9O5b3/P3iHMkq3mrTBfmfy+ISgz3aWJMz
Wfwza3eFGX9csLZBYr6Cdjf79TV7gFPgYfX+WqE9a9iEfvF6xNGi6r/uEOgUHNwH6gzncWgc0X39
liY2TH0OA56TS06vXagE3MV8xFjDIvsWeyQZWcw23v2iT8Y9tbBvep+EhjsfDyZSV9qmE8f+gKvx
iQN0U+sJbYcKkwydfo3z+cGRsBoKudGe+OniW7F/VtKY4lFalQxpSgRKwcom426jNon63aTJkti9
FAUz3oedXMvoypgkb/K40U0rAntuIZ5CIZ5yOge3LG2uIs1gjC1gC6/2lBLU8+O70fpa5qAVhuH/
1QQ3GHpN2sEZtnT1TjUDy9NW1LCEIv3Di+DQAllyCBwg/t7B4E4QPvVbV1FEuA0bmOAytR2unNju
UbblBya1Yidjq1Loq7e8yQzHzv7uCaS+PEPpC0DnmfEcZp+EKOPMhUyP9j1+9npyFtEI3hNpWfqO
p40vLCOGqYQD8UE3AYVS7r6LUJYyreriItqsDKCDDvzBpzuiYClM2IwWUEF5eE7VBGzAW49JTLo4
WABBnxVblkc9RyIQbI2OL++Xpv9o14WH7t1DDuktDS4PdSji1B+AzUBbNbNK1TuztqW7cHp0FR3F
aIqduCnZ0qkNarPhC3/e6oJcO6pavNcHicrz+1fjCYlWqpwtY2IvFlhcro2Bg8eKtfMrueP0QtFK
n1oilkYMtL3MWRcKDqLlPNBaJjJbqh21hHUKPTJM+wvmthpe2M7SV3cwX1N6UQ0BUZ48U+Wv2Qst
5rym2N6LqP98OBTjJTxOhs0+EF+YV8m9UsTurusggfyO+CF6Pn5NMERFXFAGaarOpwnRJ+4lF4br
Ue2gszM6rKU0fJku55Ow0Lxm6/cNpm9xqm6Sae1TupRv3b4DgdYTgBpyO0oSmEyDu6+g4C+6AX6V
YY1H3PWOaBNDt4swKqX5ukO5K+ETyGOgAtIXiD79oVwHEkV4ueOAEIGo5bhjFI77hB4HNbnNkEzR
8hG7WW43HZDfpM2/+AhWiCXpSpjXMStXMkBsPZuMlTfm7bqpS9eYDaivWOHyOVEpd17uxBShrzZa
MlBAiehsdWMXIq4F9xcuG4WZIkx3Gi4+e27o1n1DyRoG9uc+svh738u1VBxt68SKZMf9mtFsqzxT
ukOgPzfgoUi+FgKBaCFUm4bOAXwESaoXO7fK8vL/IPXfkAN597STEQ7LPJOLdNcfqb75NGnEOWhm
sLyk8EqaE5DSiLkeGmbWSgSxb2FFsyQk1B0haj4dv5ZQbG+7AvPh6Zhfnnn8r+8qaGqRxU963inu
kBPhwQXxJ5n9DY2t1cBDT+Cjo5obWzDj2rEu/KJpJdODS7ZfhrHwNqKQ7UQg9m/cpBizVALcKCCd
PJ47yfNA5tx1+6osoE+pPr3oTvA99YrBaynxsaUN8harnMSAZ+tE7BwkFtldlAvDRttI4H7xrJOz
5x/dAUP/q4qmGLiNcjiz04u+u7nisymBCoHcPmps+g66fC8Z5B4+HhU8qczKEwZHphXTiFwW3M0J
fqaREw/Qskz1lz/ohqG4oM7KHVBs2Dqon1hJiixHM8Rmj4XzsUn5u08pGjT0OaBq8GUIr7SW62tX
bBFhgnoW2kN4WlG7QBQArbXarePDxIoXa363YdvgOOoFX76A0XNVZsXfBf4x6GmF/iaMrON6CroN
3cY4mi3J/bGrqv27nU18LNgtt9bFdcZgIogqSkGIGsTQoqOQ2apTlTMlSfMeE4w8FcGhz6p/0RD9
+eDnpIaJBWnxKX5bU15BzRPbZ25N2Vgf+K0dFYBY3obxbGLterfv2MitsXxBJzq/piOWje0IbsKY
o66g2G2syF86uDx9b8/1j6YwD9c2p1S60RPTXSvbOMDrFhieW6S0XJd+mvGcpYlKWOQ5nYDKvMBd
ZF1exk8/DxVhPhcL6bnd9yVwUsfV5/qR3LvoXFVYdJjdWZKue9ghwAnzKVkPd9JapU4ajUg+DWlu
LRKjG9Anv1nZU2SFOo5MW8uLihL1tifQhuTGFHmX0PgxhJMpByMDfKt+dbDY1rONQXxstnnsE7Yp
zLklnjcaEM6TsGcwaBuLSa2YZL2nzUWR06x5saN5rytl/BzqZ5lIsMZwpgd6qKrjQhzKa6J3cpSb
NY2Nsl7fnCIwN+GhW+VpzL9bkPFn7FlUWFkPiUhntuPP3KqGEPutY0dl4qmhOF0Lb84RFRhoqHd+
WcCmXe4Obb+Joiel4LhLbKLVWvPy/2ioNn1s1k3uIOmHcaG8RUpFS2p3OVYF9B77vQotdJd3ZUB4
wP4vDJaZ4+EH9vyqnIjyn+6DQUy3Ng6BiT1wXVta4eCrjH4f8sdoR63qpmk32NzSJCxzTb95eIwV
Olakx1kqwB+xvgTFd5VN69CIHOFZLX3+OGFA+8wIzZkuAuuqZbFKKvXkhcHfUh8r+vMi4sBk/SeN
3JmzmMIvYCgutYjqiBAKQe5yKiU5ettAZimTCRjiF0pypaFtF13qGggUlvhMjMdDSocoa0rx8KGK
DUlVlAZNTle2yn2hMhGKUD4ynJHoJHnOh2b/VRullzbCibTvRZfW9RLwts8Mbsr0fMB34zsfkyY9
1FMsutJxnOvNKSx9m3+BI/2WZX2q20eFIT4V/ZRe/AAkJ0qZu6YchBqfMvi0T3weTaQY9pDN3JB8
AGc6UaqxiuxfS6Iq+vUi5wB3hlU+syv+ZtPtU9+UVes6zDG3mgCqtVzgyDRkF3WB5An0bOVUeZWJ
AHhLN/hTd7dyrzBvKca26chFbXQSuwnPBxZhjqV0hY5x75InhqXrXNnOIClGTSomfpNQSl/BFwpD
9dETVv6epOjN8WlpfSpZxjjDRYnxMCrvFds0gGg2mzv3HWqaD6TCuV2Q7nywKcanDoNFqOXX3Xqq
SmW27F2PQi5DmYJ0nS1hOnNvtZ9uklAQXQSIvkyYwCFfuZuL+so7mHEsm5hXWfNexR6egk1LoPlj
OXcejQdlQ4c/QjfXhwpWxf8EwUKOfmV+6x6cE180VLAbXTV/npup2hIFWsQS7WJJXyyGEe6QuPo3
FnWrQqes/IapZSe4iSyOvKRa/uK3rFYiETlFA5pK3t368flMJzKHlT1uls4GZ/euEdAjJLOzrtP3
fE7K96OpAIsrJvADQR5g6keNkG4UGM3aIKKnGhGFYq5MqI/OJFLiYgsqLjWCavTZQUzsSAz+XOpv
MRZ/3UvPW6ThICCb4DCheDK13J37OJOaqv5F9Qhkg2cUgLyIbf8/BRk6dishjKtbxK5eER/+i4i8
zCZq9j+DenMauxYuQDpvskrB/7sd9WOBJk4rKCgCVKjId2HVxTWb9T3UqPZWw2vvJeBE5O3uG2OH
5wJquGUDpQbMffGdkbwzMsMObtKn9kZalk6QrWdo6oMyzkbM/raanC756MsK2m0IqL2byHdFCdo8
8ZVjztJNpvWk92t8C1XAY8uPhxiiZOdFdT1GWA2GIWiCWZ6AH7/gJ14W8ns4le1tXWMzuoQQDdbC
8B36TONtAQz1zVGHjgHlqWLMkT1otp4AkwYzW/Ts8Unso8rYJm7QR3pDeR/TpobEMicXXd9QGtDd
ZNRl7QiP7a4IuA/CblZaFimOifVFsVuBdN6eSk9lNa2P8q3svWytUk4PV4ck+oOfJrtqiQ1NSR+i
SVat46ynuQ5mFvXbIBSpIq4K6PHGOAMn/CkA5Npga2O6ywidltYEBueIYzhEF3oEnNqKweXJN3DV
j/uh3kPGs3XDEmRoiT8EI78ejp/IJHNHcDH4qI4bpUb4oq9XFqjRri9mOgZKlVmmIHE0jO6wLFYL
5pGlfjxYgUwxL+7LFjqp4CHwpjwWk/d/h5uiy5gzW166jEKWhiz2uv0kSCUF2ETMk5uvQ62eX2M0
GzzBzQKky3wB2Lm8Dwj342/KLrpKEc9gYDFN3IuvuW4hIv4bMTIhHNSU6kF38twIH9ojZUBud8bO
urN4iWvrEDtvy1Gev843YCAx53U+rTlB7FPMOrqnRQjpajGelV7C3GI6FmnhXuOvGZS+aaQB6Ixr
NaYcfBDInkfLYmGSMy3SkEQPtJ28EqzLJtTXz0l39H8UCeBHdeNTPWSF4+GJ1wVdPW7/CrV8zZs4
LnUMmWeTE5iZZOI04PR7NPVy3bqu++mmmAlM/EcxBSp7IlBhHRQ8gtWH/wtmA7SdigkafyVMjl8c
FAWtRpwA4hojboQsKYlnewWhDw6ofy4Tg5JDXFVMc+bPcqKdadDxaavd7FuCjiZHp9HJXaiFldj+
dUYSlp8Pa1EfjuUh2YyY2HZy4wTcEsUx9dRDS4WBa3galBocFVbRvqbndAOOMy330Dd6W4ejqvOx
xxQvw63tnD8knSjSu+hJvkKw5zxlWYbf0ATlDLzvOkUZdXbi4X5UJh2ly2iu6WTfn5Qu3RW+mBU7
kx3Gjj43Z5LK3h+jM902TE29AEEZOLCEcwLWBjz5nccRsbQWpJ1l15uEbOVSAtqFqtiRGBkNW3SP
8Tf/8xdr9GhSKGYYmSyn2tVVfiLzBB+4OBbN8iT7dqmmir9A37MtPzeeMaN7jTZOcQ8VOjKYNCqG
cNf68pi48bmEZFJEx7r2Q/fgtULu5RtNB1c13A8760XJQDHxOhXIuyooAypLRonQGP/7taYKF1w0
siabs9OthOnPflMcvSBtteFiZph1HTMbla3RTr1xr10Jqx2Ey2+Bg9/maDPGuw6VUij1jgJ19Ocg
3xLohif1giUd145tDUO/eX+ry/OO19c6j221XAlgXsntdNzAg5Dx+Ec/Zma4bwb+Khv+M8spMv5f
86Wo2joAlQgCGMC6uKvgsK9/xwozDt9Rqmi04WJzJ3k6n8965Y8O4vqpbVAK8xdecEURLcNY09X/
EYWhYsh/ppDfHsHrIYsgMszD+mkKE+mrJLWeQ6lb18toDIvE6USB16EWh0Q2u8YtbaFC9822hJg1
K/YzgZL+yi07qxFu7fvx11gqcnZnNtCj/4LE+ECmpGYNTgwInBSkqrnigFZd5PBumYq19ZK7GEMK
9Y8+8t3E9y8Fv3bSbhSsoTLFEttCFkG5eDGMQmcvCM6iOkZKtcC9tABDK87h1KQ8e2AXPvA+cHd7
k5wSQ+S3/J+1928t7H/hxOBpGW3iAHypVYS/8GRaWfj+Q/phc9rFevLX9/sVREIwem376jZ75IaW
IFuyGLqWUMXXCk1/DOkqh7nXwi6QECjFNAVOgF+b9JAbtQ40muNfgKmkaTMmHVnEMkWqxhBS2WnD
wjB/jVbc9YAiQloy7a6wA8c5ofH9maR7d87N+LZDnxIWGg0+HFFma6rNeWd+tfE1d85Cxke3irl4
Fzgb3fIyq+WVPLRr3Lg/5j+aw7Fa6qwevbZs1gxkI7e+yIdTSTsFLpRkbjDlJMhaOuGAbUJGIvck
mVscqMmj7hpZ5lm8KUKfNdiv3vzab+YsAsYKIIteGJuuyWCrC+ai6fc5Hm7pmcrJ2zSin6JxldDH
Zp3Dn4vAEa2aZ/gySAxyj1HJXtu8yLsFfQUQ0MlFJCLPSjDR6L1C8NwqRrmnc4wN4MA2uNZAciEV
jx1RvPW7td+1nWKn7Zr58vnekg8dURTnl+ZDjv3vexAidA2FsvX9TDYfBQEZKCGz8SiIJB1oW1mc
uCfV+lW8MD42c/Lu4B1rUcKcIXWA2fwd+HVnw32MfV90njaZQud9QAhjpGSn/e60yWixePw3vQrk
f8BcComFc+u60Km+7Z+nT9ylLku22RDLSF6MqoC1a8vTWDUEIMlEWV2Z3qYHqJiP7KLwVsL4SOX5
F/gnK1TDhBIE+BspIw/L9ZVQn2lCtuDx/l2OwlWD6kcF0h0Aws+wIuZjn3U8SnxDFKkpf6MzjQ8L
+cL4C+H/019QW2UrmHz406UIMhSY298YyfJxrwyqhJd9k6lX47ZBI7zGKhynzKuZLTVh2RL0bKQ/
91Wc38TgZIFBedGQdSl+W8nrKBtSdYdU/En2kqmdTMdSkDI93CoKMVdMhhStkv6HWmr5vKJmADCB
NngUU//BudldzK/FcnBzujJxp0gcwuT6c02ms0PkzFOxu7GrwIK0vt7+KKCLcIH+dm49XL+L3ipI
bXqfsESplo1TZx5F5pgqDHmZQiuN5GOhO8E6R0A0+VkUE6nLA9XtcJqOXL5zkYOdftcEasBLk2AS
XqA/dkhqcV2JyK2ZL0GeqZRz9TkAsMinlMD3/6/GFFLbO3MhAap+xElbtAy3WoVrgncOBfl/aZlt
QIOGcDWjv/HPpcL4nk/F9wq4vQlHJlPRLmx9iQjYDTfelOWsGkjQTfLrwMMaUzjvTX5d6MQ5iGWX
VNK6sGPwVCKwK1lWWj55rBnYq6jjirpCqFXZIoEzbht5nzQe/iyde+ugMMRGF7h1QK0zffBQuk6a
7eIwI+AXllYr5nxFjtOMizXSJtvXqxrpkHZz70mIxcx8HFyQqovgHPbXBdI+HAQAx0hORGxBaX44
uPvYYRV7jlh5tNqsPpXQV0yAGs5I5EXe/aDKsWYmjNqyUCp/M2UEIGRjuO7dvGHkC8HWWxjsXvfM
7Q+1Cb9YRaXPz3zM6hqCGluWTpjZuFyboVZhtn1O+IOy7+r7NitiMokhRaAmdoegBCTmdkknODni
L+RzJkKaQWyA0Gd+leU2aSG65VLLqlH7oJddNjyHmdnSu4983/Fma/f+JKRAXpAIQyMYOyP3GqWk
IWqJZuvOPZLmDWnfSeesAratQg0j9HN3zfjYSsfRlGu1r7v7/TQSM627J1QFFExAw7IS6Qxw0hhT
58iU/a5wWzYleWQvXSbojVX84K2OLz6kyHShXr9K8RooRmsncJFsLKrQY6SFkH5Yy4ZxXUaGIDo9
aeV6rFpg5VGXPTded2KeEDavZU2bATSKpbdJODT/L6/v5XDyyFXPyLiboqdUjVoKeCMiro8rHiw2
+/45u8AzgCTpC6MSp93HWoKvqx4p53V/Ws+0T8vl8CLi9IZzZIv2P6nsa83g7GJ3Og63u2YoWLZf
bNSISP6yfDgbte1wXg+YlmC3nS7/iungmQDGXeW0grKooTh3er8HycXGLVui8LkBA9zxyj/Uuhyb
6qRoSz3jWhfSX4C8d+0qTfJ+Idm5y0IQ8nXNGC43RQI7xvkskIaDavL7Ri/V49jZKA4Mzs2ZJaT6
K5quR1z26SaUsnzNIpJjqGpM+MNKi9k5h7yi2OkycNK/AEhHFC7gIJL/C10dnbmR0/MumbcqlD4U
+spzi7DXWVJZSfg93fq5GodO25CFwGN5qqXB5ejKe9HRsbOZwUJ4r2toQteH12Lreuvj0magGVr+
BmI25dENMTqm96PDX35VxBeNjq1R2qXmeqdoEfSqAry7+DvuRc6r4a03aUbBAMfHBWggXJ6PApl9
4OtejZQ/mxfctSlc832KnNSdDnMqvhx05hEFNicYiz8YFATvDjX++knF+SopF6c2wrzawtOfR3bp
1ktIo9ShAsJP1CXoHkV4AmR4hp0TojaHUrPE5QkvwGONFE53S6RVXxVrxIXlgfTJc1CLVU1JT3I6
y16dE5pXli7V3S3BQMMEiAdfU8JuqvNmqeLuzZJNiCoOBVSxTQj4ML5m1MJ7iHU8eqZUKbiF1Wgh
2C19sI6n7sqCJh6W5N2sfS5po8pX4aF3Y/pio2nbLP5PuQnviSKK0oxgDJKOlqwEm8rkJtLhrvR0
GEAO56YS+Zyfefe+H9HbJyd2o31NVFMB8+SMRy1gYxbpmoFdJOOZ3ZIuOPTuw0xhrb4vcn9b5ZRg
woKGvrJSBl+G5SZoK0oFkGO2bYeVVODdRzRemzjAmQfqV2IoO3uLoKTiKZuYn5PchXKVArwbfHF0
SoWlhkiMC69cN6hMwzsYMlZ5pWMggzeXUIq55sJrfbtb2F1X0uRpTeLXXYX5ZzyceKvVNN18eiUF
tycPf9VuExIKogtmOo1NMBOc1Yldp4dLL/JcaIHAhWxsPFjnZRrjPSSxQ/i2Kv2Sz6QWV9sgBSBZ
V9RuL5s7EdDJ3e1VK14atJbdIu93AOt05J5n+qawSt7eN9kV8N8PX5gmH4SpZUKh0O3HHami6wcP
8HX0eUJhktz1Cc3cqrzpuIQaZzqrg3A0/BnN9gMyyc1jGrkJLziR2vGBpYTmtkIDnXuDk0spAZwh
BGLLZOWWAUtyg0fPYvqE7bY3yJyQdwf0bs73na3pXac3EUBYKwClRaFm3N6S9svFV6e4r4GbVDlS
Fpz1iz21pkpdhSFh0rJDiYdH2BKNopZ7b0swhtJtCBGbU30rG4L3xrR43WU4V0HE42bt9poIyfBl
EpQv2UzS6ao8+4db7aVhQ8H9tyxzwKeaKtvmh5J9JKjITbU2MdP/4KLQ8A0kj/fAeKWUqZPw7Rhu
BsrYW70AdwGktl/Tqd85mmFrNgfECKvNbyFKOlGUBRjTrQ6O5/whvBcXb7ACEqcm7exkxpv43gKE
LCSk97bIQ50+B2bKQlR3bkAaTIngHu9/s6M+Kvdyd8pEOHT4rFhDlWMEsjTvuJW/H8wR95pVP1AL
mz2Upg5KqQ7UIlxKQer0j5mYTXboRf0fu1EMi1akoVN/5x3bDP9ydvJw5Ahz7eGKeelZ2l9V8AyM
N+vygDeUVIcWWZ4xRpyPZbGzAaVoselTvbJkzNhF7dQFG+4aI+qbICB1i06GIPwrnT1Wt3ePnviu
qXDQbXuI0z3LeusYhu+0mO4kAs2hCeCNfWF8FQp3WpORZU6fdvCieT5D4EjBgR2M4n7N9ow2RHLx
X60AB8wadKBeV5twUIiLVY4F1xr6AOy4kWOfsJKWiqKQuRTxsjV6azG5XJghWGCvipq3WH1sv4IL
UFJaQMst92O6U0F13FDnC92r9ySsYHeAMl3mM/fh52hNhwydWgZageYRym3QfTfQzG4GDod1XNnI
kVqTUR6c737YEYKxdB6aeNSDKy3JY9ZGxfOQIR55CDzR+iWXV420G0RfIzBQyuCjB94xAiAMmQlq
c/Otg2boOk5SdBK5UbTueaslEd5j2AXGwZAwbQl/vLpmrC5I3lbx0fOpiAhiG4qOcT6DWMsngFme
Ve+MK18c3thAYR3fIsAYhCnCVo+ApQ8mKHg++gWJ32bs2wOuxPfEo0BoRkkpHBKO7CBPV+MiVkjW
fufZidZmEji84S6q11rlc5eTugX0r4e6Xmzqa6PkqpEStiXCbFM4mDwH6fpbkKsRUhmCFJFfqvUF
4gbyTmqn1lVDkBFy9qXLxiYN4x7zDAFhfQ7Dlnp2S7eHz3wpBUoWCuru5uKzc3q1yfmlSA5eJpmY
UpHkNMpPCcp2w8UXpif2Jt+PP9EDYcfsiB7iV4UcP3KK/Ed1Sepg+czT+1xnyjXtdqWaFBD9BOFP
gkDyCopSvrOaAdDfW+hqmcNXeWG9EY/gCYPWvz4wHJKDx5FejwVD8SLB2ePT6oLxGeN8d3eiWECt
acWpNeXQ1xcgqzhCEuiFufZOm9lLSaf1d7xSF/CcoHTbxZsfcFgxLILL6ukrCSP8Elrp0uDEBKBz
/528Hfg+jdkW9OSQYrdtavMEsD8PKnGgfgk5Ok5qlYXfwdTL5zBVlfn8iTqfPxfUPnuH/VYwHRjk
1P6bYv285N3g77Gd9i/KneGdAyjdGOv8qTOOpsw5FgmFFtiTgdy4H2lfbpKURLc7E/gsCzgNs6Nd
nPOMUhrIoo8u06vtt06JodsxmTeGciYzhtrGzCDWf/WWYGIPkYebJCT9XK8WHMvLce9MvP5xUQxl
6gHhBM/KEsg7/wAu5VZZVthJSmHXBX9+9mLCh+oS/OwpEG2NLRYSHdnhvdlBOwnkKesegd06rsvE
cb+LhYTOOe48JEO1TNJEdudIRrpUhNiM7oUUK5ftQOxsNaqjyv4+Yv992LPiniRi8krALzVjosKJ
MDsjKPj/fRFyQs5STjqUFIHR22AQiHRD5QuFntJfClFCSZFxXWnRzO07muHgd8HEU221pArs/PLv
UuLOkNnOhi6gpjthmWQueZHfkwQ/ajTnV0zvJXWWZ6kv3x9FAC3rGfI7fDw/r6HGNBdSwxzi5SjZ
6iqR83pWIGCWCL+mKzxR1BT7Y8ht9/Y/lzzNeS9CuM1TppTckfk/lQC+ZOqbqIaqDBXH2jwJm9F5
xhU0bf7x7zHIPxGOTPk8kO2aw5hRcvJOpbI9DOQyW86d0ZtW7Y2YCDBomazl5vfaUMZRxWldjkWd
vZgVkNvS2DxOwxqkNRFILJkq/jDpeaQAYJbm1ATOfm5DgFkBxJoc7ciAgCkI12N1lAjR+PWJZT9r
G+LR4rX3jwpbBrXXbeZrFE77uZRlI75Xt731RSH7ra4BD8I/CuZJRGCHxFgBhusORc9C2jMJoD4a
JRMwUVet4ERUy07EuYjnXtaFUeZR/zBwkjlQdrGMo/YYWecVGYWzAIfWFfmJsKPsP/Ts/Qs8ahWH
NiMR5rrIXvHwICMuQvCFxQqs13AOX2ZsddcWK+pThbY+NhKU08caMMIXWcfk/3pb8a4Py0Da8Xs2
qZQaQGTeNht3u5jWqX7OwCto8Uglo5ZrhRvBfXd3FCAaMRCTKJeUuUluyNzfBw+T7+TnBCNlVdrp
O4resiY9PVbkLGOq4Bxn3fjF2q5LnnS4Nw0nSkJvviRIz3lt02m//ApLxW2ZIdD3W2Sv+d1EpsS1
wvYM4SUmOfTwcEK5iW8TlY79/fkCruC/LbR+/tbiXjXBQoVfpKneoQ9Cejhb00E40H91vYjy47YV
CNMeDsjUixGOhslxXNIUPfH8BiUvgzvUdV1eU0SiRo/OXNetYdla3ukO90pYdZvNyoZTOLGQrq2f
kG3SxDjN3bFpU2iMf8THTCW58wCtucvkzRskO8HI7j4IFHgYZQjOBdf2gAk4RSr3AxQGTkkKgJQN
m4PfJMFnRAuemAHcHa3FjXDKPohaIGi0DOR8H3djn0cTLavjALjNYE547LbGsTaK4zqrBS1SqQ+8
lF35XcdSMUaZYu8kzGZksqoLEmJ7XmP/CzbYe/M59bX2EbfU7qQygozU8br0opWzM3JaJo01tjnV
Vk8GME7RqG4OUu7lbAqioXrRUTQVR+Xr6i+8j3DDMO/xIcrd/wTH9opsrKWYtLIippLF26o/r7z3
69OY06b/KT5nsWjzZr3Or2lDXwOW/uaRGB1NrE8kieZmjKoJK2QSjsulL/sTAVUAAL1jUD4nDJj8
8QMENPvNsf5xJrnWVTXY/3Yl4eKu+kzfH3ubWc8qsDpy5ZcOLrYVwkW3XstcvZl0iH/I7OjDNpJf
N14QeY8GFQz0vrK7WSOlE1IsR6N3Wz39DZT54IxTFLJZFukMRdqpYPxcVIs4gQGslGZHorIZJ3mp
Ud/IQUAJ9ZSIMGXbrT8qTMBwIAW4ji+K9hV1R1BO5vwj9zyT6GJHXOIzy2wSPhrnsPDgeE3PQj4a
q3/ZUsn/B/My/9GDSHuxskArqcmlBdorM1CJVn2anppxrAFK3uhPzvoGuTOyaS2gfnL7g06sxeOk
I7zfB4w9wHMHvMq+ubLs8JO/TDwHHvwLa8VV9F1MpthwH8wYRIRmsCTPPKaTeBVjPeLVKxBHpV5y
l6uC1C3b9x6Yi5l/pCkZdtYMZgBlF6WosiNWu2l6hSEO7E4WDT18/yHOR7McqlM2ALqGp6H1UnhY
YB5PCGSFU/b924bnjsXvH7FOo6nehob+UpzWKGn9ZIyg+06F0VO93qnW6K6ImtQFcboaEKBl5Act
7CvEd6O+TN85jAFhUgkUiA8AVRHRAYfOZQ7hXDNkw74c9VVhxsW+UKgW2h3JR2iZVKXL4+xRJkfN
Rpc3q0Bgw63VjAZRKoTy+3MynpVXj0RVMDnKui52uaYBTO45Z2AOfYZM7YDErQXywghFhXbqjDiL
i7yk1vj/ciIjHGjyGw1BJJcaRN6HUucfoArKATdmOALvC0rkHG75qrTzgaPtHuAoiu6wKojjhRpH
Uh69Id+lUrTlhvzf5JsD3GpkEqdpu0JQymrfWGuYuEQMiKTfzi49d6XHd0B8CmlmIYRx1kzrcNU7
21KFOOT9ZJWxQZjzc4fLXZTWy65pe+pvUEPVuHF2solxrzLbX1XRcBAAvz5805ztlWACAV5o5DOv
WeRw/wYnBk8QPZtYhQF/3VCcyGrHekOTv2vJMjGe8i0n3kh1NeE9krCydxDzXf8uSaQHz5mC48qH
U0N+qdsFNCpOwWG6Y23uFkiFLOAqdz8AxE8DqQZsgMiamsYrrAmgVBlS6U25aXfP+RpDHWDIVNaO
AYMOzE9MjpDM9F/DnCasI30d5vzYk87pdCSE7KfQNnxICurgBm5eNwCFsZvlBnf9J02ODSfU9EeJ
T7Hk7SeQHFoexXqZfq2vEOn7AZxzrFEmgotn07h8cbuVOYFqY5osUhGi/JRV1Y9m6inYcELxfpoK
G0nA/Z/6CTyMSSPVflzLW5aVngIdXLvaIQsS9zO4NvfPapQEHKRAuWRCyndXfqqzo23kWoHOGjal
DL4p6SGnyIWy79jLFOv6QaIxt39E8wJdVqJfGxP6nSFoIhvllVaseK2bBF3l4Q2oFw6EFvp0YPJF
V/XpKIZkGX2Yx7Pfzz9RFgNEUpvi7XRYhbJmSGbWjUxRfBF/ESljyEpRX1P+Zqk2trtjzgYC0kzB
1xJnFrnbOb1mhBLXm7d7Xh6KYv8S+zjAaGKgzMcWA3ALOTkxlUkxuSj8efLdxDx/FaN2uvDwK99x
Qj+C0VQTi+YnbvK6woNNZhtw4NlwOTY1uNAYMb8b7r2SXeAfwnOkhqcJ6SIGQr/99IcNNfS6WmZU
AbIhbyxHrMhu9tQbZfPGizxlsuElhxg4KRByHHQIbCeWU65MaEcZNy61uBDkAtLXdREbrSRu3YEy
tqUc4zWE363G8mPSj1We1TnEcllbXy5M6wEYUBwhpMZUQMLBu56GhQ7/ZVZVbUzRDusbVZmJ+PpR
X/U64GVQ8RfNKTBggj1Wz6skr3xIblI1zB/EM9fcYDSJ8c0gbK4UvGJpDN2yBBVmThi2suu8IjNV
zX7DYTsyp22TtUJc/0iYwYZNtvxFMZj4XHdi71G8h3pj4IZrMq2GwAzi3Y9R7BLB3hLLbUi1w8uD
XsfmAHrYlg2Ydumxn6igIKnocikI6/jF3dRzBKnW40wejMurBfq72qBGRD12lW4UH8yg/z7Kuci7
645LGMtIl6z7YfezODVMKAIrCkhMMs6RaGKTevx5opzdGzji64FvNYPDYXZ1HcuDdR+IixQ/HBSf
jgTMcRSC1i0m/mU43lWIB3J7RIliQY4xM6mEZJqM/2s6AeAxXMXAytADnv+eks1M77c1hcIEi8UP
LQ62Y2qAWUogB0q+jpM8UX9c8kELWKZk2AdESaH5inUm5nZjvYm38rUnxBBtw5IuJ39028OXlLl7
9r+/9m5Rmhzz+KjtmH3mVihPZcUg79Jk1bnefS946FQ//ZuLZfZeYDc5ZijDjz4oFGuwptBKqtca
hhvKNuhHHk/YwcTHDtl6Uu4bJcKxWlW+aC9EE204a8rJPM403zb/jnwIlOMi/4haq6fLNvr6arri
ti/oH9voSNZotwhRzbwUuaAGV3SXKOt2O8osQI8afKbAUXgXAL3ZBsRcdvG88M+Ba09IGBA/hSRV
20Ni+yNvd08ZmgLeSOQV18KDItT6NTFlX8ACqmU2YvXy/T9q6nHryLV1l0YUnSi+wtyCn49zdFE2
JfPu3/mPagExATItqukU5NnL4sTLENlmYNUyzDYVLWK49RGnfkrJmCUoYAyXOBmcmFRzfKsI75Gy
VvtwRqdDzjDlVon3L044DLt72CeCv5c1SmL2cBCm146Hib5m+4LJq6VvLWDVZf2vgYhX4mRf8D9p
KBNy0cLpF1h8pOOMFJZOqF+X4TXXcY1tYhdMdyJoBmG1mH49ntlUfBEDE/jMWTtVU04b7neL3+sn
7AzcJ6wLEgjIvkP0l5t7JfIpXkc+CLQBuJ33ZCXkaP0+1GnFESwPlAtIm6bOL+bfPBj7N87NE9/5
w6qtGzXAJQ2nS//cfFibXWTirLuAD6QC2uAdGfI60OAGsk4fP/+Iayo1iGH/H8BSMmR7T9w0qYau
//iFsLjlGZvV+fu+CZBm5WHZwnsymF0Vus+MVNw1WARxfQxnptgJhLYZKV8yDcAmkWeogTy0ZCUj
9l3TjAE8atJ86t6UIBTMlhEAXp37R9MqwHQ62It7DETsPr3/FO+zPQC9TopSmBg4k3SN4Sxii+bE
A6POaCsbk4+5N+F7Mxiv4wjpnbrvFukqBb9v1EtW64v2898IpcmDXokrQOWdLpic8/F8ieU0frmK
bwm0h9L4kJMay4SFNifD6EvfgW2L7sokfAv6VubC6JApOKZRf5cSZK7RV58nAW6IHmnG+nnB2OB1
pYDKLYzI0CfeRisW9HMk/YMRyQYVfBDTlJWe303bAs8nZ5CfFN50jpVKU7e1TuR196eh0Hr36kYN
5+RrrcHvQygwkzfN9QIupLbhSp4KfvOfG5Sj/4kvPQzhuEvqOLnE6sabwCYF8ACw9E0ZYWRBlWTk
UoZGPIyV2IJ3Zk5rV/CsRn+Vl/wQSPT4F69EMc3shsPP+ob6kT6/zb3oIDjVv5V4ssjkYO93MVRY
mQaGEL1eqZf/9dyB0Q2zAd+enzaKHHw6cMKsCjQBjER96EXDF9kW2nsp3aSoFkzfKOZh6fC/PQDp
3jxUagX/dOa7HLuyTTJCJYAkKVGHHl6+xocr45i4CEcBkLZdSSPUEg2VBgUA6Lnqh9dioLxqV3xu
4I7xCh2O9P7FQE9Mrz7/728qnC3JkviElDIdtfRtYlp9YFFANaaC8qpAGQrr04I/18vxxi+l/vf7
6uvdczZaxl+RgfTx87x/coahRgyxIXo5EMMQdkWLVvMY5dsaToiB1pMSWVTz6evo3eUF7KjnLbpq
zDk1HylkFP0BvGD2XzqeRkoDMelWTV8xOMBvrWkjfKTCSBEPFmR02YMHkntipW26dchFAF4Nl8kI
aHhwv81eFm80J64k6M91G0VhvNMhDXeSc9nsDT0yKF0DKFdB5lvyew871j7y8Jk+VoXZjTwDgRfN
RmZUUDs1JPys1LJhd0oZjsFJhUl9d9aUUYT1w/azcNGvae+w4Mnyhw6fy88zQP5B3FCbtswTVwWm
v/YHp5H6PGKoZS8KhpfNyS9E2dG9/fcg5/RcPt2RmplZldx1JdVkIvC0NU5/mv4BVr9hEJqnBBED
ORZvFUImCseP6mqp8g6p2mtgKU25W3LcXvLYPCiIEOIRy2U87HIyxNwx/ZIIg95fXXuwCTuxsTrI
oN1ncHUB30q527cD1Go8AV8zo0xVk7ZH+0u7uC0Uzy2MA3BVFfSH7HR7VT2iTjzqwHuJOn5PsZma
LRnX1t+8rIS9AwtFiZFPlzAxcQMFybgJIKSaeQNk9iebgPLckjBXkXax+jhe7giEKvRIUW1cLcqt
e5mxt2srFOUA7s+0LknSm6ujCFTHEMdPMnXETLAiDYcikc9JJXNTy9eYVCPr9Zszw/tTFG9YJ7rJ
Z40LPr2LIhi3zHjiTl59+MgqYk2mb2MiM5hixGbY3sX63v981n9SrvpsTYx0TPETeOB2u7aBX0XM
kf1cjiA/MboN5+H92M6tvHKAT2Qnulh2GTwR6rWEmIi2+lw+sPYjvMaTMLY0YoyigK6PbXYzyzm5
RYKUVT1iDbaUrUoaHSzXK5LFKRHbm/xZVv4yvQZcLoWAWY0Njy/xOBenhFB+AyS4iRbvb80KEnd/
v0x9clfO7Sz4S1S+WX8LdUr54cNz0B/eHIHbJc+MRhA6LfmVaz2Er+tM9EEx+sYApLT0KchnypvH
NaCSNNcLxMmBP3eQADW24os9NYz2DU614eo1p0s3iq+/xw1/2YzKhy95vr6o/T0rlq8qeT2t1idc
rK9YYK7wM9MVOJBjimhUvy2GYgJLg9D1+MLGu0+E0ZM5XZKOcHeqjsGEJduSfRfzUwpGXW5pCaJa
mnizPgEoJNrb18NcqpfvFN8grRwG17Q40eYymg+pTtZD4xplTcrE07Dx8gjJ8FybEXkNte1UFzfu
cVv3tGBUy2dGaKtDqnSP8SaJ72PpRvqEQRhnmqdims8JcAnQ1RPwKpesFFL/RZ7JGY8joQXG6GjC
NxvtQlidhAz/3oP9yFg3VR3YWH4k7Lcs+hOnM21KAPD8fGscaTg69k9YFkrTszTSs7HpiGfgEJ7O
0Cx4+1HItckPEzgn95oXno2O8ivsypdYVuJGu5HZ+BbHGBSlfoeimlCgAKGTCO5UcGRu9d+piPbO
LHUMWjsbQzuQauZ7yIgdXkxB7hA+WFn6MoscxWNkirgFqqQxPtAdNJ5zN72WC3McRN4hpE3hPiti
2lMrKYpxFCv832hEl+z1ky6LSZtXxX0maJRUitepF3Bee06mAjT6kTf8+q4/XqSVLwSAUeU1WLLP
ox6izrusMjo16z9gsnTzgQwgRmiHG7fvDJoVudNFuHIrMufWetPnPHy1LRDpQbURnVULhbu3L9Hu
EOXiCWbEJyZ73xgfOOmh9JkEoS4tAjR/JDKn9vnmXDDFJ94uNZ6vaooFINx1MEEkZOSdcEOgSnhL
+HMUX/ywSGyWd5sqQaYYAsc5rHBVXu9sJBHGLsrc4XT5Q+HBpao95ik8/Xv+lzYzYGzCaJpUIXK+
1l/NcZW9uLcjTpoaJgC3QFvjaVZRWOjHmjCuZeqQ7HV+haeQxStsjrw1qPexeqDsZGRwHZEpJUPD
UESTHtz6a0ArxXrwHlgIBZ71xdWWITrNI9WrlU4H+q343GYImyNerkw3C+ftA1VFEqgfzFj8MvdD
zlB/qYycKhBo1GBo1+X7gz5ZyUQ160cR8TmbWdCV2I26NGIKqx6Qu0tcpcroVuAsvhcSmYuZra4y
TbRKbaUkG5//kDLVw9OyHUrl58wXZ1H5g2Du0FQwlaLgOsvZgb53WWw+I5To+mSsip1kz3tkkmIf
3RYdKfI3JJTSVsHiXdIlTywtTaQq7VUV9e9LchvSu50lKKpSkxb1k8K9oV4UatR/HuIM62/8/9fj
4V35qcrq5cHHJGJnOUIF9uD4VvlRz5qedWDTIo0ewd1JRG3R9v1BFfQM7ZEy1KtrIN3mQv4HA9hM
Aeowm/Q1DEuM/z9UQxiypiR3mKkOP7AC7hzn8p6jcifXnY+eB907Bfz4x5EXGcwHlQuHpmrAI9O0
4lvX0/t9LbBuuMOHBdHulFB737pmWbQU1Nwxo5wjgNeCVJ9UDDGDvAGuDOxsxupGE7WbRFYlnQHa
3+kSwY78fQM4jnF+3CcCOBmD9rgEOZOAdQhrSP4rEQbTYPJNaj/+uA0ADl8cFA6YM8dtvSQkI+ch
aH5N3yV5eMyYmnzYrpP7CKXH1jWRww7r9dlL6nz21ANH9P0DM+t+a5/+Knu2Po5gGT+Q7JlDjGER
/NUPP2NReUvnqVbkQPkWFgpV9N9ld7yVXZED4WQhs8d2NBTniBoCg/8RKSZmUY60mg5XDStD9Ymk
OrIv3NBCBbx1WlG/BQ+zt2mLZZUniRw4AIqzpE1UstROS6P+J5v+GB1aiSLbmsXuMr+fH08KZOS0
PrhcA/1Wp58nRonWZ4j8rlCpbsOebT9hPSUapc3BuBSMYXd8/lP79v9gHWK/G1Qau/UecZ6+cEm0
9BFAg2LWuKuab8WufLlxquG0GHeEfn69bOV8jwVtGL1CXG7ANT2A+tKy3S9Ev/zggN2VbNXhwtLy
f5yIkOOhjshSmxlUmyurgZz/97ybaO8slrHCp/paan6urSVEw7vWWbzKuoon6Zst1QZdUGEYbJmm
q88BKV1tduyI7a9nMxIi1g7eKxCnAf8t92MCgfcfZn68S790luai3q2wFbN9OUGBnIpXJ94hMEBx
hudu67OiexS3HmAVhpEp7t7EGfuuTR/VWwq5cACPuBiEAi2a2rRafobGeyQZezk2Q3mYTzU8+23Z
E1cEvNmpgbKYuHz3BftHBWq6KzB4tUNF9kOwtjfcmTMfb7FBfyMDWHFi/WG5OR/dJ5tlqRQ695Iv
kqiDdE61f2zgsrj+pu9Kjud+25kf2TBy5INl5Vu778buD+JQdhoFbvk5Pm4RG6LnB3qGp9xm7++d
FCN1CJtXn/diSAnp+X09yJw1qcE4BDOrgWlCX3+kYzot+OexNNmrl7g+8dKTJwZWO7Vuod8BY2rU
BoeDEgkSpw/72wj64xGBSIlcdUhmJc0v0AKlr5DhvsFdzgckRIhac5kkazQF7fTTAo5tgwTnmlaW
sKwD7V5e8mjy3WFU7W0neNW0VaBDOyDusa0Vb7G+ESUu/i8Or58QfFCGrOjXSfeBZVDTHjqEKnnR
gCdHfXD0Miwfi8T1pfBnWnPrBG1rqyycuAeODKzk02J4QQJJkQAVwrcGq20IHQM/xdvC36Kr98g9
id6D61znvsgiQw4+oDbiihXPPgslgKSEk6XC8EF6aGbR6tlaIuBj9Q7FsbH2Ndx6ZngF1T+2QCcZ
yq1jiBMyk3NldfWtHEoUztUFG+CiNttXR+Nt/fChmdC9MYFOcyC8zWE5K2ZhTphaCLe8d7uJZ+fG
Cul99wqTNvuJzCguiO1JlZHAXoGHO5I5G6LlKXnlwRM0A0ZN8cI+DER5pCVRNIPPzqISUs2L0J2p
MELK1updw6iXIRWfg7vOTmadtVUuG368xlV/owz5NxqUaL/jAA4/SRs3Eycwy86GbzyYLmiDAdB9
YOUQoWLxa6DK5RNRA2+d/rNcU8B+ZafIvvft3RfD+vjxkJMfEiqbcZuPUWFVVcs05EEiHYlMxgbY
7OzjiQNqpZclPMcqkVxZO1xp/OVEMfVswRh+F74j4brbqGaHvPNvEtpuvmfOdV7USDDQvXj/Rlyy
7AOFrlUzV5gse5UJj2vcPgGWFxATVgMMaf4f3eZOaH4npJhzBTu070l2il9gAhYTc/as7yAH92Z9
cyHtoma4YeN51gE6kVW0Ps1CcePXgIfWLfxu8uPDDHmssWSlA+tnqWH6LExlFnB2F2xQFshg7Ete
vOH6xrFc2GWabBtY6cZAGs0eCn0yU5O3c/ffwmo8jlZBq6DYNInOc9u5rECBSZaB4HNGNFuPcK3o
VwGTPQDNykOmuPzAPosJTvh3SQ4I17ekRgsrG85JTigT0FVfAagK8GVs7aM5JG29oNCPRWFl5n9i
muLPwD0nlNamY/yhy8egyThvXBOL93QsfDSEkxiBOokXkW9dnT3LvpPITe4iLaIOWkNd6VrPxMo4
tMZ/NVwXOtegRaULuPv8jx+hV+eMXFc1evYVSIyo/HOp/hDCCevO2wuHH7Ixm2UIgeb3u1tP7rBW
XTESLB6DrGBZ0FyfXF24IjF7TgFvoHoAEe2xzye9KMBRBqxBn3SAsNBMQ1Rs+FWT4lay5VVu4SeY
7yS12CDrQtw3GZpGv7SH6lvGih1RTX5szOisgQm+e4ewwyjWPu3VGKq2gIhO/vj4ZoPG9nOzA6Aj
lCPFNg6aWeokP8cMiV+CbqBc3hwHQKCT4yLRK3yoFOkbQVGPGSrwrsNYG0BPp9OjJT1fxY9su3ID
ss85tj+0rv+5hHhROBrn91rZaVzxRFVUTcmgipHodjWjLgxldZMm1lbSgov4jk8Ov7XQoZsCHZwE
PLt2lfo2ek+eqHVbxm//N8eNPfYuiqR4GAwcJtB3i59KTXXKMeib3IJ6eAF+6+7jCuHK14ryv7V9
6Iywv5SjWcI+Uy/M+fwzlcX2TPJMqqCuFJXmY1YkMEO3BQ0owQCr74YWAaRoRd7oNfABNWhon5TL
C0QidLcCRNdlHKg5yp9hE9OolYq70+Z1vefoTCIP5jjm1cgBMVGFj76H5i2v4pY7GzeBr24QTCMn
c13x45gvMYIlNQCzpjv1uRde2SOlRZf77muyiYNJwID+fRPl8FH9DNkN78AZKFwwJpDJcK/6nOs4
zbo8zvVskZzFMDeJGTsB+I/S+ADMqq8evwrb45TABeFTNAJEXKj3lEih9qeMvmh7+YfIfd/Dnjxj
1tFA1wGkIr9jaLGi97/klkvVgnUsa7qVDTujLmWDqZqGcF09ZHCafbPR3QMrSwguQlUKDtQdQyJp
oR4yUd14c39xoL44LxzBkaqyyPIyWstPNZkv1G6KJ09+nqJtHR3Q9NxWqSiKVfsFs92DH9ohPA3z
z66VMxo9AlrSGSn+hqR/57cdnUvCgXiiIhrUb2rjfZMT5l9D27ebwgH+ohpkV5oCIBKOpVlUOnMG
m71yQVG5H7y6uAjqCDZ65VWd3WugNZLET2en/lQe7HiCA65FQenXa5y25R+929nGMcrq6b/4DLnX
XDsdRoFB2zka+hG6vdULgK/2uHDWSW3l52lFr3Um4kO0rV54W4DGu+20seYe3/1MLyDDegD+VrwI
0+xNS19YyL6zuc/7ka/Vj0eEFt5hnTie2E0sY6a6f4vpkKMU7OXTm+cMGsymyUMCpDCP3Q8ymBO+
9IyLTGxT3ynXt0wO+Zb8nX7j3hwDw5puhnmJPAQSJUsX/D93mgEAXF2krLmNU0LlsyB0oqAp8BmB
8kVT0+XD0S55LE6+DsiS9hLKmRNCRLnBFAS0Q0QYZdLoyVH3ZxXSLd+tIXz73Hsk16qYm5cv1Bk0
217B+wTz9odOnteSb6kHNNGujN0klAK6mj2a2ddgtrSAEAIHvU7zRjG/Sg18WfaKetd222ZZDrJu
8be+xltZmRMeQDfzcyUcyfKqaA6Yw95ktLSnAp+qISc6j9QQSmqgo7UMP/UjkdGxZW2qPdFFNzTr
Ylu4jQ/tU6/GEXh0ZXzuk1bkzLlcTvpcW3B6RBt1fEsib0F0QCx5qc+Z6DB8/6MewX8Fi5fU4bQh
JK4RzSRbGe2eCpiNAzgt0bQhwP3dyozcPzu9Jbrmx1Eq5ErN9V8GKy8DVWPOEnNMlAkirwbyJBlw
uq/pw794W6A1kBS1syHDAgUxDN8yA8k5yd9hrejsHgndwPQW/ezfv6/skBQ8E+FX55DjvHzg3H2Y
14QQP+HtfuR5HneTxSHEeznAIr0S6NdNjs/4TZyYopgsQFWfUADKOxxtZ/bCDVvGny5kyBIyEea5
gBG38ZgVIBcdWbqOK2b4LLXz+5U8Koe274Tx3Pc0mXoPY2UPcUMltfurNGUyB1GU9GdfJsqEz96b
W06h/BGLvBCKimCBlO23A+KrGz5oep3SG12QPIiEcSHqktOdusP96axe9+p8VC6T1tM+CQTcZx7r
bjgUztf0TCoIiZwvROGKjVKG8zeDTY46hiR1WPwu3Cjgc7blfWMXxpLAXwfEJHDVQh+EQs0LPP9E
Ybo12T9J3IDPMqgUgSHLA6Lx9e2Qvju2djHCjTyghl2HBdPkdy2l4c+npzz8qvsNKly1irEJKo17
vnJfx0dhECWMng3Ww4iI86ZZgAL9Evl0LrWNBEoOPFdyHEbUI9Vikf4/tN0SWQXSkhO5poQjw4kM
9wxKs/Wlk1R0RemDmoYAeXeeBXqWi+rmCmHZYHvcCX5dYfEZJwriikfg17LJxka+qOs6stv3Qo9u
2gNQL1NAKpYDRHR2YMfzKfVsIlG+dFGuWOOjiNzF54twGeu2OxRLItL5GhDgSL/zvIuhEeKzl4oj
Pe3UgijCTGPdhxtYf6O//i9j9ESpsl3oQRh2n4PNfb+t2T3p+AepvwtAt9Bv94GUaLQgKM8YiXDJ
e7pOUHtqXlhx7wmUzZJCAS3TJHHJWAjMH4AkXiKjs00iKQpgEtUHzHLWz7OHAWTr1WJ8N9WNUd28
rDist38kDPW/XfzWAwtqIR8FQ7Vht/+BlPt8HXhakTkreJcnajV5qNr80SHYnpjCV7WEkV9dBG4r
szDM0yVrjm2z9O7tIHD16UoRj/+0yp7d5C+4nJd2pGerbf+JD/B+87vez7m4LurFdAGZkFg5+x6w
qNnTuBtUWrLP04jiqFcp4ksPNi0zPBf0f23xXA/x1H5hsLkVfetH8i4WkFaVBZajRNydRo4yH6kL
i0jVPuqp796a3Ei7EHkn/fzcOws7hQSP1NmXn6zP/2SPXB73VQaVG7EYsJyBIukrLAJJI1suv+Te
QRECNuZBXaxqf0hbB9N3QfZIOVOMUvOah6iia8/FIxC3ygtr+z7RBzEl24j4mQAJHLw1AHYUJ8Ud
ZRLJ3387lU+mbD9mDNTJ2jXneTdrfOPCRdXiDl9X4ssWQNtyhSe1ypnkBSafUxZCtqxdqjaDW5KG
CA3Bt83XMl2tfKm1wucxe0JF7IznyGNlyVIBeUM0T5YcpbHo+JJg7edhWJjeOE2gIXO3SH0rz5Qr
R559EDvd2KAAb74CJeamRnx8Jgr3W4thPjl+YXyOPJM/8neCu2dLdMGpLx71FEguZX4AQn9AINMp
fQScCWuMlLZ6aiCjupfSoiiJeKACDNsaRJidyapXFgC+1OSvc7qwojtFeQaVxivdVwCy1rC5hDMi
xXtF7Yj8TGa2HrvMGJ6UCexKRe7kqUIvBsoUAC5j4FMC0ap1WoDS5QGUogpmNAJ/sry+3V8GoFLn
ymxQBhsdi82M9IGA2doPX0qBvKe+0tbTffp/4vbzsU79Slmyh0ybAyJD6hKmIXELhaReMr0F5fCZ
Fm2c4ISoyl1xJv5bUP2GYWrAdaS2vqcT6de967UftyhoQNo8E7NOqWqecbLugXlZr1nEKppc4brz
X0WKpQOf3nFZkkK0uC7K+jKNLUK6J8XzC/iGFMw9kcl2rB9KsyuEyq5U/cebxR8aAxPu1tti8NBV
XWQkAXFI0nGime0m484rdk//lW0mgW+F/jURVKoipK+ma1SsaiESB55r7GqkuHXiQ2psu/XP+bbk
oCJNIffkg0DiL2mRqXXY4TVZHUOZ0rJhFsPSIW/KGq/ez30g548mGL2ZKE9UxHefv3RgN5mDi5U/
94r4dpo63fOLwAdYMYDOSRm7C/c7K+KrKN1kaxZvr2PGUY2PsjwQyPG0zu48jBM/fJaLGtN3XgAu
/GCa/uj4fJh7+yHjJyRJ1zrdNgtKktQlkkqZDh4qHi8MP4Kyrty6QcGjsU4JsT/W3LpxolHS387H
HHEo8l+qp523g43pdM/5T3W0EK3AmS7bve5PWJ07bbSyEjE7FeGvFcRMHMn+nJ09D6uhUHrjhfqg
IexuKyYirKK0BDj6H7JXq8+PbI8e8BOP3G77bQ36mQm6LhbcGHl22i+1bueNUdw1pzU0DWEUX8Xp
4MKwusxVHFlPAAMiJRurHh4sByptDV/IuGahl668bLm7yJqUtvLlvA91+C+DeWL1YctXatc2gKbl
ZLBWeIOgtvtqzUFHcql43T9goFP3l30LGeDmCITqV4DNN0jDNesRD7qNDaO9Mql4wL8Jcc49zqfD
xxi7Ud118YexLl/zpwQpgXH2kbJA5yHWMfllKM3SbrRr8glULN8KbDdK5bGFhaALgil4IXXK5kBe
ifsg2xCzrjrPrwdxiE8MseCuQ6NUFbAruk/KME5WzjwJzm5WZGfeoW7UQj4pLdmS/LoC2QtGrE1w
IvomoTwvoEuJ3ePA6Nf2V8Hsk1klJyXhlF17Rjg1VfoRRCMKbD52O3LQhRLAb0TbDwbW3YRu+wxY
Jq0rbpWjQ658QyD06YI4HjQb1Hf32pyAy44UunAB8KpDecO+9ACzC6mceeiPlzif2d+zKEyFSkJr
gz8MmuEQAefIgB88Q76Th1pah94iODBddtxQrFmIv8JzEwbq0EYSOjn4QlaBxtBMXeNmh9a9wRbW
Y73jH3LOIJ/iBRr8Sfpnul3EB6usEf15qkPimvU3kYXKg22IcqWGuGMu9TE/jzhMvkKy6oFAbDhW
aV1S5EfJOMh19E3d2r/lofB2DqDk4TH4mF/uRuR8UOpQ3n8FnD9LzUmLxWU+/5uE/0LKnbq+opm5
VCIx7i1/PG0mYKVTU3Fjd8Y8c9ONbd/qcsyTKIHla43MeepLA8RbMsFcbj1j+eugtSCYV1Ghlq4y
VmZJteGJ/bpfVcMmEWdqOOIiE172oFdd82KiunHO9h4ybIUgjyiimSVNFS3HQhmcz/2Z4NVTF2pG
WmEygy3OTWBjH59OC2YSRgz5n9JnhIXkMqkCZ6691D8iH3QUsoGWQtlunGpPF+ZjnMzUIlZiUSTw
A4i+7oZm+V4KlvxtTs9v1yDxIbubDXVlTcz5/Z1IaOGSXRC3fRiy7fCcZ34udblArH62kc1SipEs
L8wt800EEgxpNVgOayQ6Ad7BujimD6z4264pEMBvUxruHF3i0ZTJFVU/7zPD5/mVDgEAJVbbdGy9
KEnEDBV0d32MAVONnvGUgW2MnYWr8tc322aqukI6Yhm1VBWY+sKxAET4ULgDt06WkAvf5hisc0Pf
9WVXMG3mkMaOggxyG9GNy0TCdalVbEbYhWJo3VUlApzSU2qORD/sfdVIcHOvH3Yuh1SdcG6VPQn7
Uo/of2kWrJZe4U12fJBkkOp9fd/RTNKdohJEoZ9F+/8div42a8Jm7cZ1gRgsOilbA4P8oXVe8uHJ
KFF8gSN4mUdsE44yYumE4cCyWkI5bfiDhfB9rEuSF6PqWnF+eCjE7N5PrzMwthvgGI5gz0G0irzL
Ty/SwSI93CM5dPpweuaAwYhPyx9DbHvEi4esFxjeGMvCEFsXT72SIAGzIjgbY5rctdsgd2WKmYJ7
aeASx/FmTUQ8qZYBo7vGhBOIrBSjjTYlyUyS4fR3ntBdBIErp0x/gMzSuMqyMHuPJFdtVYCFv9na
ezfTQzARHvAfHJH0D7VR4niTYegvMOMfknxhQq6wR3ffXfCp5E4YHN4oxuByzO80bjdrlE82Bn5Z
z6vCYLcEPNOJwKMtvoS8MVqUJpVWSZBpZbIQgbT/a6IVcL1QJeZvkcNO0F2JnzQbepR0WV+ptO8z
z6EYkK6rf5ftS05cqIi302JcLflKAWWzKP4HHPGKfO/BbV6wqyosflsG/SzAcyl7W4iwrCL6Yyc2
I4V2c997WlTpW5mE88Ksal8ZLCS03/ugWUecJmrCPRuTryGSLkA65KRc+NC888/WoVWOMbMmP0R7
xzg7z6wB8+8KrH54tQIOsfrUGThiWOKSe3defRBa8kd3LzPD2S6hxWFzwBob8bCjHq2uWDkKHWYQ
wWL6C+ckSci1CWcK/hdZsAS6Wjm8AZMM/1iSVhV5htGzO2T4Vznn5WU7qnUdrdHn6Riwycr8rYpD
m8wy5jqO52LKwX3aKl6jy8U1kZ9ZSyMkRXMdizl+WxRUBPTbCatnjUa+9pVgFJ7ESO+FM3r8AIrl
PGL+MHH/b/VttnSHTltfjUVmUfcI7MyAkSGVH6hDMOwbsCZcdeTa4HONDst1qiutlnkZx3kJ4Aw4
R5ebliosTB/vQ/UrqdhmxEYFxYOCLQuLlKjRW0u5KFV/bJKWuxXCrUsgOGnGOrxQTC8LyfV5xjmq
7hpX8UmJDR7N2R7/7pKQPewYfu6QNnkdNs70Mqr3oRuZ/8ieIToJUsYdS8V6i/tCUMf0GRF27vVl
lXFeB+hwjz50fDqIThZZlNPNWySjwpeM8eSLEesTCOU93puGU4qBbh4f+SJIC1B3Oo1Zp5uq/zEv
N77nq61MLuGD5/UUMeiapFvIwdzXgSnYhBEvRa9v2v2LH5ZUtHwBMDCVf+qCDKttSiaudFRAbFVh
bImFdb9a24iKYwin3fOw7az8SMtQwvkCAg5MfPXs2jvWd4Sjv41J+C4jNJM2M7kKrdBpY1tHbggG
5YoH0gzbo+aA3N8pYZFLyPJlp3PqwxoDZg/2k8qhB4panVwMqfXQgE8HoCgKZg+iaTnmtid+viMU
7N3z0ko1crW59kVZTbeB0wrIgP/uiE9v37708MqygYwX4nGTZ+nz1KA1WuTrlhFxHg1u/G0WtoeB
5RpkvNDgH8uqPpbxu7RV1E8DMS/uFTJPf8TE8Tju4OuUK0Vm4f+2Rt5yP5tgdkxlQifHbQql31Y8
Gm5FdiSzXsYPxWUeUIILv9iSHei6f8r/8VQ2Wsucny0H1aMmAaqkEFyCmdU3EvA0tuMNkDjLl0DI
H25foYBc/r9rXY6/c4HSEd1UNbpGNu4EE7VTRupL0/B4TnP8VdpPKuLRyoLBc0mLXPIHoXgbZ+9V
0YKfsfGQIeoANGEVr1XxojIdZRnlcd6xpLZzeic1/ow5QUqiZLeHFpZ/5uJzspK1fAFSH9o+wd/A
NAM3z4+ce3iRkF1ebbuMwlbt8QAUJsfnDNgVaGQ36kFY5wKAWHZFK3PDOzzxRNULiyh1Nbsv1K7T
c8Xcfr3U56ZStY6LuJ3nfs4R0YvzXXtUpDcIq7g2V4jHgYFbhB+h+XPlB3TJmI9Dal7gXJ7a5m6u
RcEVH6ej/V/JDWgJRGnZDohtJ20hI/Ix6jPBXyMwcHH+m+x5hRuL/3Xrxedr+aXCjeajk4WK0rnj
+he6T+PeQEen4qQ0sUdwyFNg7WT2C/VP8a1Gt1QAk/95wUa7ZPGdqSOQII+cJHBM2G+Y9m9Qn+vM
lcX3AImQbOavtLfBp5zFnQ6auYTyky9qKvsRDGcgklEV1Zhlph9sGPojzurzcY/zoCTQVC4/Tq4r
unNIvY66OoxugC5PVfkWj5W5c4/zO/tmzff2INjpWrIMf6ZT3VGE4/Z/kDhKXzCa1y0FK//uPfR+
LosNXt0kAm1t2hXAcCDo+iR+Q7xZbuq1Wn7AvrxnLbSn7Y/25t2aN+A//0z+WqEQdpxvYXwiqu7q
Q8pL/b0cnxw44xKuRt+8wpkpQ8Z0/uIOFkOILr90cZ1DGsKps3O98fSGyyIKGKA8C0kATEy6L2tv
jgF7ur6NJF1taCXJ+w5d6yoSTbYPXZvyPTkSWB7WNjlEFdUdzKjkKd9fsc1J9pw2S2dyzvMoeRog
zi6xNe42GOO04RLZCeRpF9TNTb/Mf2JpeZLCIIj2SVJji0TXu+hBRpWULXT8bxOOag0dUMkteNFu
HZnRTntEG7b/ywkDE3CaKg4YQ7AgbDjrneo2ih4JtxsXYkc+JghZsGwrV3mytphb/taNyuHo3ZMo
Wl0ErjcV6s07G7DB6s0I4Qlf9A1o2CkRKXePqCcCTN1q0dCQ2w5pqLjnyhnoh00Qw/oXtKGZLxuI
v4JRgVpU92maA12Y/HZaaERe8URYLH/qKaJhWRxOdDVEHXi3ypWbWgTFFLez71OdPehm7jWHF5CE
QO1r9ZsyStTQGyLcv06NM6wqOLU9mCtbedMc2dp8zji2BLAp8pGESbKVAxRSbmw00fGOmU9dcfu0
DF6JQNPSh/P/lklznptlnXlsj78dbl9/jOZ4EWnHavWJZkX7UwK2jHQ0+T/Z87Xiz6khAqKreP1E
ZDsH4y5EO2yLLS+48lNPqtzHCUOJm9i1HayuZOqF6axRhO15WwxJavBfRM3iWdYxn/S6NKxI3zmz
ZT07/CTC4Do36hf21kMNW4w9hEfziICcSmlYww+fY9qy2bJmqnduA9ZHxnt49zM3z3n/A6QPd0sF
1tYzNOXdUE00VyofW0fSWEZQFbcGr8XSazVROtjBTFYiGTMqhNsAkCCqVm1vu+mUpFtA0SBpzuAl
4YKkRWBvzkYarVgyst+KpUoEbSnJtRByEQjdKjWpEBapCc7Om/nZFxtdljKD7RYmv54n07Of9xjH
iwhJ8c7js7sJCEnPCGrP+Zg2ZXenb5XT8hOEd0N+rT5wREMRqQXhkniTjGxYTAta5HCl17WN+CYu
c2Trz7vyanUNwXaadS1lWnJoIVZ7U/7S13JU9Ti9nlYOvp2kIYcyKNrJ/UqBpB1qSP0N1eFlTQ8K
KSWAXDIu1dNoFe/nAxv0Xh48JsRcrwYMls0C0fkqoo+Pr37Qc/UGDiPxuKc8UPsp1nNe/A7iTlhC
KoFoAWIw/hY0/x8F0DmYYGg8uOFExYHjV6OG6DDI/XTwxEzx+Cg6hiIRNCLxX0IppkleJKKBPXxF
ASMqu7vcWYQeUlNt3j95+DuAqKMfMPC41wbiyL3+9K21gWa02jGc5QykzJwrUtEwXxXkx83UXAwN
8XenZVAGIfb6gn1215CueRMjN/AWP/42PSi4vMqo0OOBynnOnpN3f+ECdotmsg5aahabmRD/Lhmi
t6kYJ/ZJr+1u33NMs2TZAKiWoSa9JEyMrF2ITV3ZPMVLAclL4cNh/uwJtf5K0L8O3+JzyFdK9aIh
UGkoUzteK7D3gXkcqusnYkUWG7plcc56lwVY5KoF5jGe+wH0PlodP9Tv8AEbprtatedoMlxByFDb
DY6sb+MGPQAfPIQSqoUBgLaof0mu5dCR+trVT8ARvrqPsuxuyKZSW7oDVinZciTWfYl8IhNl+KOx
0Kn/C6vH/U5x4rdXQ6bFRggoIMRRDwBqmWTAXUAgY2Z0wk855+5xFUI85QdZ5xskV1Kgb5DN5seU
jBtB/QBrjDCcQAFWrnR8iGxbSLT/Fu8BzS5bS+gg3RSFGh+YCyTc9ZGDTx7t/97CljZZkVwVwI8r
CNO1hB9qgxNFFZqJowZaIcclmajhUCrhPHKVCTw5rYbUJq1zfeu3NsyuQRCDmd5FzemIbxyZC6E3
ojp+jDVCVFpD5ynaNwHZAQ3xUcc29tM/LVX4EGPeVtxg5pKwsOA9lzRiJ5HqNYnbF7ItcTba1HwN
pwkXmDhtIr4rV+ZHXvlVyHozcHEouRSltBbhr/ys778/TF7GSgXuqVE5uDsvJL0vpGar8AVtzM//
FMCfvMY9vF++I9SYyi5ANxh83d6Q7VDSJaI+OvoyHkXNktNsToD/dolk/LAsslRMwB4GqebGLi0y
CP8yD87+mI1U+f6zYMmPyh3tQTwJmNQYg5tHt0brmEkWv7DrQqIEpMlzZ741BMYXo6+AcXqpbF9J
ExBeWv0uVC2YwNUNiPm5BZRABSMPNl+ddD6S+SpDj8wnKMzvb14YoJWcfHAUaEYCioIdDhmq0iN0
mm9HLfrKDfdldaRwHWZivmtofMKmX/uPYLNbj8IcIEp6Wg2umpY/WJiZocHxk8ncJZKENmlTEo/Z
0ziz+fpLi7Nhvm1zUBPjanvoTwwJTwn7rlXBdQHsOvyiVGGNjTPnfi7D/jZBgQGdMsdBSCXYW9Vi
iOEbyIOiFC3umV78rmNbdcEUYwKPL/OYRjhVP2vUaX5BR88vH1xy6eCh52hPjdrn6VoVSsMrOmfc
Dw1dN9Bc2Xrtsli4WaEaS2AqGh5QVkP70Rb5C6XM82thUvZqelCFXXOF9TIdTBKtdG5V3eOz08DX
gGVI8rjyBTFAllArWXLIKd/LDYNE4oke52Mc56od5gcctDhfRKaQU79a2+XHYwFgQw2aCa/8Y0cV
pA5c2ZPkgVhSTJqVOzIHmEQekZGMOaZEdjtqbBS4oKqdcNHQQbUnYabXONA89Hp/b0N4B6vFtNIt
d/rWpwVecVLy4o4AiYR+T09A3SLG0jRQwKW5E9QB6oj3nK5AehYiuoqnlXotN7gp/V0LzzaRydSp
wYpi8MiQ0nT+MvLIvZ7xxb+Gr7OvyQWbtVRi4jMxVUC+aKBfNptee/4J8Y5V8M43ZgMdATunFtN+
yrlywuKKTMXdJ78/YdOpwzBXGtFW5al+Okl7jhwHqJdHsu07CJDiIKK1jIgrECfKDB9GYT0kh0K2
BB4d0MLCM/73KlhrJRDu1piCSyg65fTvwj34X8hjZUCy+ZIJryyX+740LSXRW8at/b+0WOdseXbV
ZnulcDU1tmDPEHCRQNMZbOtePjBqJ/MY4A29eMQbktmgIRzqQbb1TWnEgzsJcU8Jim9yy19/mESF
E1Me1UzqlfAGLrwcsIZZnRFh3LWsxssEEZpC6EbC1GuWO0B2nqvbw+vkJNjGsX0xiXh1PBxopo4Z
dYZpjptMBv/bwNvtWG1oqk/tTiN+GDY0J1jimiSOQa2tlX7+s1z2woAfhd1D8MbBUIsw8qu1mc4Z
m/PYukYoQtxn9bPqfYDgCcTezBSDRoJoBqJJmcLtQ9nryyabGfyC4NrKQdrq+CFmRsmOSRhUujFy
fIcFzd9iNHz6zl1cOBaRQebza8OWzpPwsvDnKiCKBwYCffnXm/TacWLueP8iIHvzwyZ7ae/HubOT
9oe08RCVVy7bDfEUqVgZJAYJ/Ya1AHp4VsSi37Hd8RNfJJ+PA21Xi7n8vd1Ky6HpfeNMtmk8exu/
ArMzOsrkT/eF7OEpsT/BQFGqlq3vj3vpD15RklpPB82jZAKBARjo+OUe0rRMb2bL2KURDoknqUiD
m0amOH2mxyoJcWt04ZLJQaCuMeJFlz6Q8xZQ7l5EInJ+RseGS/8wD3QJkZ8G41TJ+jOa72dSkuyH
qYTmZTCeN9Xhym+KgkwPTeddA+oaGj3FacMkcFWu8P86dhJqTHXriiixcITfC4vIgxgbgSU14Hve
4HmpCObJD7fUcBTxaW8PIiwvhsbfM4TNi2K2ysAjX/kJIb5DVYqjIzRFB+odE31PWd3EwNEIwKfC
uzUeDgGLWstlBnuoOnsZuluRfSNRlKKpUDzhPXXLmZqrS+LXo0rbIKFAPiDHSzhHejSFSNhbKCD8
CZAWnUEk8yTxr7nyEC+gGA5V/dG3ZPjZzjcsBdKIOlZJzyxeijiHIcaPZRU33TIwEdEpxVQC7+4i
EW/xcP/hFN0fgAF7oyowx2VtySir+Gh38ldM2vm4wugIkVDlyYdGRn2UvzmKVTiXbT2BtnPjBrcU
Le5DUlqXOKL/fCBtt+brD4Oww6xJdd4i4Xjh7Ft5WVoUaagC27y3e9J9luvCvSYOMEVoAyhfZlSg
QhuAxw79frEQLn9QmP35eyvCpXQAi4j5nNT+dHozK1Mq71lmFm/2v7GpHC7N2Zxs85h0zgEeK2ks
RlVAb0I9EGY3ysG9DzgWn1BAnXJIhDOHw+ujpGplWDIGRXlG32IrlTDCo6U3jzG/gZXSM7twPQ8k
DzNbW0Y1lHZadA6l+7aXaLrr1Y5dSt0iDLzfG1rY7Q/jnCSqr0e8S+89PpygQTP0v7oYCozz9s8Z
1GGmlW+3aIm3UuplNRTHPSLtGGGdq1BYstjh7WXeQtrgAKT47Gi8xygjPvY4xqIIcPvkEMz79Ws2
WrHb0968X6vxmnsBuXiWf3fLjlih1hxgI536nUOZl6mye07GYeqEs3xq/N/USXfva5I9lL9FOQBE
Qa4YEx3YqXWjMOI2N7WgUF5+1sdql3C2hJowIlj7KLl+scxj/ezCK8E6H2WCUU9cICEbdSAFrePN
Zv7RNaJLFCBq0Y519OksMyppGYK69gCNyQnJNLfQhc54itLrhmJReNWyIdJQQamnHpQ7A6KiCoSw
7mDeOqiAp/xlZxBnYtI3zLZ6Sk+KsZUjNjp8PqqNVRH0Daaxbtj3pLv5Y+7HaScTlwHGzu+WMUW6
PiZTmKCHlp5vA/ceyvJz+aESxCxHrb2GH3M73MBWM6/MwjKc/up0CkpVGC7rprItZf1NHI5xaHiY
ipelvEFxSXDSWbWSRWLAT04oqDTwiTvto/42vikknqSNVxergd8LTELsdBPvj5QK+DEgL7kDf2B4
w6Avyq/wuAaH/FVlWQVmv5r8TOHk3iUgBH8yxww4Z2LVLknPffYZWXxf6ZdkOdaoolawvKRcRQwt
80mbSHvqO4S5DfMDo1GDXVHWibqYPQgOWuDechyv7elCVMevvW1JMre7TIc/fWwiCICwYmiM3s+U
Cy9oekK8pAL9YWylueMk2rrfHWJmiM6ogjQ/ZEcV5V0cgEnubpMHI+E5IVeGFA+oRk6gUXjrNjkA
FZltKt/roaXljzLEMVfOPIcX02qjOs09FdvqVzLlZp9DqBn5QDd5BTzswp/vqDnR0AN5Uhz4LILh
4AJpmQYnym+8hxyrCwmIk8G+nsGJxWsW5mNnXltd61jtwavAKVqTsTKGGjrbWLy1wZaieBz/9ZiY
X2HccfBobjbwQe/mwi3Nm0Eb2y5CDIxppTihGBxcCZdoV5PgOnpcr31vmnx5KeiMK/oSch5z4V2E
FjSLiPRk0gycnMj0gAhOSn3HUG3sKZrdZDVSwPka3QpKETqvuP5bQja8YW6pBQM+r9SNNDldRaEH
8kgY0ZPyfaLGCAAbsBOjisOalpPGG/7tY4Mth1HD7waGyUC+JDRVv0ZRxoKvzxyckCsc7/HRm1P8
kSdlR2QVdx8lYYKjwLZjB35MX9r49c1Qpyr5YbNTRbvkFZvFzSLNbNbPPa2QwU+e0ozbyWjoZeCs
KAJtLOPEPYCdzldPndKfIQxeyX3IPpOOc2zR+yVlj/R5kudTWD3j1NbHdodWPdeR+6AtDPc4/01C
d2QjOz3nxoN7ZcbqJeTkA9zXj/97UN2MU+foMPxXzHBF02cm+0Pj+mDpT9HcUV1gpCi2RF5U8pBU
M5wF0Gl3wf0TW0L4Arhb8ux+35s4YxrmoN7SkEDpIKZLGMgQ5sZdEmtzQvOI6bgXs1ZC5VBReTjl
sQTb1ClTS6oMCG1fC6Nyve+oktOwa/jZ8zT24/+rkKEaIArFBgAmwPrE7Mi+M6Ko6x2XEKowAM1h
8k7Gu2FEl67qJnGNboo4p+m2Z3Oo4xDdeJOcp7z1h++AAHk7DZwNDWctJgQF0xlXH/NMT43f5aOu
8WlZbOvgVXzLPlxyr0LjCBNsxXh5j3b+xK44UZe4J9p5r2rxOLQ3367UDPFotYmrV5FREZ+5qNet
TZkyeFfs2T0Cpz1iIJ1UkxPZCqtS4UjjuGyqTl2o5s7kMhimieAAMx3l1T/UNmVSLlOdu3/3BQyv
jXqcrVUpckPW9jD6kOnwo9u7Rlbh0kREe2VelR2ddWdoCZSfTYBL4pSZs8jkFzXZQbyTJ4H52PRK
TS31Qn2Pct+mxqNIcP6IDnzXyshQ0th7bkNI59ROBWd7rlGlfZ6alOYEo8YdzmDO+soIQ0gJMbVD
o5gPTRjd8DWbQYth78kPnPObF+R0ki+/O8eOrOIXgz7f45+mfOoLeZRBfP3EIAUDlVEhM/+UJeUw
XLpv9leSbGj3UQFviQVKggMl+2NocMz2O3rEv7iUyzF4z40AFron21hnn2qdKseu3zAmddpJfvSj
HmE9lrXdmyNl1IC/CL/zPYnpxur1GwcCnVRWc1XIkAdJJLB8KirsmWUNNSMZbwM5jFjGNqjF0OSu
mJk5A5Np/WbnwZf4fUGUrE+LpcQYy8nYSv4bWf2/x6mXQPEA97BzBcezHg8/oqzZif94B13mLyx/
56IEiuDai3k3hhKYK7BU91JD6SAVGJZ5VfT+C74hIjPHhJGZdwXR2HB8E3NjYno6YS60zmBn/syv
DFgx0VWL1ajFrn+hBJX9x+Oey1xMz7vyHcV9+TU15OeQokXAUfBRBX+VDF5MB9HM0ADm51ae0AWW
Q+If+nLOUrkgPT4VGlV/HV+7U6N9RaVLcyKTJghRG1ONuaQXCCEoAfeMjpm9K7FnrtwFnCFjksge
GVyFJckK7tpu/ecy1fqh7rXnGx7s9DzMVYAg8YEA0SaBb2PCoimZZ7qiUDL67xuwWPBCNdlM1g30
7Reo2j85GawRIFoYzUvYy/ftcW8pd5sI4Sg4QyGtxVf1BcdIr2bFhofNQ2W+i0TiZgxvNs8FvLT3
yqAGAfGN+XGIZOnRlKr/fG3RdBy+QKPke7P5FFFOSqzflVtWojdmU5kT/4ZYsDuBwk/+TJQJJDwD
TZtQu9x14RT6IcMGnpFOZYD9GjnJz6JprSCOMFgJ3KFfLnREalSJ3gtD4HHsaBn40BiYgHMHvlQx
euw35Z+biY70sVgMDX/1Dx3HynmQaSViqCsoyia66IJOThbvaqZ8dYQDR+5qu161SvzkIuMfbqIq
yz9u3mmkTfv5NoLHlNwXHg44BNoQzuet1M0InQka5qiFpkZsVt8LM+yGwFHQ24i/04t83sD445sz
mfMFyvqxaYo3HLmWIjFSm6iC+ODvhruiq1Ass/Ydkuz15cl+3JBW8i3V2DaarE47ub9h7PH0HHmE
8DvXX1/UAarddLUQZaTYqqrjNgdNVW6ZeR61xu9eOZyBS4tMZ4z0qiw1MDe0jmeQnUhyExpUVYwD
3b6NyIOPDjZVMONVYAfFai/Qdh3IuOCF9QIN4JKhmD+gRF7FPyIBiyk7tROHHIKSBSdgikQ/ebOs
pEdf4xeedFZKkaO2dpXwCvr693fmJ1AkY9L4VVsSRGVtkeOfyV1VwM5ePJzoxjljELN8+QShVsb9
EIDK1MwWevJC2m8KWBueP1nDWMBV3fcWoARu0zMPJzRpxPu70ZxMsuTO8bXT0dPSd2JjFuabBMxd
pxgDddjtb9j0Y4sYEh7K0rQE2KjHNMZd8BlZfySfsN2QTHgiH7QZAIpYbpFu1xpnchP0zk0GHgHm
OXe09wjEmhSU6oBiRlH0M4sagrSdPPsTXmsDcCJ8WhuL+BkapHnxDnvJS8iZ/9nM1Y3LT3tbQoqX
XYLSrLDZHOMjcFFa79DUGmRSgwcwJ+9tZBBYYPeTobidv3SF5imTZ/4ds/9xDniWVLXAj0NjnZhU
eNCGL7xBwpbeQZXgOD7/sc6vOfH+XsZ9zke/G7qhNUYZjsFsqd0plT3nd+U0wrkUw1yMM3eDVEqc
zZixDpW43BYSXRRLSbre6xKQpdsmp2MUP+jL6wVQG8C5OAtjI07QDLGvPLCQyQsm3jmqhI/zXmNn
NEnmja37Sgbx5X3EuVpxBvfT1FRvCAFuejD1Oz7IQeZfHhf2Zr1z7R9yNDQBoArRQ0ft8Fr1auME
mpBupPfQCYp3WN1Lh9VGtYRyR56687XLXWvNZEEdgyME1hasWi4zcPeFOLrlPtbvLto9B1bB8AUL
e5KJvmOWC3PKHua7IrKg5ZgYx9M1n0AIQFcqzEuk7Dvh08Qv6IETFJQOWZSpdc0qEKyacKuck4sb
0TZ3kXOr1W/72HcrCPAGgkDMYBG0Lfj6X0Gq/lcnQiJL01DRpYUIOE1iwx6sN87Tc5Fxs1+pyo28
DjQX4pJh2c7GrvaEXxZk2w5wJJr1/LpYU67ydu7ZmyaOvLDnqfN4i4BeRBbdEHPVeDsbNp2gPe01
9IRVBADFIhPxYwasLGd0ExdqmK2FVifLEdkUGOm4yMncRsnPGWCOtyYFunFOPMO5aXdDDyf8Pb4N
iLj0Ju01h03BzGi13O23XhKGc4AhGhdBpug3Q0lxiLIl8CdbTLTD/USZp/vd9iMYQlErMt1p4oXA
hLINe6HpJksbRAeoAYIxi6cAk/GfjRQQHaWk+WaniAbGhUeLtlb0fb+gqY/35LOxkBhNaVwYXAfw
lJ9xPrnbH4yOYyE6W8Dn7VKU4iEW796rKsxiRhz6/tpYQeCZ5cLCWSQdGbmoCPqT1LZDDhHnhAIZ
qPl4jTyI9Ce5u3PskG4LIjpcC5eIpjYmUQR+9wc6s27cLBMrjl9NCSaP86Z5FziP2r8x32wm306d
LPdRiKkErf+LcJPyPHYNsKL62TNyBd2kj8/6UY0lmW6Dy3D6epJgYo94+OA2j+NTLA1ex4Ca+1Jb
B9Mu1ws4wcjV0JZS2iyYGzoRyQheC6RdYrN+qnwsK9VQBJ0KMAu0zNY2FKAqlAhZnBEXcDjWvSbk
ZSCYcHdkf9HoGyaCEGBIt33BujE3AM/WMsohxmbvnr967D/ftJMY/k8Y3EhFddLPYTLgF2QRoQUC
lhhX/+iDgh8Hm4YfllfdCg1eqTOe6Ef6Z/9ItC9tvqnWUpKmgwooU6KvQTVyKuJ9bSsdcFF375kI
trIFXtnmSGe2hVcCYdwuT/FIwNMiMvd6kjFkUQqvLFbZTknx0SRQY4VuX6iFECLUAJppyH2wOJkL
OZWrlcVRx6y7dSSbM3q8+xvQ19figEGxwDO9LrNY4FTIp0kp2OK116ff/ct2/hXWuoZDxqMdsW8x
DAKoLQD9OvGQPTR6jOzXi3hHbqObBsEDaTZmzyEVV9WM8c+DfWVUlvnADq5GinN13PWUA3Msdxcw
GBQil3aJk8QddocSPu1fK5xNMowfjQkcURWBqYTaWh3VHjUuPSSgB/yfuUTEtqX4cVXjKdzbtFtO
8nzebhYmSwEiJCrHbM7gtt5nARWMqQebB6sVs8mAjnSej2Q5kNj5cwvcrqOLuYYJGeh9oJM2/6ji
xkJmArDlc1Z64MYIUdCFIa1vv3D+/KtPDP39LXSRHBHJIwFCVaC7kL9Z1vpcPrfc9hKiI0+ta0NK
pDr5gtAuOs82kluhyjO5kBbTyZojJ3x8+FuNMNE47kyziI/ecASGsHDlEqYGfQvvGb3VWTGKWoH6
TLP9Kbjs+7eQztoAuwXSXdt0evyQjoObi7BGzAR1frPyRkGQLE02nqu7JvNeUo4fmE1TYqX+HJZn
W6xgpN4kxT4D4sWwYdILAxRG7pJ/iV+hVTpEG3J7N0btu2zC2wITRqCBhnOt6iY54aHNLALrIB3G
8Rw0NWbqbZfz8VrNJiEuLMxkQBbPvMG38bWGB2uSvzAwWinGN0ABdlptO8VHY524dV3bcTGKmlW6
zRMmX24jCHHszC/EdHvhcybr2qPq7pD7fevKlKYXCXzhUozbevv6panTlmmTcstwVXtBNJUo+6ka
+z6tQmBwCjwAlRJw5uCZEDU2WpdOY5WNPoiNRv8X2M2Zbu8YwyswngcPYu9pUBipI88kkTEEfkUQ
zpiZnzK8W0+p0hMpMb7dKpJpwyahWlK2pQDW1upepHfQQDiMX37nFvSauNXOw7m0eX+84k/6kYKs
T5zcjNBRP2udxVfM7o+Pa+SMMAJG+9OVm0VSxX924dUeYMNvGFVCgyAujJOKp60Zk4K/ia3j/Fsv
+N2Qa6cgD3277FsqY6hiNJwDCJPeH19ZY12hpnp7vCPfl7747hz/iVb2NDyW9n3hm+XaQa1CwGEh
sKeu6P9PV8HHrrFrvjt/3W+8YzW1PIVna/OAmq5h9eJcLLlrZRHQPk5/IBj8i4gneYyIcjCKKEac
jijFU62OHzAqHtx3xdxDwCi6yv/4FWRA0/bagJrASACLlpJBe9h81bzNqTptyOpyk1O/JdT3Ns+P
/D7+EVdgEBUoSf1PUV+SgHPiPCSuxREfMvAT76Hro+XeJJuHPD/S0bq6PXvJWWzZGF5iimqRIGvJ
glOy4FsEJRSfLHmpTRHcBEYTOCya9n5Hsgz+vKyrWX7aS9DlwqyJiuOiIqYL16hRAe3Ztts4/v5+
DVqHCQ7wa1fM/3DpOrUjRKb77jdvW1mCbn6fZuKedE9KTheaTJUIh3sIYRZrxK+M6fQ2qIcGqf5f
/+FpWBaMdBPaFcaGwgUWU3yrU2+2aV2dJfv554Gf6Y2eu1/PuRX6XTVfQ+WapWHa5rAyqnwcn1A3
W8Rbe8oSQQW4F50XX81z8Oe84m/Bc72amjvuSExayyqThmmnwuk56gLZ+aRjW17CZvlQcbIBqXep
U9HO76KvP4TjUhNzmdN4SgxV1n4eRwBFDT3wFD8SP4rcsHYsp6pMpCxpw5tWv3RdopIWJgyJ9T5L
9aywq3qbBihRN4GZzgkOYGT4jQCCabXKIyvMCCwvNSBGG5f6lf/aWfBDtWmDdbPDGeJkecZu3oi2
uLPAVMq7TOL5jMIY9L7DwPNewUlJqru2OdsYW8bmyysn5g9MfDXc0EWLTeYYeUCZB1eTo764+iXW
OPjz6I1vjw4PGqSUx5Xix0qcaNEw7yusGQiUpllY+3qUMnB2C5y0l4g4Pz1hwG7OXOegMe0Hrbis
rSGyRSjVdePJHXqFzbf9E8uEfVXEAQFi3kItUG9xgXdL0zRLnkxuy+LNI158SuM0vVyiGuRrZo8l
SwjfbT37jaNsSwl85g9d8rLKyp/x+wbbJBjaxKiiuocG4EtttLEkvk5NDlBpduf7JZRqoa+FqcF3
wZeW4nEIujP4lkO2b9eANqcPhZDGsdsHjUyRPNd6hvJPiNq82dvCQn8V3FTSXSjzNSzZuYCzGoah
nY8VXM5faTJTEqrjRwlRMFrFWbqkL6o6Ay0x40VLnCwBadCQF/4tjOqFsWRqATv/MGjnrZfO1o9y
Q1OaziL8vAeyBqSqCfRnNTPB1OAvhGOO7p9n6ttoeJREmkpFi/buoU0EQCYHb8Uz9tQvkwk21MZl
nxZWo0wHQ3epnQzb7OGBX+kaOW38Uz7YqFwOhcrYiksXBDsa3EDyVMPwAUf6IRKCzJXYdIel8e1/
dv+GXFfA9uq7k5T4JqRGPiJrI2/rAxlMDAxAaHeZ0Zx1qtrbSs/zFq7zbp3ivWn9mjgM/yOZ5gzc
kf0lGpPglpmQAnDRsANpfsFAiCsKG/V66WS34VDTGrfG2LZQUsb6Mj48UlvWQXjG40JYw+jbIatK
qw3HzSH5stnOGYzLpsPwGnxwfWVTid6fq7oA5B3qgm7DvFOzraUs7/ELXZAgwJHY+4Hfe2AY6kO4
uiQn6rMHllVl+WCBeCjRviSsbkJIwnVdgmaGNZTvYgGq2Na6OLOPHRJJXS4AxWBqmF6Jd+7W8mkm
BgIf9eXxcgi+Vp9Wjd7N4HPKu2Hqk5lc0pZg8u5Yh4ldV6pKNMJMWpLcRZ5+Ve/e0niheMiqTFhF
RrNXeqTbqFbQ9fNR9Gj+ll02YzZubMNd8KO7DvBWNi2mtn1/qgIIK4PLL4rOp8m51Ji80QN5ksMk
yS7dt2AKtEJF3t5bw+yO2bhchSJg+JO+zEGSnxa0Oi7+LuklcWPF26ExSG8bRzQVkwourOks3Ykf
ZLwZC1g95qcluhU9nReTUo5vJ7GNjpGSE8MK4pquRo54mf6kLs0QKdjeiYJXaJpm/GHAWU8pvHpB
LlmGddUi6IYwoKmRakWYmvrKgeAPfZBE5stoobSpMYOkJd/r43JjV02silPLYhFcjFuCSWd1BD6w
ADkQIp3QC0ddmuDwKA2dxMVMcJ9M+OY9WT9k7BNr5Hk0N8AjmsJjSNTkdoPnz509oTPmrAdthEHx
qAQwny2xwGTPOVMBL+w6izBo6TRauA4WeDMWfaFdhO/S3IZGpV0AQwSrqOgBl5DzIgHOnFRC7Hhd
Z1Koz8UDf0dPvScuxG6nZ9Ra9Uu33/L01+I1HGsakp0mVBr9S7y3h7IsNeMpcxSb2VRV/ZaSi6Wj
xRFNrYk6+rgUy+Z8P9vG6LgbPMC13YYvsnmpEKIkGex+zzP1+7XUgRvs15cSN4JWDurIkKLwrLJD
0Da8Izg75C81RjjfFWA+K9Y3T7JdEZ2aT2pz21O/DJuy3B62xRFPkProZhgj+dD/gtGHVoOfKUiE
bypqD5WovBlPcr/NTrO9VW4qfFinGVwvBkjrXsQ030MZgI1YRXnFjtdEZzmfp6dQ6Jefsd37byMd
PIKnLART02Q08rulDezIInzgQgEEA1yPrHaaW8Aky4hrFOCDchF0XQ+8BhUBACjkr/+S/6HkfQ6Y
57ht5YkTPM6fsYSAQeJYFGbfOTq3fbT6+etkOdfxToxaZ9S6GXaAqC+FhWm5xGmXULkgTMsnYLVa
aTfEmlFiQr9IjZtPy2xDHTK2LL2t8CLwmRlipXBz3R4TFrOlD4LwR1fhfQG0c8hY3DfpB4YIWKPb
rLzcuHpYBfTqRxV0WguZmn9YqzKp0gz7iB82je7xmXNQSOUwEvInXtEBN6Vf56AzIRjInL8rPcmr
kYDP9I7yxkhOLFK2NUKko0/gGuZ4oniKcTbFGZ0lf4LzVgBjg8VC0aF+Gop0geTZUKfg6JRr/go1
ZF5AL+rJIySN3Q0uV03icsqxPji7fhDNd+zJ1z8NC7zjqT7xFZpKnul9rf6Om+BiAPzPWNR8unaB
tWYrVDR2SA1Z2kARix4IMaWgtbi/KNt3juw46baeJrX6GPe4RGrn/IsE6nt/O/QvgRE8PMwiyC9a
XRTvwKxeSZc4XeMctif1HcYKQvACdUhkHhAPiVKAt6VO90YhVInciZxTCA4rfmhUzvBxi9IkM3Y1
ij0CWXiTS/QNZS/TVgVxKXK5YHsOIi9/4B1a78gFuZkbK41n3gGLXPSiy4ed7udWFUGdaBhq0n02
o7UvYzNHvHiIhBtnyJYaIbGCqWt1Ax6IFPiIRoQZrsxBGbLB6lY+iERxtxB7E/4ug5JiMpc0wzZ6
7XUfwMuoVYTIfzsH91VZtBVFXIdCxNJYwT0OojjYjVjHuI8Wl98+O6AZ4MEusKhvOIlmSuAiHCMO
953rKBcxJqXf+eJ0/wRTfEO+2H2xU2k3ik1+r27pakUEc1iNDJozvSKhmoW2HxCES89XaLrPB0CK
WjOs/i/FY7KdRDBBvtAQbL38G48U9JJmClXcko6xwh6nLet+8anLh9iJAX0DFWbzUGcp5sl5VJaS
cFzeR3XHcLhhYAr8bUn/PHZTS9sEgKE+qoIpCOOYhcga1NpH4tVLhwNm2QgaRZQgzRiYxQLekKCW
1HgXxAnVMeFIQppbumElGIcmaSrCRnDMKc2QSXEOiOgR94mQkSlui33IE5mIHs76yH9IkdPXDl0s
kC/P1IkbbvPpMUnu5JYSxn6S/WD++sy6drdF1n+iyxnGi+R4cwV8m7kKqJLvMbIiNBLfv2jfgOfA
d5Dn/NdwmhX9JJEEOlyeQIsvwhWa8HF32QWvd2196onvQiGLYZroBJ5UICT4XaOUVxiQoVlR//G5
sfI5v9q4iPy2ZVaYhAnorvoQ1N3kkT7XMkR9LTpHnWNeeDmy9trSrmK5zn6JrFRtTBfrJnxelBex
Bgg3RfHYhjWjaABWQCHyI0epgBrYaRT7qqnNFzyjPARZFHpeVOLzCN8E+jnDF1w4gFCOQOHTXAUU
PFbGtFmg+FTAQUdtk4CB7cVqfd93GUyMgmVHgtrShJMdhyEQO7aye8tCR31laRVgbZ8usJJ4vjpz
/2+ZfGCmZc4LZw3m6PwOrJGItlEa4qFV17En3kcLPF/4jT53FJrEO8xA678QjuEyZxkE7YH5e1yd
Tfyv6WhBVe3oLO4wgwhn+riMD1Hw6KcfRFv8W42Svb+pc/N2DqyQeaFt9NQJbmgZ/1b7VIIO6WhX
UXeoX6UdNDzdUqNfLKpcEWqlnXkLFlyL3oYFtCDqkRcuM/OPuGBe9rwNekJiERmHAdtgjiyiw7X2
I821sro1cxxecv4QFzzuDgcViAZuLEOOJn+fgTegcrmSefguRU5QyQDV91hLPgjeDl5rQ59aJ+6Z
RDan9DV3MP+Rbtf75DaogCuLAAeVNcJtqETeAcdUgeLR+n2J423UMgLxrEPkjs3fK/jfSLYvae07
jV1ympp5mUwiD5ZO4an4YrI5Jj8ssFhvR01HhqB1szO0buGxCoqnQuB2M8L7/QbQxZliEc08J5NW
ePg4l76k2fF2ybGp0D23lnNF/xaRh1BvhPosFRw2fuzdjgfhuwoEBvVBxNfW/WngFBQ/UsrzcrqG
Zn+RY2ybsBLw1VTzFe9dyurX1+8ostFeaQAYIRUjHV24Je73PjF6R/P0YLZzi3iZfYVz4y+bAVP0
hknGWsYkwyofJjbqbvnTJB53b4/L4CIwOyz8OT1nF7m2Sd9wniCu0TlqLxqb7tBTs93wax2FMXTa
0bJ4N/bD/sMe3OyMgjuYZJHWA5h8UxWV2vRoLDbHIZvRi/Yv26PsSAGRpJsLkQOOfcdcIUxSD+xQ
iq/HhWBF1o+KabQDWGx0IGwZEMgOfZESKw41Ag4KyOc/nmspJj6+NFX7o6ONlQiSNgonHUtIMk4y
UdbDHGhuwOdK92fEMSBLycnlmXziepuGLnYdgyET9+w8D6UZElEDXW2wFJtQCEJ671KeOzOzSYQC
bXF2Ryig5Jrh5l5hctdJq4JoN9IqrHAF3PpkgL88Mg7zSuKXlMUnhYIrS1wddb1a78UOKLqv8hI8
yE4KE2I6Hy76+TvCW++JFpZOn2VoP5Q+4yWK8v8E3/xf2smfJ8hvTVDEHUYmnHQSW8N4Fr6MLs7b
lVFER/YH/FUUoQprC5VVoTzrFA317fi3JLaUpiCShJpP6ebfmgHA83+4MvXrVS9CMuDr8JWTjIFj
hgJpWm+sGp5OagOvGIlMHMWZTlkJFx1LRMURJ4eiY22iKAoqR+xm8epuJRGaQ3soN3CVi3uivXmu
c4LMROK5VbLqj2OMSkdpyFFg+YphBNvIFkyH2dKrcZ08t9iSPVgjqr1Q+NL/zTfxD7tIRrrNWdBG
fu29SHyNuBi2jCkq9OZpdi8G5F/ZwHgQSMiYz3aFrCdmXkEDGbIiMAkopEtnVQTV+Ej5hGsjj4M0
tfGYYrsjQxFgS24dIFhMBvgZnFZIXLhFW/Y1RD3mo/vzv4VAo8UsEaYRMxkLtj/R/T2VMNzaSmUG
bdJcCz3qQEVUEx9ZmZvQkqxRNwtVWkqj25qnIwQ/iU7VaQKX0XscLFrQ/s2VXjPzXBoSXmasp125
RRTPUOfLLQICEb0R7cnNK6MwGPAHkt9VSqEPMeB8IGE0lHQmqboOQnrSYtt7ikzSmA11WoCfJM49
RZggD6PTfAjDfVTOzJsD2tBi6HAqcbs0mQdVMTq2hJCapicT58bFR+lPHqpJhsd0xahJgXYuTetW
eYruY5eycTTykPnQisrxAOpIi+urSrPb1Ik7pBY6uBe3Tbkag1ws2/Q2UtYosOBhv7I4aR8VmSw8
wXIlDmNt57vuYarnUs5HO07GJJhpb1aPvjHo1Ieqz12wIfYGnFaN+4vmHygXNl9oDcq6/U0JacCY
G1HmGQ/Cs+Av+uHBwM/l+nNNzYmxcM0pX3693FDthQoOQasVUJyivIF29wuUTLgiTAPQJYY4VK3v
jXpTsWCDzyIR+7wZK0gvJ9p0JmopirlnI7kKvuS3Y2nl2nFdgQz3dsbLylcaKzeDCkFU/bcZ0pDx
rph+sb8vWL93O+OuICaWripSGid3/2dYUQZxCSWvoay/l9n4PCMpX5TMz0m9KLEsdVtU2GxtxFBZ
zTVNrypFlvMr8+/sc62+9ytPkVQBlXHArPcXPJIPUgLZUrj7IDO11D5FIFHXk/GnI0oVoDABRv+Y
//hfKbAeorg823ioA1gq6Mv08bwrIHSK7rT8xOkvHqohnzgtTabI7Un315smnOQHpD/EtjlIFpiI
0kI7hkuyZTc3rmlUDDmLNkB8T0LRFXtqWNzvD4wln9VivPimI40C3r667/mhjGTIU0KFspVHLhpg
aeLI1pTRIklF5F6wGax1p995r2WyrjI8blcRPOkpE4VXbhgxRFuJyg9SHhdHTUn8FCvWRSelRohK
sbm3S6Gzs3s1EcfFpq8bg6qie4GMpWR2Szh3UEhXC7stE3LHKZtSBirLu5Q6WCR1g3jUU9AqaHFE
e+NkBuilijrzI2IzNkg4rzfHVc4pnczu9P7vTQAzSj/3Rd3joLD7mOcn9pkVwJJOXhZGxKF7a+Tt
oTL3Iue6awd04yA3220mf2i4v2u2RxEKe/piIP6ou1cb25O8FPtoa09HIEJ1b/fiXr4V9/zF+aqo
1dvFrn1E8SrWGgpOQ1evWdo4i5/WnNzRlMVUaw3OwN5DDV5z2NhCCngxZzPnWX3vkC6yKSShZwdi
7NAdbi0rYNp1Es9Ks3AFXUeQvKx1uX3qmwa2rdzDLd/TTulWGXCwFvl+SpCM04yV2jxPIuVInhhJ
cgsweHG65ytCMLuTgrLOxOSOciTqHk2reSAL5Xp4JMfcL3Bk+76iEe9GyM0LMHL45fVWmeWSepUE
d89fZK4UMCAKCu0z7sNQiC5B4gN4bhbFlvA1biZLtb3FZvWF1xbMZTHkO6bZHOLrXoukC63VAxIx
+5cM5/9yfvfBybKHNq1FsQcXyGlNbopbAmB7OclflMkZadQDnuthz0fL1zFwwHj1F6Ye891cpUn3
RAyK+rii4jWdctga53G526LoTsoQT4X68EBDhyMchd+BA1jShcEYdI96IHi/myLIHfXk3dVOrSAN
CfKatCEH/gpwPDuDyDdj5iSdjVYuJhugDDf2y4LShZvGN9/Jo3vFeOOkwIprydh+CUoky5CJ+za0
IRW4JRlIOgNDpXfc190nid5EnngWd2TA8BXFyIrrURC6mUfDhNhhSg+JrARR8PCsLKHrULfPkFXh
eWItUmOhglX8QRa5q/aE5c0f7hxRSxC8rvO389CwRgSt8ZKPRFy7ngpSnD3xk6v6mb55/tj+H0k5
rfqCkzS83ce+Ne/lnQrdPCUQVk63tTNQnjBZoP9EmX4Ruh3NMGofaz3mF9VAU/wiTD+IuGdV9QwO
lIZ6DRq1eclfUHymASs8RPwxAmD30ey0JBW5AYtjGR0ncs9Cb6AwDAOZQlPEgoIHS8q1Iv/0dB7P
VRIr/bbxw0BJ7tEAoSzpIXNn+06hBLh+LNeyxOtvmmxjqnmwseFEyh3DKSRjzE05Dzw853bQNZgd
JmdB4F7WznOsNdpUidw9p2aDiCc8GWvl1F4L0MW00vU2zzxc8bUXXvW2af0RGRmuMY0wGVdWgG8s
IJFCYZtJ6QgiXRYWpumywnqoA7ACUV6V9liFmWo/+L+jTTuLeBnUKcoHYiE6ewKQzlaca7XKDMwR
XC4E4Tbm9SXW0axgSDwyTs6DylRLTRLB9u5D9gyQdtuu2JZtPgCFrc9oLjlOZ+zAc0XpOuf5eMpy
xqZBaFsEGxKCqR40Hti1fIDfStWHVu+KhC75cga+urtQosRmVKd7LRSbynahuW7gkWgqHHRNr6ld
QUQx5ptXWehp6QkQghNewhDrg54FRPR5kMtvUthMi+abF7vPAQwuu26hM0I6bCv/NSJLY7fTZgRt
F1KlXHYBoFFF35U+8oovPH1hh+AQxJaxep+xDMgg2g+LEQNPvMep/rNhgG4zdNfwXoi8TtC9EKrw
hKV1sSLdZ1Z07V0S28LeyHQPwweXmz026/a4HZN0oywdbJ7gKtRwu8TuFQl7socZKh/aJXN9D5y0
7mT/cvyO/7f76hI/VSwvgJMq4fRiZ2uMUQfSbOmjQyw+kjE4ocA3ASFs6pIfgfbIaf0T7wzYkSqB
DNRPYVK4p5XzJ1Gx49FeG6yeO+sGMldOuzgKGK3mf/K31UpMRgETpjfYWUfvFeQYg5VfMNPMjE+P
V02vtW4WhYeUNRMY53AHXcMv0cjqDZn8WM/DUIEOHCxxxmLjUhgrM1eTYrSA2edxVmqVe+oJjH9F
mNeCk6HLkF+DJcrJaVLPQxdyyHK4E8BcdXtXsYmCU3g9XjsgpDmwMD26mFM+tDkYvrNpJx9hfY4k
eyfOmiQw6i1qR4LZCv52ArpwMorqeUG8AB+MQsqTjQoIbKkhBmWWeEBEYDVxqKgAVlM+eVLZFZ44
a5yMJT2bprirNCGT4OoP1Nu9fUeCFbXsB8by24IZsQcjiDRWsl8SPJ/0K3lc2zvcaHvvskyk37gX
z1q0no89xK0G8szk5+5zlZgedXkIAzItkgxtJWpmMybCjzdKRtObKycLTE9Da50by6TX0sgjgI01
4L0o/tHWB9I4qVSOpc+Lm746XtUBg37CnZxcA8R/4Pf+GF4XEuxWbJg8lFVJfIADQ/D80uzBKMiZ
36is2SaaT7bX5cGG8THnJPbhXGP2n4S3sgfDcMURRk2NhpCnrWklLmjF65dz2rmYUiFnvW6YmMNx
iZzpmdgM1KysU/yn86iTS41EmguUAYQP6r3OtyzscHD2AT/QkwvDuYZ1+QnyRBOi0OFN2HghzdBf
CbqBwwQ9utOEjEFPtLdZsT2D3VDbpRTgN9sXMF9ubLMaTNc6PXE9gZalV5RQlmek6f9G3U8+0eSD
4kNvE+56utUAfMx0FFPhsRvMVEyUGy+LcGmpdEgQaGKFtkA7O/18IOtTjCFJAiAZuikSQesO0RBv
myTwHp4ydO07dXx6aYCR7Z4RfTjYhiFSr2TBsziXYhT5bWx6BmlzGFOP+3wg9SgNDk183TX70McF
Z13g0p8fprITYeXNijtuesBLBwppRG3y7ite3vRkzrM0yze7YzzfJ6gwpdrszhMl9WZ8qjgUIjLm
A9NBKYwJqrls//0x2Eh5jL/cdGQ977D4n9H/PZDOfgI8JZyrEH7nIHnxCOJqsmOSHXpb3qGfr9Sp
yYE4IYIeHcw3Fp+Vw/1fl5qzrw5lbnOTMRHQ8S3qc/D07TIVnZQUJAb4YW6QHpiBRvUTGt0VAX38
nScpc+Z+tVt2zzi5wlVl760QIFNCiWbjvtqHZgC3xsWab+Ex0F8BNPlV7DA73EICYCD0T2wJjG+T
PZshb51gzA6gIU5hrWeEzK9h+A64DISkbAE2ry3RaQbo8hs08msCcNG0cIy9P0OK8RzT4Bs695wJ
JGvpicnqIS6RRtdB6Eb8gwkZd5ghyREgb5fNrR1ABAVO4QMyyY0Pt/0z1SwS8o/NzKYPBM7dEDQJ
R+XxHY120ZkJeaa44dreu2Wo1U9OjXDeHVWMJPCfpBU0fsvty4LBVBItkbRmYyP4q3QtiX+G0N+i
U8nSvn3Ba3s18+Yf/ZHnsQiP7AYaJ2FXLauMJPfgbFClaOOXHBQ60HGKKw/aeWRzRDxTz7G15Ju/
ol7URZaJ1f3D3zU20Xr1GVR8YrxoaU+n4o535AHtVw3dVtX9PihSznEJip5UZMjf6AtxfVJWwxjQ
Dtj/UG71wuTgytZFMKpyP6f3kQbvZodZgkrEC+ZDGuhoHfY2jaMm/tfs3NAzLU4A2XcsLZbhk9IS
dzbJdq2xm/oxAIOkhGDYkfLY4mTbG9FifZxyhrDDUOxucljb1O3TQxDIwEJaUWTsausbrndutegL
Dd5zhMIgTR4p2UZ+WRd+I2tUh/RlYcVbP7HJMDnl+v297KetNXc4PZuOBAPPq5tps4y6sBjfwPMx
Qhtj5U9SBjvQSYCHL0dV8k+VMNjrbIL9hK8B477oO9ndeGD7RIHIvmLJqmnkLd/hFGXw1VE+KBoC
1ujxTkyL6zzI/qBkaXONKlq34K9mT0dK21/CwmQcdOInpuC3gKgLOQMPZ7/qrsy2o0IWtnbVHYzk
su6dk5O09VLz05kpCuUSmCmTpyVoJ05R1W7plrPq9YSTnR8uSpy2489W/R6W8LBIUZ5b4ow/ai6r
8VGf0YzCxqsQlLtTDH2WYYY9rp+KuY/nlj7/TzNm+laNCQNGG/vIkbuctVvBTf4+Db+4OLaMKFgY
/5n/Q2XxmNeM7FdJflXz7oq0JUVEj6MxAvFZvPzu3Yfif7vPW27MC3bSoP0ZHfvkIKp1ZFez/Jmm
BA9iIQGrg0mP5yTib9jb3Ju+uC2MBziEfLwwjr2K48idrmnKkEGGajpD7wne1Q3o4s4YJSDAFr3A
ZylNfIH/6cTmr+j6MqnMqQp6N3Xmtwf3MqkJi+I5UklWPBEXRX2ChkbIG7veXb8xXrdEaOh4Vokl
FChl0aiyp9WHuJHleUbWpladAjEa7NOZZcXaAZe7d+qXx2xVYf3+UiqwuJd2YEuHZVMuSlCjHUnE
IcI5lXb8/reQCJFyUj7TJFhRApFuNLxtcNS4y1NqUdIpWPfNHRR8Vq6He2ToST5gQwY+QdHlN3Jh
XwbcKbm7aunuERw7IzxTT+M+qlp7IaJmrwjGTp4GccliRU2xf6wSyl6xjadyHlsv8BMCka2A6oJW
m0TSFmwdgrySAxQD6UsXhrNHbXF1N/md+o5mpwSbU0w7sJCmranmoki5qHyZnOxTYXt7rVB9atcK
DL2e9Hmp/eS+viybUE2vxCHJ/5Lx4ukSUjTmd4CmaXdrgE0UMcP5MTPUL4U+7oERVEGsuBuUle2h
bEfOgF7R+R/0g4Sl4adssDSDLrN8s+eDdxFoazm7vR2hosYs3qOoj0IfK7pknS1Vsu0sAx91NkIR
zbcLBVuCUJVuGi0lHDLKBj818TIhkuVDOU4c0mWP2LU2/4bdkoLbEEAOuo2/Knl5SenrZ+uAaa5Z
c6eQTEueynpU4mi/xOhwIMEYIIOkoQdzKfH5VbBUp3sIWXkmExex5EVoI+S+RHdx2l5pBbfs2/wN
bIuror0iraAd503XY90wWrkid1XolAW28bAlRWS+MVxzSmv/Hrngxl1cQeEbsUAlTzgimntGQt31
7yDVAkB7e3QY02AThDFQ/yJfwaI68x+5/l31W9HDRPqEuZwClLWqGxzeItZ7SXonSt1WfUoGvwrZ
rF0CLeDV0zq6IsdP0orC2T6ZenrwCEr2TyokCFsw4XhA7kbhSzHgf3rmVxT+JwlKQy6I6BS6KoQU
db0mQJzmTOAua/3rj7r6M/j7IuITPBl2oycUjYKgvH7W8JcTY6vE7Sdmmqt86uhXYIUqaUwkeXFP
bG+6UF7L7LmHwegGtKzuh7nmQwXvYU8zJHYr2xYfMOS/nVCFgTlP+PZjhCBAwFugOGuTgXvBlgZy
QjO2eJVuK9bym9lE+DxXd8GkT/MuLuO84Art8+dxOG6r9GONrR3nKj1Ao5M9YEVSclDirIgZ8q50
4tAnSvA4B7xyU1dII7mJ95zyVQFvu4lfI2DwXhnCRyBPoFNmGpAfLlhKkHZib+QNxDrCfkLLfOhQ
tIpOlTeMt+2e04UE0q3KMAUosLgawfMte3HnvTrQF+2rdJZnTGayRS9AasDas8Q2RGd7ldhjOO9d
nnyNaKfyGbd/R0zOmTdOB1KeAVO/ViAbcm4gqgNgy8TDLghM/yAWtHR7JOLUraxKrGRHN9rAAwGM
zTQCPUiEGlgMtM1edA00TtCvgUPVoGVp0QYZGY+jo8G0Q9hoqrjbqSY3z/B8e0t+bGogudxXaLoU
SeCCaCpoK3WdQZyIP6g/a9dlbGLWfsc0o0suBdrSXbEahHdrI3OtOSl2GZzSpdAQRLAheN908r/0
dpEJ4UQoGXINc4uuMmafVtq75aqA4WlI71AFv+aMwj9ZBO/0KwcZIMAXJPREVeDjueqQ3iC4cdmA
8NtY4O9wrlYu3MM85nvxXfXpeGHA/SbA8CpF56zpTTkX/COL1i52uuW280EZ83pgSmBHcvU+7xOY
RMvlwNPq37IDi7ZEPxyvTN79sTK4BmI5q/0BqfDQbiLonl8+3ytP9HeizKPG0gBAmCLcKhqzNGcq
wvgGQP+aPSoFxZsKjqyNNUhKqJRs8diPLypZO6+0jcHm1w+w8PVYkHbAyrTqXu+Dr/GmjvyLLzzo
CEuiElAc5hSSlAKL/SOPB/ICj5Z6zz8G8rcgGKIJLQ84aNZoUy2i+xhq2C2pmO/ikA6vOoKSMAt+
/v0Bv4wuQOxO1984rwJSq42+s3Z7QVfYrGRoWRxQcs00WdP27YpU4DK29SgQZBpYEHrsgzEKC68I
plqgM0CxQliCOBccNQDM1EsFcy6PgUIKXbT7MMYq/M5KccJepJC65eXQnrQejl5RRUWiXxa5ahOu
msru/dt5S6zhmHyt+qQBlM/hS7ebZUhJhqtoiL5AQxrnJZjM2lZ46jUza3I4nY6xXAIPy8RHxaNr
KNe42IFn6uAcki7ASrep2//qF0JrzX3iTHINyvAvL2J/fXhWdG3Tlsy5ZiYlUqJgytAiKdnjqZP2
S/Ie+dW7faXqnDR1qbcsUADrDED93woUEBNjBc7xEXcGtvrP+iFOIo+fapws3IQP3NtwWDydeael
F/3brrt8UWo1aomIB1m36vQ3++lFRyxvJk8nNtr12VuezEMNGupXCd+GQDJFUEJ7ZBWHkZwiYJv3
bv/nZ3W8P4+7xCO8sHswyfjqKtDC/hMd6sV7SNDglxLuRM80MSDQo8yj1+wgt3NNKV09EeyVdDh2
OXDfXaa1UprK53GISAxYoFQ09tC6na4Bf7W5akUYyYGw0KRg2IlUaAJE9r0NqqsYd6i1pNrBxf+Y
7bwj8RJVYTdU7rBcy/x66U/HSfmSbvHUoKlLpMB6PYZCRTfugx1Grxt2iTYHFeJGjDb7Rc/BDg4e
dvT9u/r4th7p93P2NXdYwfcZSSSJwYE8hGV4jqIWVf0Q/YT/q8RMr63XAseKlYMxAt6C13sXswYS
PqUk87+F2yVnC0+qAk3K7HT5XG8Bc2t6oIwV/CyepeSX20gOC3NP+pPhjwE3o/BuRH9k4OT92jcZ
4/rE6T01V3bXXRlvK+5qUZ5hc8SW9HrjyjHYaChMgk3E3IE5NyizBjne+OsU7qjfgZkWrEP2Dq+5
PgqcPtpc7RbsbuzAqhpz6qsqMYBwgJoZB1gvl1SESaTS6yBp1jbsVewZh5ZTikp/UI9LnUlYBWL7
g3JnFvzlAEbxEDt8KVW4ADae3609cmB3lB63wdudCYrMfOEyw66ev6d2/6Ukg0UPNuoAmzWbSRRW
VwQDYM3YtZL1XneIhStQzi0ZvVaDPp+Ncv1fKB59aKRDlbIyEUnDgMUb84pambctjfLMjhgv2N1G
NyNAedQqj3j/b++alqW4ZUFROdZf9nHAkfik1SW5WbMKzQB745RfpDIBQH5nxfBw5UHJA/PQyJYm
Co9WYs+D4VRiYn4nPLx0aBrXZqd/FE5z5oZvlw9vZvi9b0QDj2vSM0fF9miqgKDsB0CsrzHvnigd
nGRYqMLbWFggfBc0dVL2ZfSVbW1KiBLf9UtlANfR3A2Q6WagRlMWkow7+D9VUa1DjpGsoZoMWAnv
aI5sD2H4ol+iqaqmxgXeWSJ2DruYmWCZmCWCRoZaVzTu9lHXBXI1+7OR0BvxwtMiWduTB13s2bWO
3Kb8u3Mq1PmE9rlKy0WnmKjSdAuwxkgC6CKLAPHOgO5K6Td8st+a4v7b2bZa0uhhjfkALPanZexY
PRmGRoUE5xLoyrlkwUee57WM6IPSgS943N+3F3YSbRuxKrnqbsFOPRkk0vg4wod2B0O4SqpwiSBW
gN0RewAFBHPmo2Kk9hZA7J/d8ghhciYndSGQnzgk+L5Kv3WOONLGyCNxs6KeojSek1nRI/zeoGN5
0lDc/ES74GWwDbHB7mai76rq4YSQrnSVdBj531ojiwZsALUiWRopSavWzUqDOO9iXAszZrxZs0LR
geoQXAx7QVOTrAMDQPqOKUJ2dmaOpWa7IdgWK3gXrwYRJdNdsbk90qm3WfJOwFi6fg9Zj2hltmTG
KnlTGBBKVCZfupxR8qlekidIrcVr1DQ7FXrqlCSJSf6qAuuPz6phTAuWVeWq8diY8/y2DcRI7fHl
QYcvow2rkK8R6r2StER6XaCw4QZy1W5ZpFRzA9A2UphK/GWbXmQIByGpmBaLwwTzLt0SjXNl5WqP
eFjSrblS1LaqABIEw7knoaX07HBTNr1PUuvNObyrD8l2Q89ErcfDxmPeJuwerpENsQbGXiGXBBPq
h/nAWmNfhiGD5lHKcBzxtIqL2CVlgrYR83qZen8Jugi+wZPjZu+qCuLc5iMlTfDrH1qmBUIr9R8j
V0ylnMal7xufxm4dxkFjpufcjY5jrVfV7tRLKDqhlqGrOLIwMB71YbakeFlyW7zEoCRvwulYsIb+
iReHR1RClTjh3JPY7s86dW8f9KN3r4A34XzfWmot9rklfspfh2ibeHve/+2avk3ojzZHpw0jgJ5F
5QGUPvHfnFn+Oww8TlE7DPPJm0aPvqvvkP2XdbNy90/xQWahHqf/r3voBL/gR4mLyjmrzrpF9mus
1RWGkRhxnQARTwd94PBWyBevl7Y/T8PK2X0Yc4IKaLdXlYvqA/cPcSlfMOlu4RF7OR2P3sMYfvbM
9ZS0731Z7QVnXAKSR8DE0Kd++qoN+m13wThIxBjW4aqMgJ9wpIiUQyXAWYJ7VD2x0DQ9fkjtsOlN
9WZjvjHTuiEkEpPQpDekXUh501dujGWb1zdjJmKJNByXjyRFAFtUHrB82fng4pFv33AxAd2+QCsL
a0Nm6nSo/yf+LMcM8yt531s/el5Ep2hoScRrszeVHAsc9iHgZ3fy3xybQwvc2sogF+xutB8fGaN1
yCMydW3Rp+i6VZbvVDC82j7XSu8hh67E+dd7jV2kefj64fsYwchgktaYMeg4HPXQsjJHag+hjR2C
F1M0lJPS+4jfghh+TIDSgO0RaydR48iQAoPbS213tjZ1AGZ3GbEsXgkS6qGFLqMhujXuoFM/vUZ2
hzXIoLG7UD9XGVSfFVYv0PDhRVa4CCK4Ar+QgUSBpW9r8aDQ3VVZ3h5nxqd+qWSE68P17eodv2mw
dZAmQZksLJj3N3/qAF9+cu52pjEUn45DtcuecVlZeWdYdAO4qYHUuOQ0UL80oWkHFSuNBQIir8gS
CuWAc+qr+rSCQl1ZU+djookacJqWFGzA30HevAkDDFVJPEzsUGZeJdN7cOL+dqqo27y5xGrBOAfJ
/rgyHfyCGUunzOylOuauYK6JgF1YHLYoC/2PCpTUJD7h627JKE9u113GEEyqM5DI7GdElbrRcI1S
zQUcoxK8Vkjp9ecVelGK9kOYrYVBjjdR12t5y3SvJutY92zP+zHPUpMliYbw988l9KCZbiDiZuCT
9gRyzu6oC/KG8V8vZGkd9vjUTZVtkDMEAc2OXshz3mu3NqzcQ4+w1fyDKS82WAS5ebKzMlGfGRkN
Twq8Ag3hDEi6HBxU6diiUhoXIoYEssbA7Ts9XOo3Pd4/hTXfzMiAqLL9jo5PzZdRWL1ilrx0nVA8
UKjfIKBfFevn8r6O65pFEbC3XjDb9kMDHeE3XH1ixvIR/ugI15tI/tk5WnxPDQ6d1Ok6to+SpztI
bEK1pIEIzLx1IBkmhjYnL4OyUBInzXWg1xJLsdxENf6oP2wSdDHjHcnWlSwqzYSYBAQ2ZciDDb7X
3Ai0OwPzA2O0UDB8nZOSVrFoZb8feBEq0ifn8Ue5cGARP3KIHnt+r+DnpDF8RTR5lG/CsyK5JdGX
zRfF1gnh1S4kCQ06EdmP5dvdJhxcemqcy7uHBvn/LVfttMK1XRTxtulwqvJZ1GvNDjtHXf3z4itm
91Y7P8/jznEo3PgvnHC7UXVN82zwcMA9De21AaSf74Qwe7UHLN0pnEqiSv/06mfTfpyHSQpCqi0G
vX7hzuSQ9glHgiFVoXAKcXbNZYeF/E5DMoQjVHqgX3oAEs34WTWd3sASdNPVKxy+RD9Gg0MFNPBs
F2BH3SPoUMwJswo/+HWnCFmegHEb5+TEh/m/phZSgVw2+2FEqodJc9E/HW2h+l5WXYft0r1/BbbL
mlUCMX/hdZ2YCBZ54FXrRM+QnW1F7PiPVZZfADfs94WD8tn74tMuPqMxFhSsQI8MlZryulXu765H
MRTFDTceh2CUXTuhQR0rehWIFP3y8+ZC8zFB//udvB3zECKGuivOdBxwfLBmjLwiwHNjnZHTRvQM
izVxWeVoeGYyST/uUpNdR9qb1GXBnPUmPPvYSmmSsOt92GWPfi99tpJGp+B752zgT/vo+/11h+e9
YBqWvaym0AqrNsqWAZovevV+bgbpBSyXhY9YYQZqvHAOIYIq+hfe847opPs5Ox3MMHreRsVEeJi/
m5RWrOx5kCKsjrnB+XREUKbxPHIy5deVuAoHQCD6YeZlX+3VjIi+b0XwWKoid+BWA8ddvlB2Fn/p
z4uKGlIdC6PA8YSLx0hdaLehjgeSD4pfCiisBQxHXDOlHuQ9iDjA7HOExcRdJQN4H2HUCEuXDKoQ
TXkczRLq4gr1tNm1afeaqRDhxHWkJXcmNCXk48uK0a19uaI6s2nG+UEE3Bhy623iXBwPcA2+WXP/
ASx8VM2rqNfdKfxYm+NPRrBtYfZi9IP5cOuKaswJVTJWZTtuIqZvnUujp2HBWtTVYlNGfqgF05ys
xhCAOx7QpMtoiZLI4w9KzoE2h9zDwtbI5OSciDzH7A9kQeSzUsyhpzAyFsDMyrTmVaBCUkSXN0I8
IqCQAx7CFWRJ+4eCHXu1v5BIVt+DmVcaAwevDM5KYiMxAsEaDt+ncN0+CB3jYND7ijWrkYtku0Kd
H1c7EvOBm/dSOg01w2wgy4GBHAtSmTh9rA6P3lE/iccTsJZfKI1d030sCTf64KMmgYDz1IGVp2ji
7HbUkaYWsV7+cqvctJgeLDltRyDqORo+eKWs7U+Lu8xyew4oReOCEVdpXjO7p+F7teFAz0lNR+S1
qmF7gYYHQqHmh5C9bg3xkRxZKlbMNLJmKYgarjhVLn1hLaQg5vRxkRE28lcJrrkjBQ2qV1HMNCIv
lpaKMMd7m9UOE3rZGxu+x6y4nzJvh2LOVd72F/1jojyKyK6a0res999qnwjbIaJ8wsGvsOQr31su
hxfvcs2uh4sClwVRVksjtgDo0sygkv6MG6XbOjbtD6tMGg0ZnSt/M3MUvY17vZMhj024DihEvlo1
3sw92QOnUNpno3DzD9O5O33SY4FrxmtV/f8z5oQRZHc73jM6CXBIJwD3f0+Z0gtHFsWzsmbQoJBx
nD+QoOlU7Hd4kJnnGz7uESw0c3a5N70iM7Z7upUWx8rBxBtI2I535FsbIPPlgHW1kMca1mKTQ5lK
xc54Izms5DihN9G0m+xV5fCs0LvmfZGGQ/eMbfPzB8zRykMLSnu8i7jn1HeVLnlnwZYarLTJg4Ar
e0YOeGDCkxtfi96mW/CtJPeVpKehDGeGljneb1exQ0KEfvuU6dViHLyCUzyl5sQEIbaO5gBGbjQ/
IllMmzMdDqdsrXqxukE3PhJ02Fkg6je8Lr9qEWsPzmUUNyENBNnZZARvDjoWPBZeHSXOTkQubk98
2fvkDZw6MJkW1BFcaCepmxz+Wcd7fZkU+odFiwMLUhg5Y7t0ZiPDUi5N8WvQeBN5CpmPZSoY/BC8
5UMw5cxukm4iQ08dAkCUDcCUjfU8/E1rHqyZ8V7Qtxcd7y6F48akBu4LtNx7t6UAMsQEqm/pFEn2
URRPamTWze+0xltiAVoVOr4L7UU3YKe3FW+qhQ5aLkeClq1AIjdZNjCbfKOK9L+cRK27LDo9kaBU
IHtDnKMSl+HwRGCONdnNx1GjaA7LADB9E0LI2WBBNfFrRJZi5mJOsOhDjh27ojsq5Vp9d5uXSaiF
2SHL/HLd525BDyM9kOJl/sJz0gnYprdtkqlyntJIDrpoU5vIYMlk4PpYOjBCUnKwZocfZCVjxC0M
s2Y4CfVqfWiVZLSTZl+57uziYKzR6RkJ4ft7cWXfe/GZq5/KnKB63YOUf+SCBx9XYhVfVLPWOJIu
Xm5P3n4J9qOK4P7m/K07CAnMIGwD/FBphBap4tlfMfS4WEDITW0nFOejBb5YUhGUSyT3uQlHKy8J
2oVeyTWF9Xb2YT98pF36mijbH92OxIlN8lSy/J5P2dfioFSOcHh69A5NDAKr//J1ycRltoMwjhdQ
vbKthpS6I1g2v++YXrZq5X8luvs5MuIjy9bewT79ovSlM3bEdav6moGXXrSizzvsUw1SO9tXVYps
FaF3jRsuMuQg/JAUa7X9hnIkUYQ6W2aYTTgVIFN+rhVupkH99+1Pe7uDN/hCjN8AaGe93+l8a2dZ
gHiiVIBOrEm0/smxaq4WxztRkvF7N2CR9VcPzR3j/SmhQuhPusPB/0MdinCQSsKD0aCHgXShT1+l
FHI4p8B5k5qBqAF2N/s+efMBljAv9+pew+roLhshDHHcU0xj1GzRWX9pUXZfErNWalPe977EDRHw
bukeUI9sX77ELzRnULFLSNzzD5PSh5uPZbPOwj+mk87y2jYX6VbzU591x2VmJ2lddXjH0kQB8jqv
hplkvXOK7RNi7QqUpoN91TfUNA81ZBFgZ61nqtt+Ogh/dT1VENji9eKl200S/EpdfC0yezE1LST2
Zy/UrLJGGif0pd86nPPfPz5VWW45C2tLTXZ8EJzJuCMoiDxJgthg3WOd22auyD5/1Xj1uegysvk9
deVL2RMboDjLRz3FMexmoxJPZwONIHYtM4qu72E+/Wo+H5SmMTL2z8XzuMp15g7QYTypWitIZxEY
bInbDyvVKhXV9KZuZxtqb4ahJZss230Y1VwyDkeqBFmGGioh+hJxSKZdFjTyTFrMD/alWTpC+1VC
z0PJuOXhz3QTV5/sibWOH56UfzbY6AqADutrUuL6hSeMyxtWcEXq3c6Lm/rUSYuf/8iWM5xVQuZv
gdA4l5DGWhdso96NPblDHE8atvgiCnkAshQTDHTW3UwJ/r3T7bltPc1hVLPGCCF3NCmV9f+AArCX
ui9QFDV3EA/UpchRq/VOBiWiCObLvmlJ/DU8w/eJHetUW3gpKpKkiUYwTGTg1SLktVNPEQ1QoBP+
9oC3KvFWLdBrM9b3ARNgHEVjtptamynIN3BGqSQ2IvSwyOCWINVrMsJEc/FBaiEuWjFjgFC+azNO
kMeTECv7iPHQUN3SmOL1aMAvTPXOJtdoMjINU3X0W+tyKWyhCaU2stC5A5WYl4BjShs1j2I2MRr8
IUg53Wjok+Ey+VJ4F6VP6pWguLmIuQoayxhlRRATZgULjOzQ4nP/zJhqmFMu/fShz+lm0ARtzxiS
pdFPJ6KsYICtkAZ6unSblg1LqJD+1W659X8m+ZzdMY8pFOKnelhUk53oHwNmZFIvk30GYjoygT5J
hV+SCFot2xJWtMV55qxTysEMy0PKWKPQAw6BcaVcZRbFSdvHZkGvdhSqIRclznycdWnOvyVVO7rl
kgUXF7PE3l/f504XmBIjMY0TBMLL2tDyXLHBMzlwpVoZtxr3isEAj1w8c+W6LdkA9KOv/FeW5QQ9
j0YQTey8Tix0J0UKd4SWmn+CDeu9fgOqUlr3DBKooSlSjuOM++zVRzURAwM1PfIF45xS+jkXogGT
X4O4IAuyXdJC4iS+iBY12Oj96gD1akr35+A9RBZnJ1TtCK2aej+g9LvP6Y6U5B7lnzBeJLLgfffc
u9TYnndBeIojlhpMyUajyupjSAA7l9NK7FBo5Ydczid9KU8jAyZpegWnnCk6r+Ud1wzlL7jExqT0
GzXClwJhqjtXQO7aXwQl+AwIO45/qq2L4vViDFcc1WcOoU9skcECffb9aS5s98k83yA9FlvDhCWz
i5eYRb+2hNd61EPqoVUMdrApE7X7GZoDN0LlAufY9yL1fRwqWwGxwPQowOvXYZkUXe2IFiy0DJyN
ldz3Wb5FvakVdeNTQdY7yLxGykUHPuTRnjhx+6CbSIh7BjrA6KrKrQlqErzDoa6cw3a+8njtyv5z
0Imdgj6skvUDwbf9O/N0HwER/rP37m5Y+H2jtwMIB+LXDKm4SrQJI13c5RFlF/jGqY0xepHzpuK/
kmI9I7NU8w878qbOQU6f8SI6xV4A/lcgISQLR0uNBdP/VbkVntOd7sg0Lp3RWCC9g6jbfa4LggPq
2+7sN1wdOFkL5tdND5FWzfyQN0l2+KgPvUrwMTu58Rm7hNOvWBzk5YtC0gJY6RV0ryd1hMF23m2P
ix7UjlmxZtHdcPVNm192qLDvHDZVPq8VKRhbTbA+BLgO3HpBgMVI38dszzPIpSBh13h6OslgaC9V
Jd9WwSPpD77ZsWP+zlaMfi8wz4IbR+avH8bKn/mOdeTJa0eU42KBCg4FSWiITP4bYHQoBx/gjPPA
9cB4d85/8ozDWNtxySJzZeBxhKkythGMpHWT2s5MeuC50NNrfXDivkFFNZjvvMMkma0l1fK1i3wH
biLQ7WRhz1r4f78oRExSaC3LW4MmPn8u9k68ynpSA+L2JSXIiS4o0yINaMCZTK3MrPdv1gmbIkrm
TUNkYoMOhvHbCYYbtLqozT1SoYWUsilQqxdy2R/2+SQSpbwxEsxnzWol8kaBHJEb2Y3VkjbhGBJ2
VrWZ9oIWBv4vhoEDy6gKgTHtxq+IIt/kmMXAikvnhSSqQfvGAhDkbiZm0B/0D0LRDHk1q0NhbG9c
HgtfbCsc2SsfKPOrygdPGDqlzSkBBXFbyfFi7L12nohkxZD6/qyUA1SMQiogudY7TtVgjXW9x37+
JuuRpp7t8LuKGap9TnHSiIAis1lTc3fiP23vzdHDcOI3x511QxxLgNaAORDBMq922ly2DqAZ4nW/
j+0Bs6OqNFvEYkyh4Dps03ph2aelIQnLZUM5eL9RxJkEjwe9VICmH6c2Xx0/asLfZtliN5Zr21TU
/N4HHvsJ2/76WXI2r/f8ZzXhB261PgNidQ530VJEDiOCfapppyXkWLhjf3Jr/My291RX6NrPnpKu
tI0lS/M9mSr+qTSa9AD2DClNseac//5TGpIKJO1BOB1ozIP9yKUPjMvBC2TOhs5yOzSAggmlFBsv
QxCmeIjARRT55EmgempdL8b42lmJqEyLC3O96vVQlO0+lAP++tnomhpy71T94p+fHfuUm6rR2/IW
JIG5GvNPFgj1Dy1KPss3jqAXFZyzi2swFmQL06Kxg6/OjKYkySQLMQxQDESzX4vRDVOj7DhIaImB
exT77sHODFFLnvqwxBfIeBuEp++KVW4tv6TR+J6KMBUA5Dro/5QKcQLMsIbIDhGZ+sXMxr3+FSlT
Xxrb5qbYGmCi2ayMfuOP8SRVI6BdjL7DiDiVC50WsG2si1PsXCfRvDwhWmjz7h/aTgiPtONJKw4w
rK52sMwUgGAe3iBoYxBKCt5ntCC765AD5p2jR1ZV/JGnjS+DEl7wPFbyTgvRp2CnQAgog6XB3/td
R8VCvwAwx+1o2DLM8kua3ru+5aqIF/6fW1O+wr/8HtXiVWmtzfhlD3tW8bkI+U+bsCO3GGfU4SN9
0pkHrv/t6R2XOCkjOBqaCnceKH0CkPhWq2s6fg4fsxSlUJ2rJ0m3QqMlJe9ojrUwK5/10MoPX2Ba
6+dL3hqFhxjLGpYD8wf6gIBcxRwbt0n41SYAAclO5Jfl9I4LI6FZX6Qx4febFZLWdHa03SqZN3Q4
I+W2wmY5TW3rB/u8K/G88YK/62d3Am8UnL+fM9WS7h8HXAMLYxwN+x8/EeuvUGtfyErqvJqMg8OY
KqKtqcJ61WYZKzFIgsoxSg1x9Vq0RF1ekAV7HXbhnsyiX9ZPYxLvd6+XMORRnCyK0qdcitt392V2
kQowrmANqKtZoZQq7dtGyV1RlbLiGRubjKnu/KkMuoAlsXSqakClPNYVM1/mWFLYzaM5xaS8Sr/F
9z0F5WG5GPmdd2BVEBbHPxZTv636I/1jeSP3L90f59lGMf3/bWt/2Lh5FLbr6V3wZYb8jGJGjUg4
RXNpdxYWdAhlrFR8zpFRR2IUAC7FR4gbOrHjVdhWLgdSOfMUUjrCBhaBwLZv3no07Qn7JZdfjt+2
LOTk3c5+6KLrSvCXAjCevLwRemz0d45gt2h9L7BAEogm9TujWXICcB2ThDnTLS3aHK2NNmOzQ/Zy
yeJnlXPaNDXyD0q8pdwhfDRagmxtPTDlbStOhJ6aJcoDyZPhT44tl+wVEZVnYAcU4rI22oGzKPPX
J5kSLh/ab3ifFrwTDKM3wVwkcnS8S/5EDOJ7nRbG1DBZo6izTtAn3XZF8cEEIkwOvBoBo4uPgrC+
i7KXW/x531PDSU69ZFBZRqw22vHwjSs6RBzkMY83W6LiXAQSOaAC3sv34DEtwK4XZmbXtpICPo2w
tD3GPd0bKnhvNNv37QTRjJtX5J2ToOOfGXYiKD8GA/HSdIAPdHX48CABfghucfmSyazVlEYekMQO
VkMMDID4r53D1f9cuAW+ik/HCowJaW0UHSI8gqYp50g6s4BhFeMbBP/Xm7utZoVqtBA8NYoheUr8
T136XI99JMa/5rb31kNy3YdKdKB3trj6NwgQl+Gu8uBGYymCSAK77csHkO2tz04gHTCkWqPW6q7M
OAk52ecECQxF3zCmUA43LR9LB2fxnHl6Nw6zjV3qAhddalad9cPTamey++cZgYFbuSYMva33Y/x1
b3Jvec3G7D0dH3jSpWh58D/0q2/PM48wYG3jCsMJ0f4ltPvlswtGjdhKV68x8R+Qs4Uma97/WtgF
4jDAQoonXJvemn9GEm6s7kxYxN0+8BK2YEyHENyTq9IkW52bAHfHgCoM9d8ww9eLOSdMiImQRFsY
V8LA2c6fCq4NBpq5IRx3+mgcY+qzqxnhZDs23g7qkVjAhA1K34QGf5tyoWLjYinO23B0E8AD4Qfs
3mZzjr2EASQD0SYA682gu1n5gs5cEi+yLGVvoZIhf8RJ/aWhJ1ElM5f2K8hoHLatZhWLWiahfOCd
YD5H9nkPbCHgC3ExSfw5lhazBjhls2nY0NacQZacyr8eLwsq+eALyXwhsTiUDufCvmHo3fuKXQP6
yM2rWaA6vAja4Fhng//n3jVqT4Ofm9HBq+YCsj58okjbylnEMbcNDWfHVJ6Kz9kfwPTIF+fRoiGu
K/rEtjGpVvWQWmzfoujxp1NV5HrnpvN8UD0ScF8gNADV9ADIlNrtanr6lxUzpG9SJQGqLTn3ISxf
hahUoMgq8grBpGhPeEYLV+Vg0emfZ0gnmSWh0arRJQsng87zvKuEf3wptQ/AfE6cPX+mh1IdlNow
trl1cIfT7OReWX52oY3D/FMf9To00oBYXby1wImNZgaTnDY9JpxJbMFY35ZFCAADq6k6IAtCrjZK
E9UnDy8GKpQpWSxu0TR/3AKUOGJy+cI8aqmOKUJU5sQWQpMssE7hZktrO55dzRvNe6TU1QQ5b1fn
QYCTEqz8jBR4gilhDRr8M6jlt8ywzO8dJa76VqjG4eqCjmaeiCJYMcVpMQphY+4X7RtN9QM58mW9
FK6tUvTwESNt+Hrzx3SEM5ILIn/EXFBQezqp0g0RBHSL9K84zMg/AetCX4xLK5UqonOvLDVYn1zG
i23WMmlEAULRQt9x+Q6VmlSPEJo6DCjOLW3bUuRXhS4JbEbKRdEIUDF8AjGQrGuEFRJKy/kjylMh
Z3O767dMXZCn7ayE6q4bNkIK1KRU9G9uu9yGSdZv4A1KVmBy3MeW+K+5Cm1HHh74UMT5OTkmIlGq
9dO8hXfgEt9I0m/f6YQZVvlClPUPQlb2BTorpcw0TsQhh9sb+ShaQqjS4ex863Yx4VvvBHz1swxa
qdqMLBFC2CXWXtkul+HVmd13RUCpAynQ43Dio1yV5OEezA+KrTIpOxQ19x2nsAcQyvgznamqrRlD
O6geCTz5RC6BbvD1soXbQ5p2+7HlbTKvMcQVULrwXSPGGHlTBLJkDH4rIbz7rG/Hj25SnLrrpbyy
HYhueTMkusN6GkP0kwuNKSpNuhIvtBDci5fzK7my6b1HyUKqMztx8DVnQYhnrMaK5CJfAiBvCJ6l
vIiSTt/6SlP53KYYLf+Gw0Td5bMDd1BBCppYE9UeBPT62YFct8VpcnXxVqasDwVPvTfRz2nBjZhN
VIzjC5oLyGSXwksty7RtX43Cx4Hj3r5jpzgz67GtpfizO0inNX01tz4t4HsJKAT31j3+4SChuQc9
LBDd/zJoBn+2ji2LcCzjfruhQV7EqcLEA+gVsYtfSqTyO3c000a1PJEFUL4D5p2vQVm6kWZ2ZerS
PTDLni4eqBYM32E/50iPs0fl6yJAC8yKpakHOu+ybzcWVIZIj9CBg8uyv98oOvj51kghCVWOaATh
cB42ZP1yBiRW+iKlpemdWWweuY142/YwE92+RBjKWtfBeyV4PrFwwbJdmkJB4+AsUXixx/Q3FLl+
G+5ViRrasTyVGwa0QbICwmYUyvj8I6MXGb8CoyU7s7/KmnVFGYX5E/oGKa2HTNXsaThOIV4RWh7/
6/c0KRh2yehiOHuMz8Kpq5bQUTrM0HC8H3uziWFZ7uRTfaySaFd5ik2N73zUXaYwxBed6QUsjfvG
6MNkaX+plwVHBZpEjbCbgfQzWUMIB0vSfLgvyr4pqO9i7VCbvibYOxNOUvm1YR8uxK8pNscYWSeG
9KHQp4dtGZR7I0B8MlHFfDjHIU5G+G6HP0GE68bt6h7v/FkUR4rGmYIIZorXnBW2qDuBTi0fFj8I
3jKXo7GvgB3LfDF8JyxlXqwISQfNdGtgHPkjPcnto3eyEU43nSoocHZuM2utBeZ+LNOEAN36TsQv
tXD6bLVNbGhQ02OZp3tlMwXkXmbifiKqYFT9iGJlxyGk/ZbxJJA/sBxqX9RdhujdHQvV9YBRFa3f
eSCzau0GlYyTONhvDT2BjekAo3U3MGxK98K7Ut5Ng0ExIexj2NTaycdBQMHm25hb+AHET0uHAY9m
C8sWXUjh8D08GA+nlwCfIpQlPk47NeIvXzQtLThS9OYVU5lkxci9310oLXQD1O1MEJBw6o5QVjMC
wqsYgpRhsE+CVNE8DL8dc0XpwFAs0ecjOrMx+vVbTVeFfo9DHFxoQ9L1QOBcoI1jDCLkGtgxnxkQ
S7OTyf99P51EXxV7NdoGIj5E9opkDis7Qs7ZAp9+e3CSesQlH3sucz9arfyXEar7azLmoILTdtIr
pGxUo1H2Gcr/4zALK+59ceY/erMJGEQjIlxXnFeW4cwOarhwa4RMGzLBW8drCow3uXW0lkdcsE2a
O9FmQhkYv0Hgu2OIbX6WSEZW5v4eMYVeXj0jqBg0qSdHbSNtlI/FxKwd1ciScXfXMJfxDZE5vFod
gwwA8WVRnAUOihifQYbUpYcEIjYiWhK/QZ2xKyEucbEijtLgXiyYDIP8159RTnjRvm/xjNx2nm14
WfPOMvsyNZr091ZUl1Q7W3daf9IBDXWBZprpQRhkbkOdslx8lvOMb4SKBoCp0toWAD4s88bNxXYb
sJX+tkoIowJDjztlNrdKZ12KkiXTNVe9SYBWBlZjarFziAZE7rEXeCd1356+T1lMW9rbTj6ElOiQ
9rw4FRAZHYUMVQ3shaaX07rdSQ+v6hqB7VgdHLWNuYdlgmGouH6OJUh0+iYPKqhZJxm2bBxL9fTW
2rv+KzxgykpO9nf/fEe8dk65cfU2iBuNREHu/pB9p86SOJDMpJPQ4koBpO0tQXZifTM4oL7s/ei0
BuVI1NHKxVD+C/KXM9QzqV5NqCsPXTl2KxLNI8TdxsFCB1Vs5NGeJNuxmUIvRkwUAzu00lFqJk1v
AsT1LkqSVo5YZdleG94b2ASFUZRmGVFhhS/hLmPNOj10E9P48k5LAZsEZ5Snp7tCcv/KCs8mYANb
nkLUvJk731ig64W2C7g/9D50H2mxz7KRKt9cfXiw/xkui1Ms5X31oQ5v/J2L/yBC1tVA7ptfCwVJ
+gAHtq2u2JEer7lKh+DG4VFW5Phd3NxilDfThP6fUjpli+7SES2IaHc04GpL1/INCInOovK/sZIU
1S+x21azCJ475TEP8v3m0eBWW/qyf5GgAhAXVZzY7+FlWFQXqhQvGf4+rVM862R+1zCRp/S8bW65
K9z/JCLC7B51uHGIZuo6qebM/SCaG8by4HzWHd2F1RWNeGuVyoEYBdeElIMRwNV3TSx8S8DyjU6u
9uPFA1wxYiWO832oCv+LlQby+316grulmNAsKsz+f6o0A1l/MhbWaUWnBgWzit6vwDkljDgv64uw
w0Dv1JRqpuZ3cpEGlwQUdk8UKi+4kTtuPJm0zU1mz12D2nvudi6M1AgLkOEvqKmHToz9/GnO9EtA
8b/tNBohNnO0fRhRWBedC+9LJM4vvYDWtT/6hvQ/+HswYVxouJaJwntW4PbrW1rdPkegPnglK8DU
JGEGbS5TOSbU/4y6fFMgmh9b+tWn+IF1cB5nwyyuwq/hi5BPiMuYlSIhtC2PVsa5Cy+QIX0ZP4w9
9nedvaOl2O6+Sy3Llwx0LuaPQnjn60U1Evcf58OuXBIlk+yyCTIeU+sWYFI/yLCmL9hD7cvOZQQv
+zcYrBlUTSiwHXM8Gn8ZznPCq9Fht2oguUZpuAEzdIVIwsb+lBRpvfBkUVLPB5Xm/nUeIFF+yNni
50a0oXTMvhCQ7yUw65Xa6X+RFTzUYKtSZc/TZafrQv9YUgMdahFKy6JgQjWBXQwIv/aRTL4GG6Bp
5touPEblrenhYvN0LSsVQqHoE5zcfeFLiUoEJrZht/+4cYysAAtXV10e7RZlk03KD1R6sHKDG6Cm
F5mFt+jYSoogULqk6SjEx4JB/9IwZNuOp3fmNMUkAEYlnLgnZXzEB1uaaE2+C7pMxDEOB7DaEvOR
auKwL7y22T1P4ZRmfqwkXA2bdTZdLhVHc3fJvsN5+jJUq4jUuqLq5Ga3/JxkNGeBGHicVp4AD3in
xwtevp4CgPBu3ek/u/Yu+Ld8MkCizBQN3TbRDrUfZtPkjBg6B6gB5m34YSfYuD/v8HDMgGDkCqM4
TeCOh7wnJ0IQBBclicJXEbP6BM+T8bJ6JMvj598OBpmI99sQUvORnuUYFAGjrWsY1a8WsS++SoMc
QGzG2sTS/6NnYZHvdOWcu8660OLz0qat271Fum3dYyy2/62/LqtFgsgBalZswfEIKI0su+BujQRP
M8z9+bZtKjOeTMrIO2wF56XHXG/KvowSPRPnWy2IwfL1BrM+hhOu02Sx/pLJbV3rdrs3SivXmg34
nmJXo3XoH2lHd2sd+8QsM4swoKaKTnyvvi49y5nlc7vJL8hQv4u7onKAhwX16Xehqt9YRM4DA7XS
04ph076OIb/CZIUKsgyVPHt4uJKc7wlnYdV4n9bf9yGm8KGAakc8WxPqmzRxI2xvsSs3A5oNMdp2
A7r2FWB60AY+NQQEJ5eAR6FNNmk04HIHcgwLjpxVo8VFRXOeSGLZfHwHyggPpDiyVUW0IaPLhoEo
qjyZVFBIfnI78oPmMzxm8FMm3ubQe0xQ3a4alB7y+xgjJ5a3xRHfDThBO1WTCKEW5iugnuQRVw6H
JmjQvgG146VyuGpL65NY4m/ugokweuBKRdkaLiGFJx6XdycGhm8WC18lIv+mdI4+RjVcPTqcNfX/
Xer/76lvkkTZVmVQ9+VpNIEScxRtQCvjUMnuerELjxKFF/IgQf48hbkwgPolUcxue99VsoY1bgfP
DKcSTg8N+uZpJIe5kYUYjXcCdifXkiQXVmkl8HhDbw2aghLMYAgNO0w2PcOId2C1E/O7Q9/AG+au
Th3qF7Pt5E36xE+CZ2oDlFHiXTnLLxlY9SyLJAObtLw+sGa3VLUFKTZmhCAKkyxwH8SUCyzk2RUl
7Dt9S2/kqH6LSfuCAiLhYigtQ+RUNFS/EZ+0TZ8HyXAdhkKtE99GwhoVTLqckHIfqltxwsgL2npt
mg4a4KNVog4Z59s0zwRzPSv2IJlXOaW4yYvW1ICa4WFuVo7jP4Z4/4kprGYHnh4hbNF1PMAD7ayz
OGBlYkA1fCumQdUdwLZUq4UOnbHl9SetxqU6sFpiFItoyfzh98nEKq6Wq1L08HU0GN++5jU1YFg+
nTSBxrH7Gtf652ubgMRPzKFBpJsFhqw5B/IKuHPjJzUfaIxmZsOT9UMGg/7IGtHLuQHk3XAPaI5L
3g6udJw7wVSZyHNGK2i1fJw0lKCmpqjK7JxU5sFafDY+7VH8dhqe8XoaoNDvvTlJgFhAkFx5I26g
pobHhfGzmwqF+n0B23QO9ypPcAcxO6V6yBDcf4ww+pcR0nUUP5Bce482f0fUsOnahXSRJIWVQ/+L
e/rqpJ2Nh1fYaKQqO46yIXg1VPnmyIiewmeRwCU1euqInc6LSSm70FLXqR4/XFuRGd9Ok8Z/s8ZH
O26XDs0OGxGz9W9i1Zn7j9R38poA60ze7Ju1pNx61B8AENc42FJRO6P2ebXXhVZRrR2ZJxAyLroZ
eKPGLgPaVGZzvP7VUBgtoIRXXNnxZcjmRH1N7cyEPKXMils46ivrK7xOR0vyeQ9ShZ590M7W720b
AijEgwa8NI9GTbXlP7gHrfbbyUMrdngUAeCGwpJ1k5n+VECkHRkRJ0PmBVBG5EaC97Fyln/ggD3B
RS1zZ03JUO1CogXFPKduQHbsX82HJeV9HionTgTDGhQuj0wOlDzqmE9t39QVSOIuCMOnW/H+B7QI
Bb1DxWKIfHpPC6iwaPsh6tUqm98+UvImCVD+PBbv+E7vNBpxThuDvLaO2R4GJx8s9OVLFduEg5YL
TR0Vi4CyDy5DZo7PYY6vtUTq0LOy9ow+FJoZzBtcZziWtZtSrkLMpmz+KCmtDIhPqa1JY7LGd7rC
WZEkHZG++wlY741YHrLjdmaE49aAn8pDsm/Wo/nW7zglkdiFp4DO4taG3OzrmLlfiO0jpaYrN8PM
BrXe8POS3ihD3y4fQ2p8QfTTNV0XLPxLToCkyKIlv7zd/yEah4mjtcJl6DOfgNEDWTC/N9SzF9uu
aFo5+2WjlVJsNqRPMom4SAe2KZN3O5r3Ao66S1bZCOh/0sbREskyLsvFloYOdFDlozzHOYvH9tJ4
cTmZ7X36Vm3y6fV46okOc4H8pE1rXQUjKl51CveHXtIZ1ssp8IgvpcGl1zvGBAQ/7/36Y6uf18Nv
TB955ZFAbXMMUG6M4PI6sepUo5ovSXO01iiLgJKhPOWaAV6BA0ANn0soqwgO/xPxcXmeHgs/Fk0Y
4c4fur7EWHOkSUiZHK7b0XivXNDYsfTkIUaMTiyLDsXsfjW0UWbEMxuTS/8EBcCLDOKy2LL20rfm
4ZphsCvcaeRyd9VRfFlkxcGklCiF5X0Z7SQEwLoLM7xzKd+sSj4/ldkz/ZhhdJmRXrdrYiC1ZMhY
r8jarnmJu8mUgL8VfdV4dnSPaICgBzEb/3ryjZqxLRRwSR8xuJvjyRNjUxnDysapWJzjqxDneDKH
hpQaDnijQm5f5n21R704IuCIzQ9BOaWcjqHD9xpzgcg4V0sMzNEdrmjNtsogHiyfZr5hsTYwMOa2
tgOeNujna7kx9wUvButHSVcJ7wGhSRTM2iuJigjdz3V6LKkX4gc4OZ7j/1kwSI+Phsp+d6O6nPMu
Fb+4vHtPGngUUEG6/+QHels7wspE33+V0aEHwhklrrzIHQTwWupWg+aaxEqacMZydjWre2uHGeY2
3psBnok8E66E8EFK6F/TeyuueFpT1SZPKsyPSO7jmCAqGiTn2flksGcMZ2dnrBRhcVj9rhNyim6h
eTFfGMjIVtw6LqYmROv32XbCPFZFylrSIhIUI8NzZxjf6CHgSDSKxxnaZNHGJsoI9nt5LWSanz46
/Fhhfqoyuk8V1tM6e94O59mS4vmPhL6kOBVXIJ3D/+M6KvL+pz/OZgm4/Zg967bzt41SbPLJuAGg
palcgAHxFKnAJCPgwCgDIKnTfeLg67iOLnV+E1K42DnJq+YZ7ZJyuE11udhyPyV5XTL/DOf/Alja
6g/WKKu+qev7YeBw2mtN0hgNFkpbzFHh6Q3qTKuNhbwXSdNO9Q2MycgVHcdsE63rON9pnrgA7XBx
RZ9/4S+9TKksBobCx9hUefoo4z7IVWAevT33v12f7FcpSWTPLv7a4Hnv1YpEhnlEUk7qLx+MHbI6
/VkzHbuJ4AFJODOOqZpfaZP/gVxgSltOCN5jeBU5zq+91H65kdkh7JZOzP4DZUf4UtSdgOq2cEkf
ct9uEm4nTB/1K4XEW1llVVvr/wgKdxBVMA0qA+dwOstcDueUGnqjV/X/eLswHcRxYw27FSUbRh/5
dlz4hXyU2szP/ghndmYRenbQuTEXWsGiaFXwNHm4oS8umMJwa6+/NloeO+xm0bgEMGdYy7fap6wM
EERU9d5FOZN3Z0Ol+89EFIpV3aSaatPZ5tSvZmA7NU9iBIrPTPN3r6GM1+VarVamI/NXJhp5rEF2
EGoj+MWviuhyUzCY3Wtgrrc64CYGOPDIl48IkxNKTW0Vbb+Oo2oR+I3M0Oji+LB4gcUIoaSuDksb
wEgxm9GTZ3kRyCoE/Ab/hHduSQeGcBTGIByJdKw/mAiExhbxtLpWDtgIIEb9J8/8RilRpmk+0uL8
1oazIXBju6h3215UQwJxmDK1Xnb/Zu3wudRXgppnohbci6affRENmZeWNIV52/+FM5GY7gvNIvtB
9Oa/Stk8lJAAmWxmUUZK8Ine7NN1ZIakXfJhCk5C/PAiavmrvEWxMwTlZPvOSQNdL8Jd2LkKo/qj
KBC6COMwWC/+cR1i22ecrqqOpJfD7SUh86QPIQDew54bLzjjzqvA7OQ86AszUn16a2UvF0oSm/gy
LXwfPshHxlQYmcatjX79AiT2ZFUalzoAi17fQ5rk2yjPewbikYVkqtS5c2OCrLsKJJCKWB+jc4VX
jebGK9TjjXTc7H8ThgdCae2AgL01U7dwQ8SR35N3aU4sSBIR0BPFZPZq7zAsgIacIXwLzGu2a4WG
a7sM/5irjYWo6iimKHx63qb84BAslHRYqwBUcNaV91YqcAnNnVxHgle6D6Ux1/lrjSUSTZHQzeW3
tik+vLXMRAeFpMA5QlTucV06jSadOAIZ9O99/PAUsRu+IVfc2jHU8M/eqvwl7DvMW6xW79/I8dUS
Bkau3D/WvXuM2nDercDp0O6bAqAvx0CUfwXVz1/aLOn5sG746ggTJW6wG922fly8EE8ZQuFL0url
m57GTqBJUPwSde7phnhbBPKxuFF0wkw5egj3+7+PruP71U1+xZxXXAxltOgII8FNYA6jd737SG1Q
+irxq1rgk7YVMfUzBk9Xvg+mvEOyGLXiQ0ttOUREeFwPG7ewKwM/6uvmHG4zpiTJgoln16atap7Q
DzGMthXMeSrU0jTxV/wE2l4+Ciu6nQhBKTYZ7pKG1s6ZFShPEC/zr/iXDuTDwUVTlufaGxQ9OEY6
ChGkTVqqqkQJAuH9w4EEBX4tq4ZZ1mZpnTU59PAdeCXZlYUJGze6759LXNz2paoNetZubWItSvrq
hP5MrfcFC/n3hBO8WFuUZrwCrVo3N7v0iS4/tj6+m75Nt0ToVUoupXaVacirOvxeYAsTKRM+y63N
SUwcn/ij3yJySL8yfBYuc++813b7a8adpPtfaUod29nALlSeOPmtRH4RzWxNMHN9vM08ff4OA4Nw
khO8GubEiUkBala5PWqp+9dkw8iLK+qTF5Of+G+/zwkolbRslHCYBqsmEcQ3pA1AWmH9c0P5Z2ID
BWA4sD53pBplif6/3PaPXvOFEWrTYOmR4e/VrazC/7FYmUnWXVVTkcA+Uyt8Dfv2ATGp6l0gFI05
eV9HAFZFIhuvxDweTX1MAoTQLl1B7vkBP4uu/r4MwtCuzLvNhTxBG3kDvyyb6xZGTxmuRVW1pUjz
B+l3+1KKv5Juv8pNxV6IrfbfCUtwE5wtKsz+0p3F75M64XsHb65wdutv1c7YqiNOxsAAwp5XvUfo
Bwi+bPJk7O97fclDSszCrplZr/YoGwbAht09ODgcPPp3Q8TK5fsjwem18aKxUap2Jt4rV3xt60gb
qyNztnnMpXWfY2TZeVqQhbfCZNiBFKEKTXWEGCSThLhrLo/ylB7PLs+S7fjMOFRyJ8tlrFimtgo1
GcZrJrXBr/Xa+g7NdIBfrq7HrbD4Wyoi3+4sZtt70ls5fT2tgXRdfYlE+NDJ5DBmGhoHUtOlsC/p
DK5r8qCv+j2jI0/ej2WRd2BaZvDvR3tGu5piI+neMFdtzWXbD3YVaoCYWAKIY6TkOtOgoanYkqFQ
Ip77XzFaG7k7fZpeEh1dtrScr/RvIZdvPAqtcVD0GEh8QntUpk9wHdKq+fHeyZGZl0c11/j9n4Nf
YHfeUiLSs+fY+I/Y9fgy88rmzFslB7HDSunhCIipau09ZKt1zGcdW19oScXaPOJY+VAHKxuxw8JS
3xq6jtBSVCx+sdlGxpMWsPifsgE8AX+LPS+pHF6EVf8s+joGE6SqSNIwjeJCFtJEbPqHU4mUpnzm
t8QMZ+xOaz2eEXaVDaeZbBFq47tpBgrZh+QQ9oaKen0BFjMY4nA+QpdjuTqwnqKRli9YQ5aup712
ThfJoLep7C0wMrLuqkBgbNB9IArA9F9IxmvEE/d7AQ9mrGay3GTOBtgm5Ufcbi37VCWfKwqWcFYi
XI7qnyBDov6WQ3rTuCsJ9KquM+jF057/gLoKJrm+ZkfGcutNH3uwxl2acKH4YCYzn9NbwH7FIqgy
36HajaG9wRZUA5homcOPMRk/DCkYN6i8ZmuI2VL/Aoy5lRjFF72Rw0t2heDi7qPjatFyGAeActYY
X4vavduelK2RZl/ReIpB75npm7UgW5N/93+tCm1Af86lWvAfTVOMZcnqjYYgglKPwilLYhdLmXTc
lJiFOP5o/oN3nd67rHopYlzAxVPDxnWOC1wEZXP/SEgx5vGpgdJ88tGlYtJXY3NGJjpnnCW4RgVr
Xnxhc78J6/vyWRojhwS3LxArcCXgiig42cyKOwL4UD8+IUGx3freS9w2VXVMjcal+C5MMOFEwqr2
9Rv5e5rLVgz/0b573VYLcWhdWlK0PNCcwxta+oXG+rPkYYigSRA0i4bbLT8mxa2uxoK/9oqnZpfP
l/Uet3f4mWuLW6HJ864I/EmJNl/OzssHM7BO9+ZqBBn9UhapSIprXhqVqL8TlokHzNje2ENVwYA2
89LGrQYXIT4kICP2Oe4GBKcwRjawhmtXTdlpjbrAIRyb62mWm8QLCwHgCaAPx/hB6Mcgr5bImEJL
tLmZyDZQ5rQNGV4hJbJeGR/9UzbxUy4sHLSeqCGs/BrosY4xi0rj+ML3YOz3VK9SlEWHdlb/awct
+Y8nxHRrPWQjRCxj2blrw5+GbG+svwIzhwUhPgDbR9uPL+m73IrKZEUdT/Cr0RZ77iGLErEwNqHJ
ZPVfFJ/+VAgbla8iPoxPjDmgsJglFL/gJiCNLLK3AAS7UPnKhrYlnqTO/EtLJam0DxK9oz9g5bcr
ijbvrFVaZwse0Cdd9v2aux1CScBLPFSN9pWIRRoWQx3++zUCI2paCFe+6jC2197PPkBiCRta67Ea
iQsoPWAHGkfOByFpLTcKLMTbMt5897pRsCg4fZ5/W985nQ1comtFMWLDApMVb8Q1MXz7LapA20vA
G+DQnWClaTrneseNQjN3pd2ukmtOl5wZnjN/RJk6rHvrA8fSkIQ9aGIFdLay3dRkAvA80wH8mzUM
fCeifTy5nsv+PGekXRfByTXu8g/7iyxe4EoNwNkru+ZuuRlV1yq+Y1V5AQwnZFla6a1vePpmEpaZ
JplxQv337L3nZ6BZy/jRVah7uL3XrUbA7eWksatm3tGxxdN+UarlwSAzWIMueXbPyAPiGwdQx96G
E5QCW/OACPhc6DiGAjEEZddguSJQjN5gW3rK/+p6WfApVyaai17eIIMBgzEWvgZmLRVV2awRYRbO
MntxggpbhRvEShJYM2MFYMVWv0kjKyLJpdenD95R62RG1LGG9OduCBOf8qOcR5MyppvlHYBEF8iu
9mDVz98pfrtkapMNIZuXQ6K1uOfT6yiY6hZt31V6Q61PLu+x+aj66cD6ZYfcg9JtZUM71VS6VLi3
L0hq69lgJDHrNk5Z7ZbD8Bo8b9mmuh1982AZI3Ig/VOTXyEImPAu9KtJElPntNYRGakjIA3qv/L5
q3oyod1lXwQPGneKuvQRCNZ4SEvbGFcOfg0ejRK/VV86UjJ3m7+4h+PzWo99FYW/NoD0CRamPfQE
UpS3hV2XvO1u5FVIkHsWp8wTxoc85ORNisDyNEa2k3tCITJU340B6RnB6fVc6sA4dw0cPRpPT5x6
b5u82zPkK34if/xCG5pE2SnKZqMjVBfA0214pGb2nCGn3z/6YT6od2i7Kqu+p4lntIhjceu4sTst
2I0Q/4pS3dvSL7zssMknM6NHzMPXrzHXU9cRWEaRMgj6j+viQFay64l3sob7jmU+5Aj7J2Y4hzPn
P2VL2yLYFMZ9eVUrcNys7Nx6CKD88NLKSqmAzwPFtBSI0gOUID4XYF/wECjcFBj03w8ubprsUYCn
MvV9CaC8v+scYz10xESWswF6gWIBV4uXCTq7Kxh+sfIiF7EyMr7aOoxwyl+9seD4Se6CESijt3kN
r7u5hkVN3ki+IYTMFP+cUhI89+k+dQzn/eFCfCa6TLnv4XXqd+1IEMO1IZaNsCnFQYQH31/VxbmF
e8XA81glUbetaUBJrrKLI2Oj24hmtjOId3vJhDv+CDiseBXRTajUn+MaWvu9RbkqrqTuylGtpjdI
jmdIM/6+M/GFXpC+54qkggk9FZeqgHktIsy1VyXOF2oQBHo6JHwlPYphmgSInIhr2XytxBxBiuKw
aTAZJ8+easORewUwRaFVyqWhOD4S37ZtPlMsblb9PlnN5IflgKIvtT22NGlLzCH22LyH/Tlmm1em
mZVIY1PbTE/RlixEevZUVcBxUHKVcQrLm47KEAeDjK8zrZKAy9FrEX7iW2faDTA8bf4ljEXbrYk+
8v+3LHkLKgRjpCGyyREOJjvL9jKZ1odILd2MuO565cq4MH0g0jrIfscGnpClELxMfJGgdNempYOq
CSVX1Qigqg2OCMmMPrKWlv7WRU04uteHbO754a8SVIgzciOQgITHun8xOuTgMUCeXg7bJi4gPJ/6
X/mM1m4YkaW7s6Xrn0nAz6QrfoL2fa+NA9QORA0T8c3t/4GrUi1/1x76DfTxEv446ENxdf6xvSVP
OsNr2oXhAOI1GbaH29KGtOt7OKsfFBO1mXkEj6IA2n7uZZpPlybIcKBCKrvTPV5/Q4TbvQh5Wemg
6sbqW6Gb/Zgde1MNSJKs69GENaFGk7JLX2YO1oO0a7a8i/sMjpdD4uinU2WfhL2pc/jxLYXgUMWD
V2aeJo41cRVFJU7tfQp45ymDAQ7AhEf8GafZyrsGvw+5z52Q7nzo8rHJIV17qvPvwVEr2IVWk4J8
swSaZSunr6oXnqbJhPGn4scV+axJ8OcqzVT3FzZiu1ITQ9N1fbWpe/IJowmKRREHSZwphnptIbi5
EmixoC6kiMWjoRrc8D7jfAUBUabMt85obYbPEE1Y96Q9tm6bT7yb+RUYUYFqCikT0ZggVQBQDo+6
+2fK+SKaNi4HusOqlj7Tbx9sNCTZlWTLAErlt6/bNWjLdtZKLBwsR9abfQY9o1XYijzUqnm2pzfW
u9YsOfQpMEbErU+g0P6rY/3lGRJr2g8kcISSt7wpY3h4szLeCoXWJrg4W3HfkBCA+8Xei9Er6PJO
l4eHeOXbKjZ7aV4iNhvJ6rCA8U8IrSPPpwhLDGqX1XZvNPePJxTWiqnyNJjPKmhaOXfivciaKFcz
9j+vXWucgrliAfXqCWiuLz2oT421ugaiuZgF5NaAimGUhRvWw97qRh0y6wRxFPXgdCXL0zooH7Wq
J2DmgZC5DLXIZzq3iC88KikEhtPcILt6JIA1DKV69I21oYeqBl7wzo0R/Rpl0fLOHjlEi/nnQrqE
MxqTOh4vNjFX5pRrqIZWQcCUJr/8aWIUmrnL7oPD7q16Ue3s9RgzC1gzU5qXyPZDRJBJOGkGrjhW
tcE4jvMsQVuoevsQwREZY0DLM9VSQg3ui1v7ZpM1x/lBQ4yvnACTrGHt6gmzD6YX5l2spXawDZBo
eRRWwxWBghuugBAATuM5Iv+8Evdbv8gZ517OD8zjQi/9pGg1yYUGeNGakzq3ss2TbFkAVAlN4MJI
JBhdl4Ny8bkZPV4cbrgfVENdmIKpmk/6XBHa4dv/aNXaPS1TuXjF1mMzA7gZEvEZnBwJEYv4oGQy
6/mYGZ/qnAr3OoE6N0TMxg5wj99T1lgJwCmqMMrwQ9uguD3NWqfhbk+Gt+FjfX019BAWWcaGQgql
kvqn3R+7PInhUq4lZ+ejuZBNLDFbsbe4+WasALBFvz4bx5hm/GWbdsZv1rUAAfulmtRn1WxY07Fd
hMWLpSZ7zNj+NShwASTT5hroAqJ6ksHTbpeVjtrsOwhzgG5+af7fIukPtvsxkNEKhVQUy7acmyrw
BdnfbtgE/6ASQHbENKHp9UFhWRGEHq3px/83kGp06ODEZ+syi79FrijpWshRt4yxJE8bBDK/m1LK
gI6q1ICYoVPhTOt4vm8oW8tt4deGtX65KLc2zt4efAML2Rj2IL+vyhTISOeVMJgrYuID+XhCj0f3
etqeUQGSdPUxp/5A2xXJ+VpJcdwUJGPFjhwO5NNmXJkM24kMQuUkCD40B3rO19o+Bt8PNgGvmhnZ
gBn3W5Phi2ruKL+8nC8sybFFtdbVMhS8qju6qMK+ncUZ/tnh23Q3ZYGGWpLvrW6CRQHeWkzVRZJE
vI1pqnKBTmzNXW1NVYr4mea/L4elJQOeeHeoOdJSpAYdpOgo1AvTgmpeZwe9+/js40ofubAOiRRf
kSm0tYWq1pU3JDzXS2wkDSY6Czj+4ocuchf4crN48NTfyM23IdWBEHLVxF0E5n5PhhRQsOUZRDCy
OjxOiwT0vYfEq1y6FB5EGihXz4NMkvoK3Yf0rbzfIvP2LR+AQzgGkh/u4tlcqlBE5Z2ciT0/QVTW
VugzVodCS2PIHQbs2lxEjHKARgNM8KTuiZl5W637wga/JNgKM83tyvcAhcp8sdem8C3CeR4UzCDQ
030RGqcqfb4WisoUczyOBneDQdq6gZrwFjnwnJQChoy63vDosYVxRuOZ08+xAaRHeGaeBGYq76e3
TqhnP8K8DHZwiipUZIWIxhCKkFrSdhcPuwAp/7ZFPDRBh4UzEyJ9v8qF1k4S3TYnWprcE553DMHW
SWS4xKHlexh0CW0NJDdRWs48cFIZbqXjWQ4JAZclYEbSDsQ/0TgZX5BHqZNSmedi5+HGx6R2WK0L
rkLd70ELPT95iCDqzVhXRLDBfry+P1MrkNGlOMJy0hdagEc8AeSvcb7MsN/P33G56uthY3BDv4FX
LFm9JQGPtDn7kPFGixq8C7QcEamZFpvCVpvtk8Q4x66/UIbluxRKohmtYMroJjoppaqepbYrQJF0
0ig4FgyC4vAng5h3aW+Lyl8ihQUXxcK7yAoKbR1+JNG7s0gjcExAqu/hOORfVCWuAYKXuMZB1x1H
XHfqRLuFkVcN0CGsVPyyqvz924+rJRL6d3/D0WRO2aIvR0x588ckkKLImILF0fx4GBVm5XIiV2+K
MHiVDXnrrw2ayQ/Uk5JtbfssvsFV7B8i/WXiZcVeScVT5PwXL0UpRK/LExxI0ZeCtlKpgT1Dze37
cHcFRw2CP4pxGMx7mEF3vAPUpYPVu35I2nRDwFwUs7jg1VlDieUAQs0YwBjD2CsIAMyFC4xaiOLQ
BqrQFbWe6zJTwL+27Z+kPMt2sIhLZqZLuy7a3pNzBMrFr+h0Lfe7ZhMlSqFC78dyop8RWd7RCo5f
bvduCb+uiYYb5FdX1UWYu4psYtp7qsByjK2arQbmtmTIpx5sXc1gMwHyOqxKYi8JLzoBFfoyWwNl
rtcrzIRVSR4ym3Ow2kXyWM6f7R2VCD+aStZjXT3pWDN0VpSzjEOzswG0xuGHT7tSI4Mk83Bhaqsj
h55pWbOoOT85QoZilC727thody3nlZlhAFThZ1a1zhCYNW8H7eMZSupCaptC53+r7Xj+xi3F2Rnx
RC4aT6D0IjAa7RtW0g+bg6n8beFNAJjJxkFOXIvtcvso5YeZ8HbTDwK0mWy6UK5CEocHb2bkm+et
XoZtYlJucPZEKD5rh5bJWrcL0DInbdWwW+W8Xx5cBv3+mQkqvI+JIrR3eExJIWGIwYzkqC5xJjG9
nYoULuT/W8p/5OBQHsBQpfxJB3KXsGwGCkWuIKR86GOhwD2+j3OftKWF5NJidc2fxRdhEU+6X0Sy
qAhMQMtiBiQoyMRFF9Z3ELK7yB6xCYOB95BUKoZI/kdi+FCzL6Xrq4HSdgc9WKHr1Eg1NIsFRJFi
aK6my1E50HmfzehbpdQQHz9wy6zW44Wq/FdLlYtwF2Rjt8MlT+bT6xUaBOhyIyScEs6AY4QjUQbv
pVtdXMplvrf6Ijk0gGy4pAfjQe1eDYq/sVyN9S4KErTOHYWZZrxmXQObUyXLF2sbONnPmIcWaaCV
V72I7FtvvRMCyvDiJljlbM4Kis1Ma1YQ7D8Q0zn0pL69MpUYCYEpC/LVOvNrXaHy7A7syJKZ8LLz
bUIYnFBLeIFfKm88onfEWzKomVTSY24aBA00kdXK204b2wQ1jrXcn1dQxe8CPcbEDohSf2yGAae0
4V0AjmiWutvzFFtqpzeACyeemEFYW/VZOZ28y9d7yx7ltNGm3s6Onin+g4x/4e6lt/jzfYZvSFdh
rdVoP2BNeKTHJZ4TxgLhUUr3GkBBCRwnMveGovTW9NHw0lGQA4mTv671xrRHkrdZ9kbXbS1bX4vS
b7Xgg+mP4sDHFtpjOxnyP8ib5oJrA4hDorcSUnDIDAxHvxx+4Axo0GoMQQSQWE3gH5K2MGKc7eG+
X2wJONypqz6nN88NXu/Mb9/kmxCU3FwzPCHjZ+cWyTrY5NCnyN7RpgkDVFLsE5hPTt/BjarLNIVo
8ET2DsUaz6BpGnd2OafS/S650xAgTkPyyanPb0OJW1KzD6tPU59BEiCoNpnnnF49YmBsSN4RIHhJ
g9XfMjmaYaJCsWs/uBW8VlsuZkqCXjnWkLDY2QABdxnksIjAhpzWWnqk7r3y+w1RaOkoL5QfcnVi
ntpLkwVDU6ZvtvIMXQd9KdOCUyVosohoOEuoFRStzm2rGA+or5QIjeY5d/a9eC5QYos3NK8k6GhH
I5ADjyV83ZCTP1WtTmPc8Vug0Dnijstj+cUQq8mZGSH9QzhpOX74qgawoIjfVDFKfcDPWC5hCqBo
SVKLtv8+Pb0ycXIN/0gSREkxjh1hXMI5U+386pQ31P8a/YsQ1VCi2/l0tzoTOTnlzp+A2sTdJnwX
SIXJP1L+Mbnh0lDmtUd7Q5L7nw7qIb+qAj/6UTFOD6lEBOHGUxmiJm4npf0JymWsROuLtiXi1sFz
QU6KPZ+a1kI58/grfTidbiQmPtV//7sYujiFegagJpgGIODZSM8zc8oOSNLWnhORouDwcMse8oy1
wQWmmVH2aGU4VupiBgHU42olmJryAml1IDGj3zXbS2EaZFI2bn3m85ET0KVo2hbR4lkAgf0ZSRBW
6ppWkNMJOQDdIJyRkNklHkjJOZ2mobtJHgbLobBDeVqVQNQoo5VZmpgkzTi1F9e7dL63bdlHkFs6
THTYdmC7cSisyXtn6Qz6RzOTM08neMvXoYYD7YyndyFXyJALu694aOlG9xXs3MHwjtfl2Fxarvta
a9gJo4qVJzvNx2hHf/UvvQt9GVimV/uZsYs0U+6DSZjsEFM2JjaczpSdDeJej6A0pdOpKea9ik21
/xmyYjkWKtX0BzvgWc6YtTtuczGAxyGjGd1Umen2SQCQ+RRPbTQUbiFiNeFtoulkenLnGy5Vczig
q9ELdcEGHE5A8A88nqBFh36lDNfb96vKfdR0rKN3bOm54LW0VhJ9rcHeUAZL+5b0MsGt+QdGPtMg
QL0iRiZPEuJSM0U3QF8PIn5173dHqd5bsTAbhSj4b0FigKaeo5RpwxefQdXyksratRy/zh5lZ46e
tef/mxiAVHl06GZaQnyZp2ZC/R/6SgJL+uPx4W/eqkVXNI35hvp0zMWpAjFyZdM0skbjsuBG8OCe
Da9X5sxTWni7L8lVjNEtKU1zrs/npkW4owuVo+FhzusjvJL0wF+lb22agkK6nkdc1bsIco3GVXMx
tz32sLBSeWQkwNUXN+wmSMSdQbZ+TowWzZmT4wZm2BjBDQ0/8PkDz6pqll0xaKzI9c34WePccJpF
/fADNISnolDODUYVlspaip9gcCdiBF7B9EKXgDN948fMGb3m//DYSRdbr6ptyZq0ZX4fYJN9m17b
K7UPwMjTsJ8jpcLDkPYrgofjdVujBTzNSi/q1byNviNvTeISKxwJhBtYiimeVy9M0B8A6sBGKbz+
R16ksD7eRxsy0A8HK4ManYWTXN25jkLJmDFNlQHhVpkJRorFgEXym4oFjqRQs7di0nkVdaQdiL7Z
Ir1k7RL0fy9QurVR7KXgbgFYw5xFFQtLJfPDL1aQiHkijEGMEX4FaE8Gg5o55qpP3kNZU7LPu+oC
f71nji9Wrzt303qyTUrupMqkzBt1FeD5xdP8TphSpcnCFShQiGkMgZcO8LNHuwbPysyaDyRRBibo
4xvPFl1P/bn8c03cUHvBWbR7Dt74ec5WpE7xMhh9DBGeXsLknmvRwEbSNhKd9c/mfoKilWXuZTDR
Tfdh9Oi8vPhSWa/iefCA36VA86w5cgFytg7VxNTBGf9lvH/aYGrM2aTtxmyOunlJCSPR7x+0LKAt
loICw6sXIHde+FTNA1wHKySNueoMX3L1RJCas1ZQFvnnIF6jAinIB0naXn75gHQTvZv6o5Cl3HZV
Mqz1+XAnCgdTMXDgkIPNPzHJ5LWBbC4JUxHmBJg1ob4Ix885SPGoRpda9RHukV/IexBgNS0KBSz2
+LyvlZKSLYZeJjcU3dDJsckQmdCmEmRx1Xdrv7IYym99M1dtL8PEoFFDgzUUYlUWUIm/oY1xHuTw
+N+aIdwDYYzkgorfsi+bKC0r7q2n2l83xi2zC+ZahTvp1SAQPtGS0ZPwymO427Oy3tvs7A4BZDbo
yk1DoqqjZeUyLjeXyEPB8XVACRVgGOGQWVrWTjNNvWZQn7xWF6IdMqpVPlORMZSlL1U82afA+9Nl
zKoHjjr6v5a9wBxbYIngqgiBOoFrkPXdBb0T3cfDlph81fQd2WX9yt7V0wO1OcU1uUkUnUFIhy7o
BDCvvvCHLl7s+nWZgR8go1dMThEbEsckzMozrnRarFJeBHiNIkAK4oGMI64TRDVTIRbEEc1jmLdO
hzZituXmQWi9OZZRvc0nkFtpAK/285Q0U2+UdJUrvlM/6za/56pEpDMts7vhxut2KHOPcLidHay4
xcEz5MakMlDAL1N7GpkpGuzY0+UaA0JsnSThQkczBJqS1/NZDl/e4RPG/gkyxLw6Og30wjxaTpo7
Wnt4bHctXjRZeIMIN/Aii5PpiJkPoLftPGvO4UUhhfILVV79tlexKOM8ajcg8Ny5Z48/Ib4AxP7c
bg3qVe8CWyu/y8mYpbtTdZXhHYdztAf+4ASN/OYAmJq1U6ACm8z70dUOXVOrrMCON3xcz0IqwXj0
UyfMB/Jx+QY4Bt0TdG2aSvYNWSOgW690SLjl/kpLv9+7vhX2u3FzBCt63KqyNhH28FXiyLl3VcQL
OY9QsHHzVtMBV8xkk1+dMFYH4NSok7Wnds2eEfnObvFfeUx6bq0ZYAPpgfodxiMb5bYCXF/yq1fp
HG0Uio/2RsVDMIIbFrnZsYSmMdT/xlroWQZjeOKjbKD6jVLus/HVgWpbbNCiBFxPW9hlGU3h/46Z
MXc4DxEXmdWppZ8BYiJOtyjhD8eVSMfuZmG2YS0zGxbgtrMN2u1P/NvxXdXpuAInmt8mpP7L7EDk
0pEWZ9iKHVcNAwB6SyIQt36+SjLato+sTuTJ7uc4WWu8TtIMBl+2t8dN+wj2ql7s5le/MnXPU8qp
+BBJVko7sHPs9UYMZIG1oAZ9Ps07ZSzMdZvl5ZM/n0yAxpc0LQ3M9hwsRDAXoF+suLD8j658TlNf
tAkYO1Cl1QtjrJMGs4hnlvcCpX+hGtoAWuttaiPBjzHyChSwdlJHP4UENUg45GCZEVP7t7E/w9XI
dQ+O5SZM3UXVI5cJyWudcIqua1TdKOBw7dJue2kL2/VSgfmcqIOl2uGTbQuBtH1rZ4k/16D0lCJ8
+/MK3dD+vDS812V45wPXenEAS/InUU8uuvMxa5l5kFrqc5VVz4Tj9pTRUKcbCOdoi9Vv50AXy/7a
E+FhqZX/cyT5ncYPka14p+ZE2XKzNQZFYgVQkmRyQCSicetpW4+43RoZwHiGd3XA12rsty7aolOh
EsiIQLgClUByTPyGiAQkEr+g6SymFNlh8mRMHZMX0RHsXjcL/5cn44+ju579BcX1dEnceYZZBW2F
Rv2C9pRxXvZlpzo57wlK86//QkM0wMPlfFPQHhmcLpFvxOIbcPfVPI2XZtjxAlJpnndJeO5XeQqU
sWEQy1YmRK3ulO4jKxYcm5PLuAnz7HXw7SuRePM2hR8Nf5JeaEqQ7qg5vrNLUyVYPtbVHJ2lmLEN
hDuXf4oQ5WAKPNH1/9RTxu5pC1R1GwEZlSoSssdJzSYdIfUHTMnga1LvIwt3KXaiwYkZWCpo0143
M42k8LzIyb74SzPVTZy+VTlfE8eQkHYR7GzjtqWui4tvREdvInhHEIduBSmaQhz5RDyvD2Uql5zZ
krcaGKq+2mml+mOBF2BgYP+WTj3wCeV6zGMq22qSGyUMU2YNKeBuzpfIFJixZzp6ultL78mCQ0cp
krlL57pSA4M0eZgporbgQ6Q23w2cY9XxVwdf697L5JkPc/7aQBdweuWB1DMK4cgo3MKwYkQeVFG7
QUN8qBsBBHzWOtcU5BKlhdYPFtXw29OllYshQCS+MLKrp9x5w58mHJ+s9Q7VfS6dgvABtCuE4imN
mCorm2hai+No/H0x0nr7uFLhymKLblCZU5ZoffF6PuRX/lUYEBIk3tQ3tlmvBmrsKP5ZkTG6NmHz
EVsiCYeZQlsdizss9nMGMkD1MHEbPo5btR2eh9L2PpWdKi8d/YSTpJf1FfpOBsfCkzVsM7F8l6NZ
dlmZ/sTLunKS9R3yaJotiIPA9F8Uv3lxZ/QwEydcCowTysOOOOUxxKAVn96h/9xOAIzlDs63d1Jg
dyd9jDEPCBiK6Ln9FNG1o/IwvWJLZEHh3YPYqs0I21rD1uEt5XMaq3D/Wdlmf+Dmu1VD2dBEHqC6
kwb9qeZ7EAkumzQq2GtgF/uvsUOpsfGW1j0r5NH1rI8tadYccFj4WsRxfCdKiIAFFUM0J/O4pZaz
2hUDU5zGJO3ECYV8qu8P3wdLBlLghPxou9R2dkv1I9viWdcnNMkuR2kDDW7EfuaWU5lM3ht1xzX6
8ci+lr3oaFgOO8bpuurN9/R0J+z6TBnVapecz70/VBnjPgAhvvV312ofQ9ysr9Y9ww+Oq6HJCsGj
o63xvLVCir2cSAsQICQB68d3oMrRIHipv1SAMItkvHRadp2Ua/a1kk/uHwe12CKXgxygPaGZVtJ6
G6HE6aib8x+F0qnE9mcwR1J1PL6JkEnUJbcJdSTfVc8QWktaUEWxE2ZOkfGZtUnM2BmsXfnTZawv
2N8wioxWLSlj1pLoedJuAd68uITrVvbC4P1xNC7VdbJkC4h5XDBGzvtuS1tfn6m6n6Y5qEhoB+8Y
ysLdlaCCyXD/lJdmCUX3e1Zs9mWeCEGZSlU0icPM0c7bPi699SOj/fCznoXSauF6hL0EeRcuqLBW
mlbkTd2SsokLLYrtv+w7yk9C6p3+JqpUF35da8Y/0E3S7ddXZHNzx/HCKHO2OG3KjZ8K0tNiD2PF
0Wy+yT01ejz14ekXgSlbXmEAurO1+d05ayBVEZKn+zRpouSoxg5pJtFbXWHJeh4e90WVj+gOV53c
T//TQYFjnSpkmT6KfPuBzPqgD9HcgGZHAGtTA/5X3+1c5X+97Xq7xqFN58iex8/+ufFA10Bqp4Ce
KouL8Mj2RiRKcn3z1ZBnZeBQ/Czf2IhcNuEzEqNCccMfcxvjHAmVaEEyCSHi+e+LcmiEcJcOzBjL
oFUk1FrOamkd6FWtLjKxzDH8HDbAhV+Gm3txI7kRqhHyv7WjlyZ9Aq6sEIVHVGY7OAL8/ZdS0WoL
7Qhfc8kR53VtX66QDY+5dnlYhjT7Iw5rfdqNdiFA33aAd+cWJZcQJFgRth+J+IGtF56Md7tNHeRW
ZtLsUtn/rbs8RtIf4/+vUNz06SKoHNaFbPsZalxGjFmKCvvpGzN5RMWjjf75Pu900Jx7BfnSXGgs
rWitRq7b71nQclvwZaO5UHCvjRvCdbN5Oe3wea/pv1R3CbJqyLXG/fu1+dxTS5PR3APJ3r7YWosK
ZxINgqzjNs6tAYuCbdsFo8ZQ3T+bI2hn+x7429uAJHlKf7n2OVxx1ITw/RzCx1PqT+SZ654BERBS
mkrLopBQA7k5crP2h+f5gpgMSa3HTRzJcBb9SlO6xUnmpDXcLBjGJIFnTSDaijIJRnY4QuETq/pk
K+puLLBqlou6EVOzTdLPiXCu9fno+9rDfzDqgnVY3SOtIQfP/m6yb8Og9pRuHRuWdx5GdDdYueuu
rUBxubCYxSdWJtpUvkHabfwi1SwsS1XJM5m7d4toD2rDBq1AO1Y475ZXEbwVk+hA6uHmC1JscGt9
tAw6vyCAYJpEZgLUawKrJ4sIayWkPLQpsefcFTprS9vzWG3XMVqOCBHqNFWJYopoZ/GjGx4D3XaK
0T/y6OWgEVn5JR+Cx8H3do/BlP36+iK8B4ElOb+ztE/YU3ds3xHgPyke1v3e2ZE0798kujYNYxpd
NH9b+VHpbZYIgUh1U8PT3jjUdY+AMS2SpXaaQSAbzB+ituw/ed07NBDCTXy9iADQj6C0G0FhnCSu
Rz0inwNvokj+7ecoWd+ZnVvVlPp0jygbK2xrrxqtC0epApDHkXIG1LHZxIxO9+3wuh7K5QnEXzbl
OHxO3C02M5xHGRURrc5Q853z/otp6NcSmK1bc1DYqrg6KBCjdgMgGRy7drffpiqDm4kcez52vPTr
+554xa8BDkYLXR07MqUN5tv6jCfdo5z94Dy4I87ygIsrliWKPdhF3ra0cxuNGfO/z/FVTXv0oOXi
I/mO/0ouPpwydpRJpopZbzWfjBXD8+PsS4iBnX6HiX2wU+qeHavLywWLaoXXUetZT58GFYFoGrQD
kc2EOF1e84QcUzth7rVeZ/fUdZj4ztqUEgCjdRFiCbM0+8aLMu07RqXaF9+XMt9Dq4dUdg+/924J
W6Yss44Qlk0xwZPSBOLoA3akD5TyyUqS/OzyJRLbn/SWkFiq/PyJQacTrC6Db90LPZKWNkNmMWDI
tghwOykjtug5WuqcIQpikZob7BLLOlTUPOSEpouBqBL/AMvWIqrqQ3LqMFncyAaciqf2qqkEoiJX
TvtxHhggj8escn2paIizLt1JO3am5q9Ia+GK9iEAW2nv/KoR9hANQYLiQB++J/QoRRi8b6cE5/FQ
Ywntpzm+bFDUmKPNmmW3m61kOrrNx8QkaF1mL3LNNPqd7JsWZr0AgLUvkfMHhh7dL77fZSYi9dNG
Rzaa13dInEfyOrS+JppIsgQajqaXyJp/tHDXYxPa+up91DnDiwWPCArFxerSer0R+GxFwqFt9bZm
p3wSxK105rOQyQ7KTxCKdocKWcleWWx8n/M1Zra6LlITvs151RddykJ+JDcSQWum1G4DMXqCoUhB
J1Rxzd56gClQflSWWMdWNmJElrH4CK9z6l8wtWtZRptVrWWw93GftzTcLJnDFPBJS83owrL0oezl
+SOU5c5QGZHrrSOx2gG780rG+new1ZFIGHNd2tU2ZlSbuvRyQiFxA7ml2EBGX9AH6GjhndbSobcw
CxGycj8iO/XhDATqN111wzVsBXshIyHvZd2AX9lkQyU0OozQZYebeV4pwDeTwlV8LW61pB+Z6uEf
117S56e4LkXeUKvxRjfkIlw1NZ9nGHOtvZcAiKgS8/Z8Kn9vrSwDhEJTVjuahEg/8zNK9fHemixo
FcGW1HrjbK/80HBiy6XHln70zVTjMSn+jZlUYGI00NIGp91s/8JufFvHAsOkUoMAPasawnc75ux3
p65ktzRWBkUYCm2YGt4d3zs0oRBNT5zr0xeZMy3nLRXuTClLRNhi+hQw7nU1OMB8c/cBMR5uforh
R+c/Lxl6CpU8tNL3UhL+NY24+ftsUQmXrQgfCW9EL+mlxj49LhJ26KqxNBmy+3W8fITiykKJ3gJ/
sEyDkfT4ywtk9PrVH6dJ4hqBDOrVGceQlXzY2m6UZ622l7RTIGH05ISv09MkhrscKNW+nzSyymps
P7qcopXJ25lJ2Dfrxq4n9OKuCV5joncE2qOw1JBIl5Rs+n33oK9gP6XVRBUVssNFf8+XiMmMaL9m
T9k29Edw8GW1uCeApMIkjiWclPo+zYSGD+LL+W3qRCcxQk5YbpOvs/+bEW/77psijs+bNCBUF+Bk
yAfZQuJb9tMTC6LN68bsk9c7606Bc1jWo2q29S7bJ1lmuliLYhzKOUhTldqDvQ1ixo8YyPH47yYe
OulwnUfVC7fWj5R4RhORSM5jG4HGujae3zOAjNncvK++LPr6pturudwDHgCQEKvir48iKWFfvKIH
w+R+Ut8D2HFDbCukkX4H0vd0TN90zKoxOzTYKjOpjFyBteayX+CxOJyBmkvJN+B1vOOmV3WN37zx
apMx4U9v+9G7THNhNI9TSSE+einAfyWy2ZfpaLIqtg35XvKZyP0mkl7fijb+g/oWZfeLhELy/DyQ
VsuFMErcYp0pxFuvmCJ/f7iDGGJu7/UvfGzi38jiog0Z4yFv09FTzNWciKU3w1iC+dlZt3xox98l
iGpFHihm63YRvmnOogEoVAJ34tgLk9sQRA1b2zLna8zyIw5gfoa29r7riHdeXlou3kcX0/G8fTvI
wel8e/fQfhudwoZagn+1WjgK3GaXsd/pl3tS6m+hs2b0hE9WmCMpIrbgsMRK2UMAP4vc04rrpufw
h7fkf0DIn0GJ+aZ6cup6gQLq/fcyPRJ6uNycTbPUX8XVc1xgVUswcioNAlJ0Y9VVcJifoh6ZPOwc
utBcCDs+JW52FB07pmaFqf9BISoeck3TyaUBU5FN4Vy8KDCuj4kgRRyZt7MS4RN8hr/5izO4I3I7
NyjnT1foOaJQYE9o/E3VWFjWltgUgS5ju4GPH5ZkiRuJykz5sO1zeRwRIU7x8cQsZl0x+gk6VS29
r0WFBoFWaK4tB8CewRORRDhDFax6m5pn3+6RgSTq7OsvGJJavdrn8a5CNZX10FGqh3RF1JrE01Tm
Ozpu8aYS/CdZoog5CBJv/GMOiyzcVdXhKR6vQY/MOiEuBGzJD02itn+UeD9DsAfuFSlA8naMmQQC
berkgB3Hacl9P/M2QHVjrISxmHPmMrbHzDXEG8xDgecmZNuoyAO9jcXKSAOQdS/Qx1fVw5ZodH2O
MhJYFhKRbJNqrI3IKub6r2oO4W0bW++Ha3o4PMkdjlTsFkxfilzqPFtQTLzuvRSwyUxYYW+IBkUO
aQwutP1Vi52SU5QFVVmep9dAmwJWJ1kDAicZcOL6smR9M62JYON/4sgEptTroSx9Aw/wTkQVW2pU
hGvEsMAL1A341Ao2+5rvy8WzLTza043pqn5hdVHBzNFEPRPS+eiZBtpQjDDFuR3EduQODn+k86F7
2yxqC7meDYJpDeuxqa1plTDszPTENofxoVyiKTX/aktNnISWhUivnAEKJ0JrDf1bj/XqnatWYrqh
MLd8n9yECjP0vLsp2fGEhHxQUa3rD8A22qPTyHzbWMY7W/jweedlvNuWUJTtthbBkkexQY6iV7wZ
x0Noz3Qa8nXQDzZaPp5LQpSJ8il2Pq1LZUCaLcXnO5unFUCAyvxOdP/05hTrkQfGXWvyDz3Sf0gE
3VmQvF8Nvu7BFeZ63pcCN3fQgHuyYNpyRXBLqAeoyxNcN5xAuRzg48XlRJ7msE5INaxiVvyZgRuo
NtbP716SKnMVgLuV3Aj8LtE7C97QTFQmwdol1Kmk1N7lMsc+51XxHyUmYMCz7Fv8is2GV2l+0bqO
CiT3WBr9Qh2apTSTkhI78/ZL+Afe1+hWN4x9kDYhJ/NWyLoqYHi1Hjj7DR3ly0tPhoO3CG0+bxy1
aWHqkRon6BE7+FpxF++qVZ/ygzB7rUKvTzGSf9ZU51IiJvhY8YLKexDjJm6Yuyr8cw8c1CSIAD96
M8NlRjpLqVkf5HZSpXB188EZTOSNJMlr7AuqBO4qxZFCcOW1/1f1/hd6dopKbB+bDlElms9SeG7n
xelAjgyH/hsPcz/8M2FwyItaAz/giUcCjfR59UaOzgNkeynUTtSc1RQKMW43daCurCG2n57W4aEL
YFMlEHilF2QPZHX8omy8EDL6fYnK/R1CT73anxIYlco68faraEtpwOmTIxL71ynBOrRgb947y/bl
3bDmZo7XKJlr5BmNvKrGjhUErxC8hUVpGo94DmwIxfCvXCRQ+LhegTEAk4EQWxtRJmqti3tTTUpY
sLrgltM7s+lJlrSWSweRD36vHADH/khmQrdD2Gxsj23YIvTLK0XztfNd7DNxmX8CG0yg8OLl4mCn
fbd3aDW/r7vx+wY3yAp2u56oY6eongLu0j5DneIT8TNFwb07G+VIsqrTNwgsSFAxD4atpQGzoMN1
+83vZj3GGK0Pu0S1xHgiXv+kJ2hDjR3AB2tIkh9lJUfWosM3L6OmVLaxCXYesNDmckLRFmc59iGq
wVGTctiB2g1ylrBvzTr0Ur9OcSQ34gi2yfc+Sr4Ue4JAYGYvBoiGKPZZmZa7s1qF9ul8SYFMBpkr
HQE2O5Nu0XmdL1oUzVXUtBXBMRVjh6GeG0Y10GoLNWF+TBmkyDJ1IZb+JaBe0J8XW39iY4LbD3SR
NFXvPvF2434ygjeuZgUEil0DpBQrr+Q6Ps1ybolAdOynsTgTX0eYnamEWGNrzHdCEgY5ZmqJgKXI
idNexf9eKJw6sj+aYodgwR20KCw+Kjg1GWwK3VbFVyCuL0IrdymHqQ3B/nJCZaldHedQSmI5U5ng
QuRnSZFMiRxd0h1M+giYigYYHOT2LUUQ5lEzWWa9SZlBfh5PN01I3DcqjM+GMw15qT78u2/u7xs9
5Sw2czCW+e33jOWWFnGrsBMbTum+cexuw8ol1yTiFO9wPMSEdxQ+cOzLb6KMpI1g05TQJHGjMZbT
1Wskj1+ceaxG8P6z2zwoXrSpKIZ81njG3pwXBQ7QedaVOn3Hby+O4nvTGXeu8oQXqmVyfa7CgUE7
FukU3AyO2eCB3PEon1AMS8zGTlmEBPh5ZYo5uAzMRkquBur+6DGWN+P/Yhd4ls+n8zONs4cV+k74
K9T5ZolRkaA34/LIdCKufeqP+1UEzYw6HD6MtuAC2f4PGygLDbU+Z9LBdi78BfZ5DX/FQEpgJTGg
ntdDWD6v61BzgjpF4lQ026JHvYmQfnwMP1UFxh2wYWVxp/loFr9TPJ92zd1rAIgkij6S4MHlqLEi
Qa3fzJ2koVO7Y/7alXyPmaXcJeh661G4jkHON+HIU7ChlciorzZE5bGPoltEWQm87+SHMYzgkw4B
x1y8jn+pMxx36GlDC/PiJWxrtGuRJ77rcgtipYUHpC/YFzF8gPohfffekCrcjjyaiTlQkO2PzPEs
yCdTmAc2yKr3pvEc69Mk7P7wSvoJWtmw7iDbzB55r+4X216Vktxg7JBYBawI5CVPEZT2MovqrCWc
vHM0Bm3tbd9rH9GEY8S5dSaZGN3GVjawX7xDMfbIbaxmV4kN9HHaLP4ODC0tnEN68JUY4sfW1LLn
FzYZ1FhUpsuq1WZoipJKJv4mUdHBdqh5rJS3tdw8J0uZ86dyB5NV9M5LkcrLrvC+PFClaDL1enEm
mFNUum9kcGr6CPNEcnUbiDD6UjHkY0+ZBFhA9xZ7wq8NJ+694HaPVYfztgDfnJhkogZg/iNfYJOa
FDy/mbPe9h7uPOqP7Z2/Gp4a6uKlF6ytTI9sCaZCbtDopzAtHkW6Kx5gC6WfwZBfW7DVAv4z2CUg
guLcgcd7gQwXz5OD6bS5eMnBWS9VDmeAWaipXl3inCjCYh1lSzB8fkqWzYjPjIm0PrrLxj8F9w5L
SEkUklJ1dM9WQ2tFoMGwbA02kx8aQcENNU0L2KDYI3EM1L2qA5Auqb3YcIKy2eFIWgO/Fe2utUqQ
XrAunwWoRALu+6Kwl2UoeERe1GNADxvTLanWVs5sUnW45DTCQMMi45MXnXfy4wleirB5AwrH5K9P
q1U2160fHeyJnunGPU7bP+IMgHS8H3R84NpJ8djMK/Pd5sZdSR/7emDIs/fMpTBnuyXN8Ga+qwWc
BybyIa+FglD5YLxQHzBxxgqhJfr2mzX0EeK/WeSzMejVmfWtFEPDSlx6ryOS3sxuwckZ+9REa6ut
20KK5vdIlMlYrhDb2ovm0Tmpt1bvDQvB2RgKnh4+JywbI67HyuNlpbg2v8/SdmsSItR6VV26D4Ap
RBagdAHkR2FtoUvHMn/hh37WcvC44RFcAX7flPU9eNZ4E+ciQFBcChJp20XyfwkQ1lkNpQG+bBpK
+pnYelcRCGuBrQ2DKPFVUMoFRXLe4rfEMmrx45TvBdav9oZRg8rp1XJHqXy3nZUEx4DUZrm1LTRa
rqathmt9XKIV9h6oC5xX1L6mXYVkjxJ9Mx9wjF3QuTHhS2M20D432+k0Q9azC9mk6Ar30zKZupTu
MHE/G5qTk+N8UIUg4g8YfrSVNH3J4brGdYyk18bZ0FXS8Dp7yY6DUWSiQydjwkr1TxXJGdc9cy6t
vIKMTYF+Kp6vISShDu6gZaQkTjOPTxQxw4gBJExzUsLWTQzW546cmv0kjGAzwM4Ifzvm4dQwyEPg
Dbn2yxoKfXODR09k/RHwZ+zox880z8B/232/nxrTaeRwJKaCXmd79X+U3ZENSz/yihejmpQRFWHl
QFlnNEnF9IqmTYe1SaQuz2mKEASoLTUFtsJ8Cm3TuxRt3/CV/J4fKzXnzu1u24/hvtDHja3H+LDe
hgUu0Zg9QxMz/GhoVGESs916/iWGi6WuisVB2PUmtzrRoodfoeSjfA9fYH0/to/z4bP/s5e2EYGE
9tGTgjIJQngU1N81osghDNBrrpN+0KbGHUbDKFAed990LQO+G7smC26it/tIVc/vHV5Z2v9i9seM
zxzUY6Bv8yM/jBivkdiY4vWHPvoLRX8JDt0ke7R+IHn11iMc4njDC5o2EaI2A6QFlGZ3UAOyKwQu
NmS/sxFye3dkjUZEJ4THF7MxHrumURrDnhwiG2ubpepRIsk7C63451S9APafMB8BnXCL0zYt41JT
1UgZBfD7QuhkFCL6MLDjm+fnEsziyCzmjI8T4WSbtBHYAs8qa1Dnq+tdXRRSIyKa1zw+Yqg3DfuA
om0bSZglPLxD5Tk8GXfkd7NZubGBrKGCETu0fuFGLaDU9xuRbDW3qgQy9C+kH/F4UWPElPPxas5c
p2n/YWSif2FBAky+PqVyuuprk8SZc2kDqEyNkqt3QPb9YZl9oAKT9oFrQP9xmsjZLeGR9ECic2f4
FXNKcAXSr4r1nHG6fd1KsOFLGazK6NDY/QUCPeGdxgIzSLrelthIXFkDCBy7c+8LLWGQQJvQidjr
iUvwWN9bT6fcI5tP6uVGHLWa+LqofsiiHK3WZk/MF3wYKceNCgbXN/IuqLx0brcJ07kgoz/JRSFy
BDC8Y6UT8vHj6Ryqzpon6B0Hhw0/8T/AGkfVgwC9hbkw0ckMFi32oMMsGhOoJy1Kvm/BrGILsKH9
YuKOij7owVX7D9wyem7cCG+xkYjuVJdDMBnQWLHM0w+mLyybhRCPNVAPIz6RHBssq6pv1dGozuld
K2G/8F/kZwjNUJx/399te6LqUV16UJcXdcdiS87gy+O5uRZnL+EHRpDqaj2Qh565U/MyVG4eJSBM
3ykGeeDtjQbigwcM0NosPW2ad7sr1g5HtwMvJFX9IWXRrm40JDuuwx/ZmcCjhdsx3C4doEd3MEIT
m16MCpoLBdIH0OfNLLA4Gf0FOd0QuxDSx8SXuPuC86xNn1dLMWDawy6A43oLV2c6oeL9MyOzvl7n
znQ06HR5bY4Je0F741dl1MGTzXsoOCyOoTGCTtQgppNDAWAqhNx7B+WuxXyxvQQVW5nYxmcHYCv5
xFIGhyjdl95thuWPGZ0EGB5eMFYYcZrhhYY8egq5wxIE3CItuNATa79dRveAKJ7h8R2Y62yzJr0t
o5SZtKrR6BVCXXWEeSOFoPKpS17rORrLHfoVFqTeTZJWErUBMPgdkh260hFdb+8dmS58pozNNAwX
rfHofiPF+mRkrXa9Xq92XUeDfNNIOe9XzY4BjnK8IxbGxRkKY1CShBe7yPnEkpJJPprcDM3rjdic
xkpmx8NCILZOgk+Cf9/o/uOZgqYvb+kiKpo/Lnn3dysUDkGNa3+cRlF9nLMpxWFVGj1DdLWlqkyJ
E0C/fBi/UO0xxFsoSMBptzn9gR7wJ5II2AIiYTSiTN1tV+KeMOyXuHRcEtvEhI8k2FX6zBu8ngLE
qdDBOa7YPHUFRD8vkzQ9Mdf6p7z9rDnRyA5jngsb1v1qHEPaS3pHloJlcjXucpGf/QtpJLoa20iz
tqgAncqklOJXBhBDOxr61Lldi1Dxf/DyFoHsFxsMb2Gx8cVw2xel3H/LwT1pHJ3kxTMNgPg7VpGU
LsYmbplp6qAg4bFsupFImjbg8red0YV7cHHgEcZDehnjE0BbpLcF9g0hf7wLLQKD6XdJ4cbzHp29
uZmUuiacNi/U8BdbxS5EYLHoKi0Mq4ZpgZ7sIAGEM89Gyz7U6Gxfolo0pXNeBPR6XMGNawEg/NL9
RuZ0x63rsLRNdyAreAj5UY3J/v5g8caetIi6h6zVHgw+3PiaF12GsSP2zfz5EsxHfYx1A3MKV5Q6
RT9vu2AQnG3/amI/TMbSSgXuDzW2GlLXi2y/k34nkVQMptoB5M5D2ujH8QxUFvfu85i5jsdgEBWI
jEks/est6yo5RR9dtsh84ezOcfktPjF6NbndCiVVEr7SiBrkcMExbMEMne7Z9vO9MlPgySoRUnuy
OH+Vi9L2sDHxX94dwodF7InZ6uhtbLk+L16L8Ge1BU5UUjHSeYN1a8tsFrB6wn1fKDrIzvtQ70aH
gXMxUmyyBqlM2bFWs83EcqOj52tKnLWPkHiYkWkXsgYU+/GiJv04TEfsJGmSS1m7NbaTNHRvBK1B
IjC9ZxunweUsbUEvXFRC29dm8xpXsqkKKAoWgao/PMybc/a9gu2WJ2fVRBlWVRnz1tmnnTRWvG5i
/Et188Oi7mLA7Rv8cRINT97OPb6Co7UwnrAq8gDBh6XFCFFzsryKgaDUXY8ky28A5zQTEtUUM4Ls
eyZ0XZcva4HthTGOk00359FAQD4ShN/YhrrRDAXjYPSW//xhc0IW9YsIPshAhHTFVsd4ADJXY71W
8BKnfzEpCDy4XqKP0Q0/UMyF+e1WupD9yZRwA+O8cO6eOIY44k6qRAsyYNynJ1joFvOrQJIDmrZ8
YyNHHHX4dAsa/Fv1UL8ruFZeSCO8fnQAUKqFb0OIt7bxZwQPfxzB23NPAwDR0tbK0hKOn+Ym7II3
b1aJFQOotf0qyaPKX4esnX1xQAXP5xHlDnxPBF63wIqA68ep4FfvNuXzJCrLpCRbECkML6KsmTzB
EPOwjs42CkpUrkzscC2XRKbUP8HgmuJGGIBosSe9H7v/AOoi7/9+gq0scZUQ+DnzK4NJbP4yLL/L
yXEar9BtQ0qAIDAwqzoBpdvM5tF/m3Hd82whPd/peqYfaL7Lax7siorzRyZfiJtyI7iZn6Mxk15s
vqWsCKuENdr3trxDtX+Z9gyoNTRRMUW1AaJxb3BUvQilbqt/M/rqnxfURYSZKvfiB+R5mPkcRWY5
soE4ml2fk0V2MQcib83yQAXtn1CJXmkEhIKV6r0ka5EjIFa6oaDx/XvkHdW60tY9GWo9osAgLMLo
1LbwfgHI0ctuBxNjxSuA5RPPsQwXV5LHB3ZNOE7VSUZh5JijiPpj6T5+Vmum8s5Csmksp5iGl3he
weBKaMFamOT6PiLdwJFPCPG5LK1duusfiaOweNic8taT6mSPQ9caIGwdvVbMddTIrpx8oMgFIvSj
UyAi5b+z7JKPhoprTT7SZ/0LeU0m97YIBhbhjp5DECN8EwJZSTOh+JCMBmQKHgKt1jYHShc4rl5J
qNgtlTP5fbmy2VErDyIsa9QvV0W8IY7+7DStdXxbPtseMQ2emL+ISYTrRHZiTPjdZB4J0z2ymyYc
ZrScrP9SZSlhfryuEyNA/WmQU+A1Idaz0FhmYDsGW8+zk8ZWW9Gj6ZzbSVNsma6eDLB92AcVnFxf
ck28Ll2ljZGR2FgtdXUvRbULMvaQgZ8PwKNE8UQsONrPtwG0OXAOERmbLE5m/5mzTH9EmxpX3Wy6
Jh6pmt0ObQAuOdM5Pz/vLQkIyqQ4zHm/2D8snpzV+Ip9+NXSZeVvz65oqCkiO5mO9uVWiS9Ar7lH
HaPEhnpqLVAm8glk9e449N7LjyM3CTLzfvPg9/OYksciHB122NtGc7RSTvK959QzrQU3+7FqQ+r9
Q3Pxfjljly98+emMXJGpeocPfTY3+BxTzDV3Y5udcPP/gj8e1Fro5tanP4nSVK6F+S+MMzZhkE71
YuDkVVlpwGRynwP3fQC86iobhhBPE0YeJKv7pPck1gM1mNGc4f+lR2ln+LZGe9nzZiJsOVl6Bl7C
wvgb7ckPPOdONyUUvYITyo+nQzGfLXfU196wAgZR5P8u/HoPlfU2cVIIcvpOivkS764XuAjQSLkM
eNBakwNjuXeusxf2pL49coUploFdLLt/ZNJEFK5MjGugFLPK/1lVvuCx9XoRL1tjCQGG5K4EdZS7
h82Hh7eOyeDgqn/2caLS4k4d4lX8n1xMymGi1xFpI7y0tS1UT3T1lMf2QDOB7EXEjEeUmboc3iVo
1xTjf4AY/X59StrFurlH3w9mULpfvphBjVml7uTd9QNE9xrAwUtyF7RyKYBcZngULptfLT9+DDKo
iX3RrE7YUJZN1WeBDNaJU0LhMpJbWX01olR5PvyYBwuagtVKDk5J1pb9YS2tKg6RukQ7/jpSaaAR
S0ZCh6RANSAegUisMK7xExUbxuKB+0S39rNacat8ULOXPYtNIa1/BSdUM87ER69a5+QHbv6Jv1LB
3Mb60k1Hg7hh2eUcQTSZBU4y8kgVL0GdfsjsnCbXY4L0am51uwx0o80/xEdApxNtJxEQsksnw+YD
5Oi/BAjsRM+O+kNiG/ubcVhDRlpRvYyxsFumDvpjFK8BNAFVl2mtg+IxDa3w4iToBG+DbDK33ieo
LZWFLsklUMR0huNDephHzIZUTrfIYqPc6woORuxBw8zNTbqXtfE6BDOJU2J3ohDiym3y2vPno8Yo
L8jSC0mBrX0jdXBDxpdht6w+dyQelFLFho2OZzAuOw2GqKUidzWsNQ8n1wSs6szYKGJW47Y8PEJY
5NZSQTaWq/UdBY2FLIEwWxK/KOE04hwRH0BBZMR+onInQOKRiEgQTRAgnW4zqM+jDrSLCY3NYjp3
DR6CsSVJMSwDhMayWZM0h0i4wGkCKQ+z8ahm6hHov76aTqttXpXRIPNQCWrw8ABc+AqGP4rDjiIN
xIM3bA5kR85eQeTCu3Ei1fjfpYbboKGYqYy2DrPp/jXORxePo2mKHeZZ9fdNmjxwJLoWfggFxsSB
oRU3l32F6DmeTix8rqfzrNO4/dh3veJNBfxdXGZ3lHfETdTQLM83JN4UtqVz+XC/+SO6Cf9geEzA
vlnr6JBRXVXLxFl2ehn24J/QuljxQdQXSDQoi7vOA5tk/9xOG/knaUqxTcO9598g/MKz9JBBzpxC
Ak9/pm+DZXwMLm50InjwzwhRW56Vh49A2bz4Vij/XmttFJbe43BcRCDB7bqevy0HLn+SE7e9EsU8
q1joWDTAJAjYPCb9FkSOKOU5mhmJxmcO56RIFp+duIDQp//ujOmlsF9Innl5/Av0L8XsSeFsPbst
iRfZ9e3QRBRXEvKBJ117kI9zKyr/B9n2Rbvr/UIx9S5ulIXBAOIBZNMth4yfrp7E1qo9jzH+Mj/b
rKALhCaAZnVkbjpv7IbWoPrEjmjqFvNS2msPpU3qRZYiSsaa5SvWxiu+0TkE5JBcUe2u+HEeAKdx
7dZNHdAtJf/qzWbTGhLCxHG78gihSnu64+Rj1qNIxmcuMh4u6FvhZoBhn/ulaVJWGkmoOEwEfFaP
hah/ZCTCaNoCsQcpaXw73C16QnV/pvayIIrntTzJFSaKXxziPABaqIWmULuq/HvpaXn5Em95MoEH
Y74Jk3ir/srnpV+iaJWFarfFtisXWhsaRTVf35/dosywSFBxSosWZ2Lp7Wb3O49FcxzIljHIVD1P
Ew5GYAZT8dzOgR3rl36G2I1HtjZY5Ep5EVAAq0MSNxXPnyjdFeL3Fn/VhgF/xlA7/hb191687vhx
aN4ehSHyb8fWQGCn/pJoTM1+LvrQQCW4K5aIQcUisS2FL9k/uVzvvy5Bsoc5nOh2JmslfDDdqsKS
vYWjtyiMK7x35/kJ3wYcXUj1Bh9YP1ARzjArs9laoBgPEaRGLPAzhc8zIjo2G6Y5Rp+eiARdr3q+
GOaW5EdQENXKDcwectRA50jVtUKp1X0YPO/rdAtqg2OxMAr2WctuFR1nKJwaaIkPVqPECq3DS+/j
vPlrmyGJkTiFLMuuxQ0M99y/9t8/14qf9wAzxOuc44p1/n4lo0GLJMaEogG7q2jSmtp1AsJDi0fB
7c63yxqDuID7hHcpYvwDVZsQH5Jc5+t1rqHUbdVyeqsbvoxuDucguOXOYkNSgE6z1rTJAWJMveI7
SGJI88o0ZipYBJs4L4KNAUOuZqOH4b/Ofg/m11nL1T8kKaETshPg/nV0CQd7TGhjuGHLxSPCD7bW
a2djoh77sTgfg3N6usFxt2xjyhuWWjD+sCWJU4X2CvSNicviIIPCgOy94bi1lF6dEbUA23tdjufu
5vvhrDYvkfYkxKvD/xBvSlNSGdRKswLTX7zZoG7WeKN1SwmsmZ6pF2oMl+yIFP6T20RImYR5ITha
FNOktYLY83RQqqYjdHvTeMdVroLHqm3+PFqG46179R4R5objvDqRUpyuw4dByd7QF+PF2stsnVSl
dM0rYCfpc24z3dbjLE37RB6XXRkFIumTLdzFthfmGyShUfxCHuILm1dqigvwn9P9mP1XcLAxroGY
MOs5mp7VKKyhwsySnJmYs5L2UgNoePDUcKV6KU31gJXjnHGjUDX7kLIonm8NpjXLM31mf4vMFuI5
jtep5A5vDUb0ukGlN9tDc4WIM+NuvAAE0JSixVQR35dPn/W9oQJ6Z+Uz1fQJMmIh/h++27imLrLj
9utWBU06NcoLi21ApW8bvPwIwEPYENwhz0oLfbHrY9gNoifEhurPgdfnXkV05rXpU/+me2SGuezg
PSzE0oodl8lm0c1CniuTik6FZeUwLI6Ro2L56Zgyu7M/RjGnHDOSMHh3mfxdqErCpF/1hildHkVv
5RNXJPBD0ZpvA2mAFfkw3W2Jc4vVWkTqX/NeKWL9WnQ/uHcJRWqbxJtp9YDiXh27TONZ9b9hSXbB
iicM5ks5KQb+Oocw7KVqmbAh7FsOVMUQ5fAJq83zku0kpDzgskSlZvbqvCTWY7OrG3NP8qedCcTZ
lAXiow/YH4qxE+ia7yOizVFgcNweBZpimgVNB3Y3LnZ6CpPr44zQeJqYfyhQ9miLil/r+o+QWiUh
uXNFwTE9QMuZgUT2Uqbyw1O3GHWg3eH/ChILPEG8MaxLnvxt7uBXHysuIwIVZ4/IByyRNaTkeq/S
xPiSvhCIpgiSPhWoQ5Cc8HyoBi225pZX2ZlaeNsskpYr9oE8nW1++rZQ+sPb8B67otLuQb9OtvjH
SAVBUqTDd+ae0FIaOodnh8jxXKbIIyKz9Gre+ctgrh+GRxopZ1d1JU11TuRTDzT32Z1bvKvLHPDS
HETETHJdmdrNUw0P2rp8JVkcAA3OjXobO5ARY4Q0+2AgEo4W77qSZUkaD0cymyTwn/HWTeaVq3UJ
WjbAuboRus3Ll4i2nImaU0zT0m7UIFtu7NEFZOjv0wpkn1f7CmG1u+gm4yeudjz7QwSmKwUA0Xgt
HKRqw3O/DwLCSpIe7p0o7jOhWXrBHrjotMGA+oftlk9pVpG1iQ0uTnymyeB4n8kJe6IDMPVcvZqx
ndiPr9tDUkklDmvWJFxoKoJWXIzlS+ndkUaETibXT4q33Qy3vGNbiVpH0+lsyKi2bXScFpjI8jg2
jpUzFWZoM8/xpJ+WHCGr6DCZzKejjgeWoNrH1g4wy8sfgzixveGYAR0mtkF+VlcF8HpjgTxmWjnt
i6G9kCxBw+YuKRybRHFUkLRIBSnKgPkJ2zK26h0dO7wWEa37Cm+uA8OuaSFsBYOQPCIJDao3Z4b1
i0ns3hyVXbBMV6mXmYMI/+EgmDHI/4qGZkSNpSIrqxEtzlIdK6K8IccvqOQAZq/n+zKk2bCUMstH
rIimx/JTu9G/zvAM9OVms7pdkKAPxx/Ly+XdmZooi/kb7PpPVj0fRcyzpu8J4hQxlr6bPlifttw5
g09/fnrnP9jt9edhUeNTVNmhz/m9ljwC7U+RqnQR4/zd4UzOEgvpANXMoAAwufYiqg4RKQT0qpzc
NTk62+woVLvyjUZg92OCVie9iwqrhn/15iLwAJWGrNpdM4MxXckWrBQH3M92NgAWOZRsBYfsVgot
BgUewA/46pH8vY3GEF3QhfjYzONFra01nF+ZtGzybWES1jvOBiu9ah93QCcL/ari7K3tvbkOYpT8
JoH9kaIzV+E73sd6AuB3v5DwNmkq0ZZgGyWzcAx2FefBqzYB3UdIRWTeyTdbT/vKCGjP8YCM9a5C
MoLZe2/VnKp45j/Gs6Pz2KyfLypZywp5ua5cXVoCli47QyGOxvBbohRgf/pf+H1c2JIuQXntiKRO
xfiz/ZsM+de5ktwPQvz+3cX86/lFMGeJJOa428f4Jb3qYU/iYsl3SXIvcLatCpNSyt6CdAO/K9/r
qjlXiZDiSFBaI8oDOHlw2Td02NyD/29Elfx7JxupXz0AtCJrGpDG2lPXmbtivdM33RRjEB0osMb1
G0kW/vYiTBYacsWgGlgKlsWcELpwl5aKXj+WOGj0wZ5oLT9uZoYw84PF1BVm4o16ZUwHZiUF6GaL
NBtlgjGC6LyVAdLoekxptNiEHeBMhUyyr7QQu5/vEmElXZOAMGi0OEXYZjzXDMCw6WqAT2pqhIiB
Pgd2CqrBXIZsZi7ym0zbqUzzZLNgJ1JxRr1v0RTlKCc/RAT9Ttb6/JMlWPVE5rPXAsFZXP2t3J0s
iA+vK6Y55MrKICDDgoeGqt9J+5HygmhBWOhdCt58TAt6aOuEmT6sGp227yjb16cfFhIgTXnkMbZh
AhS82AcImXCjgPxCxkPv/Kqxj5JdE6aPAhoJFE1AGgQy7JM5AVGNAVveceFeBaobIE2fAGEQSYdZ
FhTE15+DNkKcoW1Eqvg/i/t+9uNSIWtrvZ0KyaYY5QlktNS91IuGRKlojTCrdkjcxshKcU44qeIz
YHtGhARxdOThFFjwaaZz8wMzPTOpLrt5SsM/mVxdOi6OvBdIoZi6zPB1prHnNsa0eQ2At1/PQBAE
mUGZtrq2myD2zDidwcmhO69DaNkdRc5uublqn6QFH45RqpStI9I7JPro4VUoQE14A+7uceNMYUJO
0yT5A2lH7mnOHNsPnqlbjBp4qLmLFTVZQhgnA3qca2D6SH3L+mpBJZPNRkX6OueLYcj3Cq8GGPer
a+DamSP39+9NlBoC4jZ+FLpHtFzLtWWyLgpPPjjYRHROhiDcLT+OXYALx+KwRt1288kSUICGAylC
i+trrk9HBVkjTTTBZVDje7Mw4/LQuViT3KhQ1jnjG8AwSB02pfvOitsTz/o0MnCjU5vZwHfcuYDw
9Bqq2NcCoqmehA4YOks55rhI27FM1P8ARynicuxL0cG40ipi980+5a/k7lDycMQVLZhdS3ebBYBB
DRaDQhOvJwQa6sDhbjk1cMS0P/bNhvqyThFaXtFTB9IPXJ5yT9wQsgnZUlzkWSioLxDEEzgmlu8o
7bxyxkwMgYMZLIm0n0P5ReoMMMiLWSRzFykMernUziPTYJShTlIpe2Zg/W/6MrwI7Eg1IuTs9OeZ
R+rciqdr5wBrOnJ9TktDHA31rpJPmH5FLe638syDkgIK5i6UK71l9cCOPRKpoRYXWASEm+r8Zy01
joC7FRAMl+djC1944B6F+7K+Gx8NtrCwaC2OauxTrrs7Z3/jGOvHvDPBi/hkL2mVH3SOfIP6UPFP
l0Go+axiNhkmLiIHI7/IxgoVxCbtCVY2CTe+LwWaWIJrh3RFVmPfrbW/+5lKHLRWB+zAtGzshU8b
Yr3AhKUuVscPSvhw8iiuxeBHSMeZ527isi1B+JOGY4TWqDk7seJIBzzLpMukBVPqn8raQwjnF/Lj
jDUzMoOOQ2qXWQ3YB4YYkbslEG/I2OWpjt9OGeBL6qlm54MUiyvGvBN+0J/zm0TBP46AQW8iBW5B
SXTRFJ3TdmUcl8CVApVwJarPmdEvxIP2lTHZZcEUdhiIfNh7VkDuRiDv/axrbkQS/fY/ux86Wmg7
w2fszus3nFLbFbi3ysy8oemOK4MO9XIferHHHENm33iLx2ICT5wqDX/kWaoNAPgph9QJ0mZoQZzT
xNbasVB7IpM6Br5jOFdcspUzT5bjPF+ehpzoA4Pk53B3p83XnHL9bRkeSUkNBU0mBl3gBOmKgS+F
KmMOEIZVVO06bopP/fnsx/5uOI+K/L2xJ6EDhUssRlpt+1Xm9UnrI/bqxK9MzBtyuZynDbz/NjUN
OaB4OryPaxKycLZgPqAdllf5DfknBfDLGaDkHsxAVhh5WW8qz5x9mhf6w0MkQi3QLqZiau5hqqL3
4/0pyZZrRAXwkLDJuH/ohwS55En5eeqDcU+U+izhjn/4Yn/iP3qifOokG0DtQ/kmtH+YjPLKMan+
sjiPAOyJk8Q4lpTlyVhNZUnG1rbG5/bMwoK2uL+daso8T8qxRSsb030L5TPw70oUckH4jzXw4hJI
RDP4O6dyAsnyVEOhXYb/b0EwZTJhBWnIX9SeEJ6SPYU3m7SdRg95v+deVAyNRWvsUR/ebtzteNao
hnayJbTqfMPygse2tU3xO/VMgtplQYA2jIkuAHS+QMk+xs0z61SmMogoc8xc4EmhAHlKwcwPB2m9
PjXBWDtmaHNpzOojU7ute7HWK9hMy+Xm50FZqi7UGHG42UAm58PUyoqmfr54iBPGq/wvCmcGBPEV
3wsYZGYS1h7pZTekE6sGC2ApcaYYgCMF/cxFTBjR/TCCYi+CBFNTCYRobQrnq0c0MZogCCPfsKp8
HH01X8iCPOun8sGdIN1sY3y02jQZWxUtfAx8LtD7ZUPHEzfYSa/89SBZbakxE0VPVlulufJ8Fuee
AYQ/MXT85PkJ3fGDw+1fM0e06khQaEr3GL65r8X/A1qJyW4QXMmGsTRvB0VsVdd0FFukvBlqLJWp
1ilcegp0z5SNqsfgtEG2m/e14SBCrYWugs3lqprtg1fHwAqPQUhmjl2I6aglbNc2skOlUSHHZbQh
JHtxmO1jWdXJfnTyxkWSPqeETlUIo0e625Ls6QBu/Abn0DTTb7CQYwnYskcmm6gMOYiu1YUMnqRK
ZEcvgkP3lIk/+crW1UMApmmnkM0Py8AGdjFjrVAv9us6SR7quvKMgaKc5OhE8dg47G4g/GsEXKur
YDLqsp4rBjXFuUY3y0TUZp9uT7Hdt0xhmp4YJpxZWYSXNCfw6SKbuzwaP9GfUoiDHfMVpP4ovKGV
vrUgF0ZBvy3zse9mD6nP7o6xTIk5qUJvtU6CeyoRwOz/ARECFZysWdW6Ebf013BeZqJ7vJVJd/hy
Dw19EG3ONgfP0o7d3KZHR3pCBtR1ph8JV5ROrWOSTclMtwFhXuJyNSj0dlKcP9+HBEr8Q/q/7HRf
V7RKjHOzP0ixyI8dJWI7xpmA2TwvRiJQbSIaYC+/e/esg5oZvdVVzPBahWuDGkRbyVVu2fTdZi0F
TWy8c69Cpf0XIIY989yItjOrSRU+pYHh/s53BGpOi+tFC1z7M1QyxfK5t2PHdCKzMEHhg7dbS9Xw
G7ANw+XutOAlQX4JkMpgNCWAC1C2fsdn6f8eIhEUfQxPXZ49Rt29FYpTP/iR0CrW2KQwDZWs399p
N6yp2R2xecKTjr2tuWjRaV1Fgo/fkxbOmqyrr7Zx53qUCC7s2rL6E6WdIgpHyvLCS2oI5pww0ey2
xu5thiPSmSr9TaMd5MI3pRrVffORK9dYqPkD2wPuy1ZQW3mnibC6zYz/z85NEuoPF1L10mA/uw27
k8LF4DGzHZTqjNN7IVh8Und3ef8DsSLbh+nTeb4my2RAD0aMQwFZPPNo9LtFmWbKBYVfoSBsnmqc
e2/89A9/Mkh/uB7UJxw6F9KiiaL0iXHvGXrb21b/7gU/PNxK1MqUubLeBogcOu6OkIkkgkFVG9Cq
QEW+Dj9zh116vGmpwsv0S+kogvmrR3OCsrpHjB2wmtLkjlFvgd92ronJHSsr/ZVKhIaGeYie1iP3
zBePO9RVhJ94m+i8nZ02TyzYJrLnBOsZkPetkRwet6lDKb245EwjqhPhpCkc8P2Q0WamP18bu2Z0
W9qCe5apo1XJJVa76gUgIRFY4gT9vM3uTw8NLii4G4xbI3OT+44YmggWHEooZvcbZrDr1w1cRgeI
WFk8rhdRsCuk5hAbOjKh9mTnuLp1KNveLy7lWY3GHFYyUmuj/scoM7Fm7xomiYBwWhBnE+rTZqTN
AwnHU/1e1GseIkFd8ntbUEKvTNrNPkDwI60CTbATIqEUV+2RxgBSQGfJaBNVlCPFyZ4e4fVyS0O4
xGoScgnVFs9N5qJCdNAKe3goUNCMACOFHcj1vETGa9rlz88eueOElx53IorrW8QsJHPaUZ1KEX/F
q6FLP7CD0UgJLNRMUF9l3ITCStZkCE+9kXkKw1UKs6/z5Z1lSWlb+R2YmJHO85mPqP2GvY1CDOwN
/+0mKrATsJlDxrrUjl+0bu8D2pV7iVMo+O3MMGFJbjyl1QhY539Nrp2dS8pvYiM1gDz/V7A1xo5N
22u6rHKEXQZg905NU88w9Fte6gysJl9w07sSzPOu6mUTcOVoYNg6DHLL+e1bYm4NLkDm7xAj9H7K
xZuifMEKrav1EmwKVFWUjsTpkHmqMvUya+wxbCeLQYO4423UIeDNY1qCjB65j/podQZ8VIWflmvV
i+QQ1crjUuNU81GbsbJDUr+Zg9BkxztJKs6TwLVJCPC0M/qlJMd/t3Ebu6JebgwVWcJJAmAyiKqC
z1Dl7qDCwwE5gQQnuGC3pLY4RebtofcF2AxGSzaXHyTubrj6Z+B4jv9bwG0YA9OsWfNoG84xgSID
XzLhmzK9jJnXu2gWMREhNHJ6yMHjoZyUYHADYMRnG3+HwzL4tkLuDklu5dBb3ybDRqQ+oCOR1VfC
Z+O6euq/ybtQncpvf1Ko3SobaFBRxX34uYrqKa9ADYAL7/MBahSqcyX6yo+0/3YJKUOkzRNGXTKa
8YuHgmNXq0itZZqEsOO0HYQ0a+MD1EQXvzN/MVqWii7S+olQEsBBXeEH2WhLPkJbNIGA/YnY8hzv
YGRJzFQeFWuAp3jdC6AwNoDB3YQwzOz2PSxtbp+xcDMwgmyfNJYSZ5Gf0gN3VYTciJ36mOoCOO8M
nMPjuOCNOklHmHnL5rSKcD+GjPD4JXF+us3FKsGU7+wMJC58L5nnLBfWItCBu7YoKwb/8aBEuivh
HoYSM1m+7anb+WL7qejebUeDAeb2rb8lkTTGP5aCgp1h/nWgTygJxNUP4uYAECE/Kt16llAZdP4T
Ab1kZS4bqelLoJ86uAI7j1/3uusaKHOB0Efxy548UM4+utBIGr/J2a4XoUzC3jMZ62TcjnlsuPDm
Co3aEMYa5dlfl7iyvzbsNX+flulfIJncjnZvIUXKsKWVOkl/awfeElDTme5R2f1yyy/9f76IGFyR
HpgsOLLlfQF19fZjkqQ0Qa7FZxUlI+gB+JgXcRzIgnCb9r/4dQFtdzFGfEzwY9GqoYRzLI36K6PJ
WbU84P88Cbzqjp5c6p8uXJokK4Ft3WgluoZuEG0lt17nG6CrUjAxufzdJImLQMD606ePBWJo1sCY
XiRSkmXm/WgqhNQyV7SVMpzKSW4FzQxsA2WKGtQHFaY0WrfGYSN7uGkOdoXSeZOf3jqnRQemho2a
kwV9ZQ8vgCYvZ+PCiado7eTRUmGFVizvi/QzpX0v24VmRetHUeLDg0GycRmsEYWbQCeFbjuezenf
0eOz2Gq3KmaSR1PZGN/Rscd5oaysZcX25Wze5JMpwLi2BQZXAy+3eO7brJhW01swbkecJ/N+nSxU
QJ9g+QEWZw+JIirSt8LwGEQAtlvELLwKNcGg4H22DYaGX8QCvVLGePaKuBL6OveLo7V/PnI57TyV
5/9wFbFAy+NHkqLf2MM652V9kevXgIEEgdfsuL+NtUImewucchRmFKI7rEBaMd1e8yVjzaMcXiRv
qyDyZYLQatzW2Tg2GIsK8muxhBgBCrYAC4yBU9d5H13fBD6/xtinEg4o4JjwkyySXwP9TPSXrlxm
LecBbC2EfJHUXl9MOak+Nl1bxwmIKTJ9ReeZfElXXpJMRjZJMKnar2P3xZW/6b8ySXZ5xMJrH0U4
EzusO/8PNqMGI25qGykzvtJ8ABbNzWw4Z1xax5fu6NRpRA3Cvd7SZxZlvdoueHmZ7tThXTBCG1Iz
xlGwbKUj3yoP0ubwMOm28tVNfX+sUn2Uv9qKON9C47xR1uIZTkLRAuaKbt7n2Y6K9ZuXpMZtsM3A
JHsElP7hxrqUCeQ/efd5Wy4QiPCQshXEGDkd6YGbfne95U9D7V3K7g11RdUxzbAkr8KqT4Kt9HTh
8xDf6RbAIbxGE/AKbEw/t7ME5Wsw3eu/OjkBwSIAagXgRKGt7H9sfQ/B1Aa4M93eD/SucmyT3JUM
+4n9rlN9vM69PN3dJtfCWIiNie7sCxx7bM1nyKg6uEvSce4lfmX+qTWIWBwVOkY4kH/V2sgSoiqk
HSRYmmciCfzYbViNZfwZjz31TzzlShrmeGk+0kb+CVrXrY+guUgAyK3ppD45iOex2Voz0OaTBQkl
21D1zpNKL7p8RrD7ySG/iKUX4+Zw2ODkf2xf+Ra2cYHykbn3MUbX+Xx4CNOV7/5zwKmItmYPb9Qh
BNxjyWtti8tphV7BKdF47Ha+HvL1nDxj2nR1TaFFYsbIMXQ5KKF1KbJKOV4B3S5L7KIJF6AXqSxE
h91UwOouWeqK8WXVtSNvX/DmUB5y0+y9/fLSfiIAb/2VbsubcrsP7awUu4YAgR9A26asyjsvMIPb
p8qrmcv8Ro0W0yep8YImOlqPBtI8xFnsKGomXrvCNGeREESdAIhJqbLHKsB8sZSC9ocVaCCy7iNe
wFzDvri/jKJWZGHxg8704iV9snBwmHw/nX86k/diqOGoXiC/RlLQcZ2madQfHNxDMnZAoORJkS//
1vH47LRoe4F93/noLDCQhUTOhCJ/0PjN4veo8Tj+IDoh8f9RJ8btYV1UNgrHWoSWbk2Kiyx4qfpN
O0hCcPPzWHpRSPaNXo9A4OKI5gM5xSlI1f4hnUF/ts0ZDxNqL106yAwjIftLNcCKeepSBpz6/f6I
D+8SoF82BoaaKZzTy4fxZ7kX/uywxzpTiNNt/Z86Y3ZaJoomhmBsin0rOte29voyA8SUIT4ivyrx
Iy4uSbkwljG4l8/RReqF1FkcsgKamAjzWRH5aT5md9dFOslX6WyCTq898UsMzvU78b5925vfHD5r
bi2Ah3jNpzJav8BWt4M/cCw0SXNQEYGhDgwJtUecMzsEZVSipZkQUVqhvfGrGOtLz4ceP0900WTZ
2iTVHGU+DS1Q04IIO3oZbL+ttsPIBfIOz3buHs10LGdTDHfTvyYGoZSnisEnaE8Sc5kOH82sb4I6
gpNYrbcCC0+t7mypNpmcSBt6Z7BoUoETBYejP23sjEHczuWlIbDe0bMUDHLx8iWW8ej7rXIPx874
ppB3VlHs7NQLa0jonPBA0tWC/qNntZw6+yQ1sklSUFnrSqGeW96Cd65VU6xOrk2y0DvM1ncGWsW7
8MTKA4aWuolzAPioBoLzth6y4MbPUrTVv31jChCGL9Ep0afG3a/FRAjKkR4nnGIJLxu0Vg399T/X
BUPqUBaX13EgG4sm6//zmQIqMf/eNFhTnmrd4OZ4qtcn5NseRGZ01rzOcCB4IcvfHt21ZIYhrU2T
VeB5RCtwVMOcE7dVGG5Z2eTYmzxf47Q4t4mLjSJmCxGucZa5hdEhCfTsjX2OigGEnUphvhVBC4NR
Q/7B/wHt6H5kfSh0XkASL01xhxIlGvdznhmLsMgReFAMq++TLyaaLsLcEgGDPG47h4smms1O0ruF
+vjV9t5+JPJXzjLDIxd1NhdW1rsvcqllcqwgKO/uEem2J/5aeoe2RVe8TkvWgBcIK8VmEaQjWcxj
R6b1LrgQgd1e1FlRsNfwOd0YwNr3f/Mif2W1YGU2M1D65PMs7xn8R28zmkUTa/DjWuA9Ts5XuweA
jnu/CqRRc5Z/TPHCxx/yBepLNN91BPdKQXDbsjMBwZZESiyWXrIQaKldgt8YtQxCDDoT+hhNr6mA
iThjTwlWBNWIqFLKpDT6XWiOUN5uz3kLtUug47+lxLIjD0eUyloZ/OA87ZbmunSrgMMZx5D3iadE
B3lr5Zi4Fz8OK5/yf11kcpkJbB3c31h9j0yEW0/izpnrwFwNVdD0Oh8ovRA5d6VzqnxHxZpNZlNJ
uEctb9tkZJvh8YQIzM1Xig9v4AhZkh+HEn4zx/52OuRplipkQKnofV+4zs1tkvV4v4dJxLNJYKEM
isfWItQYyQFBpeaSopvXIUK8SaYRL3jDXiBzloLHTtEDrq2LpcxmfPDlOW/9r7TM0xJkx/AZpUFc
TEmb3llQM+cmbrfY8XZ0EVRM2yohNhoS4GpTZTRO6KVPtTQO2VnlrEZwJgEQWhz3gl8TxVFAt1n9
GFcbZk/11UIPffC0Kkf/vcW6+bUEmI4reznNzODwNxRLPTZK9ykQwdOCvUiz3byUGxfSTF6sWyVU
/TDme8/FHNSWXUGizHJdAMei5A/yqxrZH+IdXIWrr5k9u44dgeEAGCI5tPiMOPuCom1+9JzNWoeL
YgmaciCWsDI9qhoghIW3y29ePyeg8faOmCn+bPcVtq4RQk3W+x8J4MKS8T9L5TKc0S2ysEM5dNxO
0/tdChwzimBJ7kNtV9L4NQOz3qzJMVLywS/WUHBVjXgpSCJRbzOzueEY0enNd3XyzBz8+7JfCEPg
1hPa7Qx/M1ZQLCZDAu13u0mLOfMjawrxLzOLMSlP/bjuou1tAm9X2DCtBZC9hRYCtXBSQhxEvxB0
Y2T11/iqAtzWCLN49LZkdLt1U16yp4qmaUH/vQle4EGb/V7QYfCu5Fjebc8+sCjJTnWx8TWAmTav
/MT+YVymcI/FqiaQPTjWyQ/o5RPwq6jDLNghxkO9ZqQWgRQbVJnzPULuvmrg7X2cZMbRrUMNkoaW
qrXWlPBLsK6nhVvq8Ev6mQTaPMNKZ/4cNGydfqY8Te8Yh+mNu6Z8N19irr0YhuiaPpYJnjils8+B
7x+CJl/zgmY6b2Djl2EthrdJiE0SHfoEfRB01OXVR80ZmlySdyF1GfkEOFjOKO4RBEJCCFSXyG5k
C1NzdLfZajkKahr0afL7h7VgezSPT9F6SyTUs22QmGUD+iFINGRR5QjVKrov331fZZprGBvHi0oX
fuCj1QGJ2j6XeNgXlZw5HSQDRizOb0EgYMP8lJ3Zi+lOxBpyNPgBwRYaxjHK7jNurvtvUBMrqCBr
AoJbKSDMij/kQRKMBiImb6DBVmFfoOPKfz0+9AmEzL5j/jcMVrPGAuT/Py9H8zcux7PfIjPOoj3T
Rka6LdI43x1lgjR67Y2j9xhtPElhI7LIm2iLc3oNLMfuQbmUVIAwfLR5QU0fYUtwiqd9UQNTwGri
Yydj+Aub4px7jZlEcCrj0LmYOAXnz4cBJvDjdOF9jE2DzWywW8L4t23BuysfJVfXiIIQfyO5LoFP
gXMfUVRCJLmu8HczzaTUSZQSLHP2ZphfdnNG8a2sY2J6XH8St39xNioDFPJyKO4emAxnim/iQQzS
MRmWmU6xm2MH38VE8DL9NW6SE1CODwTVAlD5nE3l5M6qmT1hjuGGAUXYFjgA4NDOBBZzWPwwmHY6
zcaGA6/P49tQUx/22Sdg9KZVMkqhb5Pz2Hq3a3vjuaK6Oy3LqtBjwFs5Ig4hdmJX2HSxMy+HfShJ
ARNoY4uoTviHP2onF7SfQHrWO42yitQ2raaV9BVFD8CD3dnhxNAcoI6+EqXTCFWyDWQ3npiReTWa
pw0NW5bgsetrJCnVpTbAP2XCl3p/JDNzeaOQBwyZDQ/wxvJdzXpewYmDc0dsCMNGgHH437G+sJ/C
PpAu+ySx5z65KKP0x3GHcp3KJLYyB6aTpQd3+UOMX1Fz9q41m+Zj902mOnCvpPFirO6E5jJm6Vi0
VoPBgDbpffrlE8ALwOHwmD12H+eDqntwADH2HuWruPGb3GwqmMeBKzC3twOupE4nV77Md2uzFf2x
aM0pCY3634Pdi24U94MgPWP7kr28ulOMMs1RUiV9KY1a4ZF4BS/ZfJYOjc5FcqlnLx2wMsBM9sPF
rZHaDoOLU8IGeLsMS4hhL3zMCqHdgJbY0/2QccYp99uCjED9KuQneqv8pdKA1DqXNWyi42LwIE3N
yw+u5DE5J4QcQ7Yq/GYQKMLVMFztwldzS3I20V0K+htroSyCvrt36VzCwhJrNlb060O8eovqgDZ9
vMLY+mp53vJja5wkLlTW59pdGKdyt7FEz2FDoi96xRw++H57KvYAaYiFIn2RURmirZCQpn3FQ85c
Nf8mPraWuzhiTrtjRqcnHNj6FMLHUdiBH+XSrHzbcYmB3/wA1iMW3xmwxltvxx/7wJdqaLrSjlek
dpyAKdOEZu2Y/mBy9XXLqJm1BoOt47zGrrN3COm2QbxZoSxbSIxByVOfeKxUg6PvJGMua2o4Y7y/
lcY8rdpXN0MvpgsMdCFeH9p+3g4UTI/IKMmj/ov2qC/LhFIKcAqKvbVUU21eu7OcF3ReEwIF/8US
BLozsfn0f4uU1VGzf9bGCyfv3iM4k1Qm9ZxcyNDiUyk45L9q6fKWTRGOSEiqN4PGeYd1tXRKkRX8
nxh1kKHAdMuiF7NlFFqGxl/qoKqYwyNJ2i57fZBiRrDRo9x0L+XDMHiOJLbuVaT8HlSYswMDYknU
/+EC4qbFDzynR/b9kZ0fVZGyNk5wrBmGwSlMf5xq69ZNIX2PWRnr33vdNj7/v6QaPpHEUHnOn3cB
ANfGtueju/IAArB4yASRKvJgGEu7kBVBop7IrSm4FI6FAurM8G15sx6wsGIYbv2bx79x7Fq8go7i
sei1My4VMC2cyHM2wcInhxz+mP0S1YW3hgO3yPgBvGYQ8GTTpH1RuSt6Om2nDQduk95M/vJ0cqIk
aObloi7DKk6Dd0KO0ea1vy42sxLFB9aB4Do5jQ+diN9CZm5ez2RkZ5l7baqJoQ4oDZzh26sn0PZD
gI3V39Zatp3FeNKoPgwt+gdJgpKk8HejjkxtGeAnH9+hJZHOphN6U3IBl7uw5QNm+6/FZ9EklMf6
dXV/0yLJEzbbgjLXUiv9dw+GEeYhhkUWRUqW5R6O17n8qpavoQizzytR6actsUWfbumh+HPGgKgS
sNN2ty/u+b7d2eL428MmwkZ1QhoYxM9WqfXMMJzHijrKKfjDdYP9JPCU7LiyeSSiKWJSQKb9fsB4
lQNL4ifq6FTWZDBVNTNp/fOx2yi7lc+g4yynav52xhfqUE5reT7bHnZdGmmwwu5BrbUonv33rDps
U/4Ep9NwqJUilVDPaObg6/dowCC3RgeGFg3Lr6SuhxXcHZroXTA6lEwEcciFJGhCXo7B8+WTc7IA
3QvHpCnioa/HnW4In6GAA4uBJ0f+GPloJqHL2UHFyz07pQN9wRKFD7mikggah5LvZi0xEIlixZzB
r2RjzPf6zV3ZrzPdpUElp5+qG6Xeom9dmkMS2nGqpmAQaMy4xZiyygZDLm2hiDjoJBZSDgWerDDU
5TLFYV4drD+fzYZ5mw5oQrajPA8bsXqNoB1S6edYbzAQWon6g55xMo0pF4cJ1hYYzfgiyGjkntfm
Iou4mlXlx0gzoQe4k+wxqsTG/tCIXNtZ+o0QxMeKB3U4vAkQjBECwuoaL1zg+wLpA7kdCl2qP2TF
pCVZcGEyvtX5TZm5l/pSAW10E2vIz8h9HbIF4vLYhcDx/seEfUQyQnqHzTzvEuguJi9q46LgYw4E
97GCnNb+7+WM0EOP3bCSbuI1AbyVkYd/sfskgTvLQYy3yQrE5WNDt9ImzfQwSx+bDZRwbt1Rwy1x
Cwttyofe1P5fCnm605vZNXNOYS/55Qo3RdeqyWRb0s9KergtnxB2Dj+GeLDTK4HMn+SxPDsdHhsQ
8SHIXZJ+6qyxQT012HlPe+co19BswvnLxT5Z13bxS5B9YynHvKGtw3CXY54BVZoRhce8ordKlsWp
X8l9vd4ZVA14qQ0e73sQ8fc/CTi4KUlLsgXrtG3Jfkk3e/WC5RjwZtCme+pfo0sex/Lrg79FO8oJ
XuyNV8w4bTBdkhRA3d/wHvM2b4o8dO+hcNbAE1983gWH/OBgZeLyqbFB1LlwAKjVS/p6yfyCHvNl
UdROjY9qW8bJ26/H1nYo29smFy06NCr5PRrJJ7dTpweItMtkxqHsoOTun//Z0kWuuFANwnd4MRVa
i308bJEAWoVUs20TJ+0nV2qqGqF2x1InwwQr98KC5+jeUWD9H/5FX7yjRUJNaUe+AlCKM8aCfAU3
xd1VMiup9YhR3v8iQcikPvvK/pXYIkoDQpjfvazKUuf4ClmypwYxBEm5DbB7m0CbnjIRdLIRRKYe
vhRQ5E6tb74NXsS5SeODuMbXaSiwg0bvqGkgx/9xgS1gCUZ0iGySLNXvTnE4V4CjKAk1nSHTRUSK
iEU/NZExsI2WNcupMGn86UxR/Yf0BC0s+4BRSDrH5uOi+24UrAy/F1JrhYAYLBU3z4Ms9xSfFR0K
jeU469aKRc9WnVW+fFTnOBIaVLB/4iLex1SWHTSXD85HDfd+4xIAp2p3SRhrhw1zpTaDoxP2mpaI
X9u7PPFPE2BcvWzB6PghP3iyI9en7wAPkHX204SAWaNaYQ7HBg8Y4uROdRCaIUY+LB13tMDyALsY
UTaxMJJogMdyRedIVmw2MX+lx9OawpowcIvrjtb/pvcdkp9fQzhjHNkl/W87GSX8oL0M+LOfvPHw
IIgh6sQt2sZCmL/G3k+dCPlc6s0tK6iaE+ppw0oIDFVE3u61m/LIAcUvM/nwmAYtlQlLgsOwbTtR
mZtZhaEWfb40EHEJN3EA6qtxIWexdZY3PH/OiLWFGGdzOIBNaAGbLm43O7Fehpu6xTfHWtxfAC5E
g1Bs/0wxGxyQxHOIkRfhCWMeNflorxQelUeMJ9pJHpJtOI/uHvX+oZHdfWCOlOnxrdia/IestiVD
d/G5TJSDjwf9QB/LoF7M0uqHTKdb9PS2qixgsQhIO4DcKJfeqd1OqycdNY2o4Xnt6eDE11eN0fCh
oHGhNMd0ExQ7gZdVakAESHKy0PRkciBjBCtSXe64cxGzIxwqZV1GijMccyBNy7upvB96kBUwOrpR
z0LoTz4dYwJmt0UA56IrDgNygieiSD9/5zG7ijsOdmpMqfejMxTyiwekbkjdPcvnwZw1vvmqVZMC
tMJiMF9TmyX3WpYzS+GncIXf/EziEnUj/2MExMQqtVETZwGK+HQSwkWPlsqBcNJEp6Hmv5G6jwD0
rqOdNuKSWMoYdxZtF48aaGfSJsVB+cXfLl7pDTOmIy2odDHzwkrjA+5QqMEpO4eB0FQVr+4GVjAZ
9RhUIkImOqtFZHyckLyfoQeJQJ+Boz93FOrKD9pn004S8ri82McyxvtxT7krd/UXv7Uakhenw4rz
eBAh6EgxhgwSGmccRBPE0GNmVtBPq04Z+7Qry6FjkKq7HSbwrQhqVwodLmdp8CUeikIAjKAWSoN0
0BQQGmuAoHrieZKDg4t1I4H7bjwWRpn6riXvWb6Q2hZVidgMQv50hAc537uDCBVCDbTOeolnNZbJ
Aydhmx0JlOMsMcp5Q3SLb+4C/KA4I/7Pfqzbwt4gILAQQn6/VX7lUSZyvBGnPw68oKNYEGAD/++J
xMP/8mxUC0+iSo2rawJAxpGgQdo5mWTsTS5TLf2XtqVvTEF7jz5t0qdscg0WiwurBUU0Fhc7UIt0
YH5ptEr6z/PhdiGbPkev825no7kiZWZV1WqCbKVL+bVzSARXMhaI+Un6sSlghKKedi0S/IA7tCIK
75E5pQE/gZMA6hB0T5eKvNYlhiHLvFoTn7msrCDKwGUMnayafTvUhyrZ0GlnvuiGrdx8GQTAwT2e
g8iiW7OOVQwDVxZ/vm+rpS1L7D5Ia/yeIt9cgITUyDhCo6YqlPDJBpVTlTzxg8E7BXqDrmjZM7z8
p6gHnyIZNjhlcm4DbeK4jaazepNasLfGHrjUQtRQE4KJQ+q0QxnwQCXb/sUjl1jBqTPp9J4NrKZq
wB8xkTOFGP/ubYm7juIUbxafyb6yb2PYUy/ULIhCGqJYmyZrtUbEJh2lvsetdiP/0ddeNoKrYuIT
et+OlEA8ol4wEwovGUzMk3D0D5HGqZJex3V2g1XlJe+iuWzcURPJTb6B+9CmBBTKAE6eJFTCVcR/
sL2TX6Hy/YmgjJqrBju9QITJaAMeAU4eINX8HuK04cP1+jS/C54mS/NOaJdGvXyh8Hgdi/KKTzMA
33xvQbXrEo9zJnQA2hZq0uQOM3LH3uUZeAp2YXQtQVniv6J+9vwvyYbIm39VnQc1UaBum0xDlE8A
jXWq7FMbuSEFnL2lqKpTYDbJAp1L18I+Dhkna11M+jb4YVB+HAASpeiEIA4kZ54YN4/vzV+w9Dc0
7y9h5V7OVQ664zhUoazXvQs90wp5E9dQzOTq3P9p4rSVvMyrundB2v8ZssmrrOZ8jG7Vq2s5MTIf
zJj7B+bmAQjCrJgGUbEy9g+10E89IQoNt1yao0l1fTvDtCgd8/9RbvXiSFJB9MT+kg4UL+f4wuKt
vZBxPj794iaTK/z+V72tXFuz8sWcEJ1w9+ukRe9NuQ2bv+RKY2OoKbmRJXaSrAIqwnGWovss9fDI
1mGGZLVK8A+1lzUgDH+K4mNuRWtIPiVhkSHqKf+qQ+6CUvjWae2CoJ8OJPBwuaDKV7IQuGdtuINe
L0mUnTksvMNHx0gu8IWRPfZJTE3NEHMUzXXMKo89bVHKgvdXBaPYsPshVgXDSJJkTmql5hF20FRC
PquZAayZm1ssxyNRk2pw7wnyAZjbRhrhXyInt9gSye31v7/aNmA0EpeQVLtnZvYVxLs2ndabWm48
NkfxrlrOZpkFDCPa/sS7Z6dsVsMvMWtpbZ1yNjdyOgfq93vP0hX8HNQbkEOl2BqZ8+I/qLpN1NCn
llHvmClL2AHLwCs6og1/0SXx6g5Fzq9wJfX7NoJUT2LA0p2sCslGWyglSgdjwhpYj8UZ0QfIsJdd
cJ/p6vDfcHQhva8bW8mJbC9CCTYoQmjOfhhD8w5OUYhNaFm5PQga0HtOKQuWlZQ8Wv/o+rx39b+C
ClKvf48pV5nFCsqz1dNuQkZoIivxTg+OqkKWOhgWi8GvwZRqSqX074CCmFmndJoa6MKFb93iXg7y
EYOhpQbpUdLb0ihyu+pXMK1Nywynm/Q8c47bsz2p0ZCL4PAjpG0k/ICOv2S6mpGkgZpn2ZzjZH+Y
yIgU/OvB2wFCJCcMqyCu1Fc+6Ios/1LywjGZMeGOEpsUipVS/P8wIgRoE3gfQ97bP6tslnR96Kqr
yL/9F2wZYKJSpiTUD903c4KcspxPDrx1GwgJhjJ+BDbhvQa53yHB6WL9crNHBPsCFKWZWoDo9kqR
L9W9OB9TQqRi0ansuHjUgo+qya8LQuULuYJWO5IaXhUWb4fkI/2dscjH0q6KxCwtigHUmJxEceZS
W7Fid0nl2i5UHsaGQz6++itqOfvGAauay45mobDbdjaEI8PAYEprJ2lSMBWKeIp+CUazmdFNma/V
lujcBN8asvI5MVNxLqxmiKvz3cJ31wRLoz0msbdgRbDK0adv+sLJHF/P7DzAnbAt8ftSdjhmevL4
HBsRsThU5c9t1RU9nJ1tbb4zksulaKwfTVGyLn9GnhxxYtE4WuPxQX30y1ZaTJvTaRbVyBScG0EC
QKou+CrUzAkjWjt+tkBj08cQyy1XinTVCYMHxvYJhN8EQxLcnEC9/h47OwGLGrmDyVGDA0hMPkuW
HR0/1h/F4NalMbHV9EAkmNKXp44IkZCFvyfQMa1f5ZaVct/OR5hL0GWAr5UTY3gvTiAANIeYcXSG
zbe6V9iCGqZhURxhdw/hj6F6pm7Hdo1XjiKoovd6JnIX1S+6/UxH88+7ZV9NyGr9ieVlkMLosoAa
ithTuVu1tfY0+0g3dCYXsd5LJm+NQV5OluivVBdin6K0z14d2SpuKchrqiC93H6bWVAa9LBlMmEu
O8ywDNQh+6ehQQQrDOz5Pbm9uMiZG0C7lzOvRkUSgZAlswyPmWc2vNjLv+Aqcu8XUfOy5kF4ITxn
hqoyyjNxZJu+0LviHEigbl5fEAWQWOSAOr6O2JoQhlHlpJjaIxNF0cIEzPv8qv6N5FOAgoF4lsMl
IiPHWC8EANa6Vp6G4B0a2z3WognrbqguJDcdejYZS3I564UlHh6zgogn56rT/jnfZK/LOcRzV5kY
dmqm3asVlXxuCuZpZ7iIkCPwWVlVkBznvemY294jtHe0wu2+tu1GUVUxGBmjNP51mEnWwjiADX+Y
slyBHlcA/OLVzDe+oP/ugoDqClWg/N/MHtLLrsYl7yfsUmvz22yNtiUsOgrZX7Mg9BcgsB08OjYI
3UXYbl93ddRVYTfLXSSyQEfq3w6K3UJsSuqaUKCgbDmnwDjFxWGf488OFJTbFM5n7cUS3cyByJqg
JpNx6B6N2qJKu+pOzSzZBElRkTtWqPYZ1A1E7I20akfCs4vXqLyd/2/huWkAU1e7icVRFB74zFR4
azGqVEIhAECPWvkxDYbLJ1Y9NVB+hAFQSK2ELG+W0DXc2LUIVBqlHMoUw6Em1czUr/uj1Lpezlw2
QfzFd39N+cGCepkLw/rsQStkFDb3iGHXpIN0FL9Q8xNFT5z7DT0iUZZJGZi9yCHupPlyevYd5H+W
x0K77LhPB86s1tYztSJZ9PtjwANSgSejZg611Z2rarF+pjOAYK4v8i0D2MvO4/ioSbEC4YlOLgK3
IdfBvsimOGo0oGJt5STkE5+zdTmpR266zhGLNqm+ZTDso4/IFtU6fH6jMrS3tzmwxe8hwAwzsD4K
liLhgsDtHfZnvMEkiwGTSUvc33fHDk1FZ2WxgnzWjCpxdkUaIBT1IcfiPsJyvheezKSRLPEYpRxs
L3qfbxtgzibM1FE/Pc2+D/64TpmNvnkxqvsKJTaD329Izlq9/2pqvOIOQoYT1ms9NSANXR7HlcDL
3KQDjWYHEynDYNnN5S3Ni9m8w5BMt5DRtDE9MkQkXP9tIxqFZI6hPaq5iukRjsimLpI5HnlzD7zn
eLbedHUtP82mKghTpxThodfagxAZinhwIjk9S7SurRfbMonAiH/yImpgy8qE1ruGBI8li6w0xq9n
HqcGYZMccnLk38bzxFfGxYB78x7McghXNmzynqHxfUo32IDubYvX3b13DjGsmZT4Efn5/KCPWor5
fRSc+KTmE0fH0LufXsZYrgNjCH4dQTlrCFvFxCE7YTFYHoZ4B6tEWAhnv24d3l4+KdU0Cqs9inmM
N0PiXSOD1vaMty4jb0ZRP4S57A+3jaR9zCBrKNPFhHktLCQ8+9Jm0PNeOt5IZTl5owz7kn+ctVM4
nqXn8KgGTJBIqBfiEPpMGsXtM2P+AZVJFvpXDXRIclZJ/HrOiW11wdSGn5kNF+o/DNA8z8g/ox+H
0ZQBp27SrVwox25xYDCSwn4lR1tZq5GvbOz7ngg3Xy1vdA5FaKZviZjKsmoCQTwlmT8K0xddb3Tf
rVjOvo+2h7lq/5fSG4d7lJcuDJQPF3O1362eByWdz0ElZ6ilf5p3dC6iUpZDyBUHAzaAcbTU+/CV
oLMSX8gVSPCGpCgPgj1d4rUU8ZdBuhleCakvC03LtMt1p6CNB+EhkeEd+RD/OJHKknOUkRaf2Nik
Jq1Ud/lA2jDFcKBKwu4YRvfInJ9GXGIDg7d56h3EQJW3Y4WOxTKPR1n2KwH6eOSjzNX3sSi5w2dT
CCankT7TBlAs6UExRyn2+s10pDOJJc+td3TyMv1QunumI/9Gsq53+2ITuBq4PWyHPNSEtom4H3Lm
HT6zDNyHYjndY5fTHHjN5pHYIThphgVAX31zEVhgwRU87wDq/CjjOnxGxKqurm/LrcJxzPXnbtte
ucgj4vkAxBj1JEV+mF6anAd2wZs51Sb4UKPGORLO3g0jYgw+BfeYt0e/SroURt7M21XeTY5ZRDaY
FDSbN2L0JI1jEpsOREzuiLAmcrXXqhgC4/GpygAlFMZVHji5Wltr3XsHdRst/OPP11bKISj48Skj
T/DlYxh8v3nAy/Wc5UWzraZlFV+ybGw2WGD+cImt8IcVSqlE+p4Lyy2+Iz9yycwF48ZFmldWWrqW
gEklSp4/wrWPKi6IHeWPxb8ICHQ1AksfCSaw8zwHI15XlqqiWSMeqLUR1jqoEgZkckI6mYdXw+28
5/6nb2X3pLYWdCjVszZZQAvGcILOapBY+CzutOH9dbVi4KFdN8j4gzoWpTbFPSquu3OYAbHe0ztA
CMB9b/Apinzu1q5wHNXqmKx5F4ztQFomRT08dmpq9YDc/8DvsWTRff68hfN2KYSGgPi2Exp/pz68
/8vOWLCf/mLUxZcihk4ddH35tycAT2StUROjIt/6yBbyjM46ayDEmsjeIRKVhBfOdi3uleYLH5Kr
7wrSbVjHCvwLzbuebfDL5TeiXjQsk3A0qobVKNQisMxzEparID48wsKj02ZGrW8/66Q3i8RFBU1/
i0pjENOkbuB7MbTYM6GlpfPorcU1GZa1RNdOX6Y2EOL86hu5ldGyj06oEnIK6nwV1AbZJnUJ+O1y
jjiEJO3z+yCmBiWvLcOlzcWb1foM2uf6UNd/v0fv38WRuaMBHRq1oP5lL4YT1FbULxt0SVtsmTcd
SauaoxCEdw41g2gmExRsNfBXT0QTFiYImExwy7mfMMc35sYGsF+lxOof0r8xsk4Chb0BMQtteDgq
B6q9NUAbsgz2xLRjIOcRigjFwrCm0klK+vU0+r5Cz3wfYEGtj8SW9M8u1gL/2nkWrWlOoPEwhmiQ
PidGpS+iP3UbyXgFa6W99i5lEhqY4iLYtuOZTz2BlHQj/L1rzuuaNueku+RbrP0nbyHG5lhbV4Pl
IV4fT7S/bGLNu/IL4cNpxdKpDlefZV9v3v+sGmaKVe5+KG4p32U+B5spTKb7MyQyRSBkwmNAhGOG
Azjf6Kz5RlBypCQJIG0+TjxIGOzCX/mlDZkc77k72PZKGKQfeZiyXsN3WcGFboYEnPmvZNuNFwGC
YCWXEv0W+VnnzXCTm/epRIzvsE5CC1GqpjM4HnL7ig0yDIIa+FwhXxyQm+7hbDersqtzwX0WZqhO
U+KnR84hkvKTjFthO0nGUSZzr6idnBmbVklH9/G/N8NS4jZ0BmFj5Z3VjPouCm85eCJpfN37Z2fm
dXf26yZ4VI4C4s11qSIsH/uUDDmo21fLfqhdBXBo6j7b5ykWS5FKlxJdHbeYZDujp8El9zlOY/Yq
mSR73DC9Gtoi89onHZWFm+WRU2gj9p/d6e9wrKW34npfyPEu+DOsRx1L/S2ugZL8w0xkJwuc7Ho/
VfuVzxJLqtz372Y/DAM6136L/wiFcv+H9lweE++2Sn7tRF4oNmOdOGaE132SBHDyOvcTNyX53QD5
XiHD84yStDnfkuwl4RIE4v9pezwx78CmzIEDMHW+czFMYO9IaOwKyd8jhgWFeA+dRWzjN7PUY+pZ
Oas72PZnZBXhMAyNzsZS1z5ZvlaW6C3zFPGEIeQS5XSwAaXzB17Fc9/iGqRGa4wTAmxtEnOc6+/8
PmaFQ8l6+oc6kUx5j5YuHjYBy2qDQq8HNeGt+PHyrMCrm6kW+DbXOkFpes+yhtCwymGHwO/eM5QS
SgwBBCZUjO3IeWrm3jLey7ScxBhCEndzG9ookjcbiB/FjnIMB4xGPsJdZc+ZVrPIkpcnKiXjRU2O
F6TtHBii+j/UPMRHQbwk1Vs3Btpn80RTNlEetiyCg5apyhYW7Ey3YA4iXuHlPNbjaUU2WHUsZQ+j
dzAxmeu4NT7J3+NMv1idN6Pt4xdEJQVrZtmZkCWjHSzEMKwsTThRwPPEBq/DHWBRfr8bJCbNCAzj
RdK3oTk5PUm28UzHzgqQ/XUbuc5w+oTNNK1Shx1/ci9hE9Lawg+oMOCez8GRHR+0exX+yy3oKWXH
/8XWDUWjs2PHWOO7kqn/ya1xj9xBC2Nhymd6srjJN80/8w1PagzFn9u/NKnX06MRIOBtCbTMX1Nt
x01SHKnSTlMb+MRNSkB9B2uGdcBaDxVM/3kbd7thlVxByVN04/v7TJiREyJGqT7wYzRK/bHG4YXf
Cqvk4r8wY1BEqggC+/CvdHQUs78Bhk44rvExTpQGWqWreCdKId0ucZNPRP567Sf+wNqXxgi4g06Q
HFNURm+R7OE6fzUsnIcd6qEq0v31RUOtnMT5Gdx+5CnI/2orhME1lOiZ16810pkwgE/ersUHcH6X
hM2eXus/P3djT1kXbZTtfhqAmIvZh2lDo0EBXk4Br0syrugIyiskI8s2DUh33DBJejR3Ktl3EQaG
EgdS9j57GWYnbTiBJvjwlXKmPnKibrey9anE4O6TB32whr/LTUq5cuNWHw0jDcsaWimBSKaANXQq
2MTlsu5bAWob97sW96v+dCSebI2tq4v5jbFrhCcCiycPBskxzeFhvchHTm1QmNT0w1RC2U8g0fwN
016jEORnMGfCgeaxabxp/UxQUpiiQg2uooVJmdJkH1Jp8QhvUzoaIy8wkOIHeaSoI1A7IeTgiZvo
dF4zlvwUxLnnbY/PdhRv5L8VXd/h5gBarrIthXB7hdgpcz5QpYgpI01w/VYn9/0+s6l5mCy1x/Hx
zsBN1gbBQw5GbMdDJ3yOQ+vJVfOgNdmSpRgnqAWWtVnpyPYTvZPI/z4Ji+yKpg1cPUzRQd4R1udS
V7PVkQ5M5dr1dSvXvnTwyEkb6KzrOaKp3y96H8cXqqBdRp1dqJfJVryyPtsrzPaXHjcqP46NC3jy
4BDWAPbojzi7UERVD5o8wBamQLa6dqOpUrhE0/H+OsD3t/o7fiDr72DKADYttmBhxXaJ+0A39aq/
E2JzpiqxRJz3DpYHihA9AOmuQXgv1lY1on7IEaEfJqtrT2/8cKCLJLk+qV2cANLhbzFWZenx9ave
TFTL7KAiZc3IHbqFSRP7HYjYHb0mA7UwoTpj8MRXnSgDy2LGUkRQRIH9N+5HB2+pN2k3UGuRjQrH
XV0Ia1ljzNaOY7vxdcj9OiwPP6/tI+ZCifiq/+Z+EJHPMgmlanbshfO3iBr9mYuc3PQZc7S3A+bn
d096f74b2LLD+t9uX7trFiXo8RURe2VLxqRLy6zuQzoafRWC/pZBBZn4THtExjRUesX6lcfJmW8q
Pd5GKQKg1OJVWciP9zO5uKzYwLT4bfjBpF5tPrS8uKyRaYzrZ/Jw4L6AlExXloF3hPNNev58hDGh
JL9bUlbj5dyjFrH2P/XNj3F7YSWOeRxhfc9woHk4V/jFlD4Mhtp/7870egKyz7aOZ7ra7Wzh3Tqz
ShHLfLfZoCN8cL9iLscQ0raRZExJQfw1f/hXXtkt1xerOAh3dcgp2BR8biEYqYZG9ExjLUVXX9ov
vMP6Q+uYz7LlFRB2G4ZL0SjQMjGUYuIBNqnYBvaYHsmTFVNp7dLSDYrj/FUGmNWzvDrNQpRnpQyC
yEHsvHOXrfwNzBBiFTN82zxA1/VTi9ZJoeVFpffGu5JbzmBkoC6odRZ1yIFDp7F7FwkBBp2JMzyk
+MApFYaECrYdbw5ZD96O7NbCAeb6XoaZYuOyHrJg/6rlbAfs/BurPRfNt4JLT0CqcPLqJcH4WIxP
WX/52Bw3wcJ+Hed4wtMX0mxsPzup+SzFOhYXOnYSCQ0+U/2FKpLlxQ1iy9k+JjwPDz+f4vg00HwW
VCh4/UZcKFSaa8Wg95PsccrqigRLP+GFeMnBjoh6tVoOD7O9vHkP8eZjThAjfd1nOXqNG1SHzlGz
2LW4TfhqFMJH7/NuQB1JqsTs8rYGAAgXQRvlu986ktfHPoLqqNPozZG1Iyn8bFA5V3VpKXSVOX/3
KjjIGGEmXB5yKS7lTmiFyEoJDL7pxmVuxk0W47Y7YiKERM9E59UlImiHl+GoBbobrW+8XywiobrV
UopyQ+46VrUmWUoI3DvktEPqIGGDxRrSww3JA23SiEfHqsYQxiFalobM2ogmP8Roklk/pkhLsFrL
LNoJp8htQYeUQKUqpZmmYaXMen5SiBAkcrFjG1jCEc7i+4Du3ei2zmw3dXORZpTBgTJHyBGsxCC6
qu9zx2MeUvPM8OMWAi45Vx6WuAx7RHqnaybmok0P4xhsOeEh2zHni5J2Y3lE/8p/skJeOXpXoocZ
29ur+Sk5Up0vmgsJFQGYlt75Kxl6bgirEYpoiz9hBxhfk4HLGSK+kCJwaupsFZ3SGXmFtTj+XrEq
5m7a99J+29tqCXJfPXf7/97QPGLYgOIbXWmJeyBaRCq1gWPG0UlhMJsDJvys3YQ5GLoLMVCuZ17A
6KySO9pbhM2p3VA/x2oLm0m7YuNfpstks6JJh2kDan3H2s+g0K42UaOip0qcyHvho7LvRhoYyBuD
V5EBGVhKfJIctIHrEknPs07qJ8qTz1XANy/DAe8FPb81lGEyRIH70Ls80OMg2v2csViq3N1VVjDf
2brbktDOaQp4e+b++Wy+OtkQDy3wjPMpR83EKqtYfZXoxuabCx6o+tw+2psD4ICEVFixVQU7Dv6T
PRrmqaeg3OuiR4FZBLks8PEDkfpjzJxMKZfl+AtxJjR1+x7oqPEOyHQPJ4hVUBGld6Y1swNR0Wes
qJHXR5JGNHyQfuIyc07+LM+cA3CuRELrwbXJzmEGdIyRuVQPH5hSdXOUWUjOyj1LSdS9XcCCANso
xExSMhwcnoJEaHMEGdd2kIrkQM8NYyYTiKooii4tSXAHZJrXv6yBzWE+wefvs66a78xgD6YVWtCk
hb22dbuzLxtYne+9yTZKfkPUOipBpCW4ENaQ5myF8dluTLdFHZMTaAnSVF71ZXE67JD+OcWNfCDD
5YSX6VBOk1p0HKfgtxmZCgEadXamjDt/0Ea7le+7qOgHEU9MiePu5DmmaOMixXT4jffXY+UhRy7f
6Wl+ZyU74MgTtz2ISv9b+WgBeE+WUvFGafjfgZBwzWKZqdiPnjdAhrHNGmwDEbI7udb2h5Scp1Cb
8Ffr1dTK+Y2L3McDQY0fVtwfbuY7oT3xPMOV/hy2+YlXTE9Tfegdm9RhNW1/HzCyrrsDxXNXMFaA
tyiOL4+EXFoZ04HCAtoyrfDI2PyLgisltbayjUCAQb564Rp3b+L12ZuAty2DLN7zhAF1Y+FiaQjQ
roeSRZACxkNGT4zhzX/EzT1YL+ZVlXmHSr1JA+jMZI6dahHt3do5SVOUdZfss7mA48uerRwyDvG9
PUTZWSOjMzm05ppbElq/Q4pxGyNDI9cqpssd3JxW37j1REsJwnykdya77TaGg0YdOP5Ydi26fO6r
SaBDDbmKAnWpt8aZtAKF/1Gbjk1WtXu9uSWeMoL0diY71wPAPdroC7mEDKSCN4JwsooPGnIvu2DL
cjZ59AViofo5pMIwEnjyPuXxaWCIAQ8CMTaM/H5apjhjtBXhFyrbYQGTILAYUW32+4ucl86M1Q6I
I2tAGGfJoNdLjhGob/SJ7G4+E219IO4JsReYjy4saPzWrvbUp1lMU94uck0TNr6FkOUN1IShnIXs
ycdRh02gNNB/vtDQQuICkPYFPsm6uiObsxyMj6C9gdxI19+l4rinN5ZjzLBEZCvubzkKS+Brrf12
diL1SiRB1TjxwIgP7HatTu2Va3A2DonOX7n+T1ei6pVN8rlE7chxR4E+Pa6ye4pciCaTVkGhGLZU
EVs99t2mHs3TB7m5MOSDICvX7SbYgXujWtaQX2jQ9Rvg0i7P3iEuL354qZjWFrR1kVwWID/iRocc
Vxa0OkxGLhjGlRz9b3a2uCZRJNQWMtBQrzjVm7u6k90HPTqj5Lpk0yk2zMKz0BOfDWkh2+cZZNa9
FPdnjC6WvL/YSsxCMzJ3w775Ymuj5+Rv95FYccpMPsoElByExxt2Vh2A2FtD2o+HyflKIfUxX6ke
8LCdTx7TjvwaGQjlGFaSJ8AES78UtvJfLhjA4VWZifarj/GVt5s2hjsKJ1M1a5hT/xn4SGZ6bEQS
bDdu5nkh1Jci2IFEliqAJI6DIj06GhZ/PsgixEstYb8vhPde3FKR5toutTivk8CIwnTsn9b3110Z
Vg5FO2AluXIRerc7EFQPfHnhuD+iSVa4DCCob4VdK08QG0IzJ+mwJjBLxCszPEHPsnKwV8nv3sBu
GrQWmgO2ubTptZ5RwfpRCd9lUxJ3vP0rO+BcTanulrdvsZTwosyU4aD/JPmZnKxoIkKNqswY3y//
SJbwo5UOMXfA3M4XfWnl90A5PprquL48aCv3jFPUi8J3xaTRMSJ7cLR3Qk6Yb1slYV5jjwlS91hN
ILiOZan6Yv0yIyYYgP4iXxy3fSi2EVlkFbw6ZI3r3++xqD+F0jRfCFxe29SYkrmlnqO6tfGt2E1Z
gjLzTX7nA6UgwZT+MuTGoyoTwVMQX17wbv3f6v8NsqkkbNz9/3bMFKj+GLl4wWWG73hhO1fb4GFP
a5QYT0Qp3THbu2osR9EaMpmWywuORZjBnPAGdzZOrPSRZTdtYbm7h2AETK4EmlEUH6AxdgsfQj51
xijFVkVrlRoKO40ZbOmZzNR1fO/SaBhXommt4H5k2BP9dIIvHrCzJrqmAhgKtN5DdEk9gPDyyG+9
cmlQXVRNTAwdE4fjOe2IF0hpk5qWMo2I+Nu487+DWzIuVdGqWo4EsUS3q1ezUMfuQ4CoiBw0ZP4z
6KwTu+UtOBDstexaY0uJHWEtLq/CpzeVF8UIhZgEJHT0Fw9VYh3c681MMppAMZPbGbsI/LNcWXuf
Qgax+ddDT9auyMxk2wptVkutTwTZ3RZtb6DDL1cm+4j0PwurFju0SWH8WrEMOUc4jpKpvATN3QXo
xS88Nx6ht1U9LsJFVr8OFZya0CByE5e3wo/cCZtFYeWoQCuZdiZvrxOOzFXpSSA1FonqStPk9OHM
vGNu2P/HGkA/ha3Q+SGO/8KXaPFDDBX0+y5L291GADkg40XXCWL515zKxUl4OB9ekvF/pPq/N0uF
8lW9OX1QoBySjce+MOvWc/GOwEe2D+T400SZWhpdIFUzm/d52wXN/bgIjQFne9IAyKChtppohmLT
WXlpLBdQQmxoy4h9U92XwtrprYwA7Wc7VqOPNsGbP4xjkvsK3GIcyab9MQYn88F1muNiqyEiRCK+
r4hbujHr4OGB34RbWXDvyah0Igk0uAqn4MqjkJ4eRnVLsv45G68Ps+I3yHkHvrsvCkCF+Xb9uKyL
IxdQ/d+iRESgIORGL98G081QJRl4roFHuvgOfy9+UtGhUWwp5Pu9QP4NhL13Tn0LHnsy1R4RKY87
i4dqyQj/NP40wbDes9/a93OqxWLx+AvBoyadSre2Nl+BYP/UgJYc5sy+laZB5EcSm6cAUcl4wEW9
xtYSqik+O1L4zfm3WPK2eAI2kLVh44HZtvH+cREcmxUN+wwRb1aaGgZgNZn4FRkxs6Gmgmb6m22C
LZ186Et0Az+KdtI4Ksw+WgZYly991xY3h0iLJ8tK7va7bOAjj/tsA5NnuI19fvuZFBn3kBV6sldo
S4I5XDP0NZbZoraE3cyqvCM50/XTlmc9+08d7QHRcB7AFtEmurbmpy+fAUvTjn7gDU081AwqL1Fs
Y2Ts9LmpR0+5VGNY/1nSVDlqnU4o4CKmOgVz1X5WOBlYqxH3W2HFnxqK5OGxzpmbIeQC/X8HRNR5
DYuq3/xGUHzAWXEXgbUrToC/g1rk7QAvb5bxLW0zkarFHfJO67xFcsWRD2/zJ/N1mvOf1edDKAVl
XBB/J49H7UrucI8Jc61KjY51vSpIM2nTG2N7+hVbbq2S8ggStyFT1GZ+8JSFEMb04bDD5AJtlYmh
cVY8BjsNHElahwCzNckLvYzf4YHNOH3Dw17baqUji3Rq+33i+THTF5colHYM9OGCtyD/c8a7lpEE
A+Hbyk2R6b3ZUsnfPDSMRswxRfP1ZpgdvzcoCA9Drwoy0e7pcOXi+69j9a9383QWlWdnEHwV1I+y
3cdpQXPpotO0+4Q08H7gQHHckTRs+BS15VSF9UwQ/llHrQroe1ioGJTqlBLnJtML7PJeBZlcRxJP
t4HHt8NX0Vs6/uj33A6eCIdExFm5xgtoJtQKHir+jxPBZ2m+fdhfGxGfRdLEn+pr2s8Y9IHo7hzo
NYj3Vji19hyrYPrzkYQSEWNEUs3PoU8CKXkQExEnUF7JbzjHV2PhVM88xuqun+f1SlLVa3TWjcaQ
BKF1n459I0jH58q5T+5ozjMRp0/U5/+91ghLva9fIZ2iZHQqDuSInNNrC1JhHpZl3O83RLH/UyDj
xfMPlZjAPlunAF9xh3ivup91IyNMmIxwu28rDJI7cGw4OKVq2WKtTSb4cWbDg9Pa8FPJHp4AP+ds
xqJ8gNP8JauFLRk7oVTRy3Sl+BFN3Lf5NTQiHRop4FgR6OoisFd+kHRfFA3FI0jmKjmConIhjtXY
2L3jrpVQmBMs+MIzmBd3MLp3GFAgvoCR0ZGJV6OuoG1vc+vYDCDWGJcciZqd9FbfUujxWeoyz2E3
/+4fqAfos4mN7UsF5ceX5Xi3dk3hI83XdeRSLUG4dmvPR/mnIw4JOrLFbu1pczbynzYBJFd3WQfo
YgtmAR5bczVB5cQS9/94mE0dkwU0qKxhllJBCqHve/rzL6Vdkn2zXNHDJ/V5Y8zoZxDDSRLLtWmd
5JfxOSJ9dhERPmauedWhtBo2UP3/vJPtBIFSA787TY+ZPd1TWM6db6p4QO7d5L+LaYiAK2cbDR3l
8FpSb4CtbdhIP4s7eHD4WywSW+pTCXA0tisoTtGU+KDFfXxhSG9VrbpLOV1KDEdH0cNM19Xhbyw4
zm8UiYTgHRqeXhpmlfozVkcY86w0sFkqBagbYK6DcOZZd84I7xvZ6jWNdcI324QOFIS2BAbjdY1d
gL2U8Nfja8O4heTNYaMr4crvnBOHoAfO5KLZKc6N14/3V0a7zFvXIYDZx/Bxfb2TKk8y9+VBdIg9
nR4y+t2yIqDyEORUbNqA22ozGP1Nty3WQNwgIs6j1yEmkO+NiGHNNnBqCqVLA0fT7Ck2Dk8tUvz+
CRX+v0n0KuciJLlaQU3NSTuKETAFi1Wjnd261gRZSh5eYpFEsnjXmp3mSXQN6l51jtfWo6pRwFCM
SrW6+EkDhJpZ9yTbFXhtx3XCdxRA72FCibNyCQQaWLd1VHnCoJjIvSbpxZ3Bx5y7Hcmih3OD4/vG
+vK4HZmecuZF4mHWGQxXwE4MPd/XGTreK74VHXDJzS/OJhk7jCRn4WqD5jk+0a693RbMqJPhGkrR
Ctz6188CYPzfk3xWcb2Bu+KWd2v16ZZeh9HVTeTGZNLQw+ypM6eVWHfQiH1O4qCMdoa+oE1ca09V
da8kAC6F5ErSut3In8WTkLlrNKBgy84YiqmbaTd1f0au/RZENNwvOpbh5dYb1TgudhvH6OzVJb2q
d5QWb2fUjoFNDjG5pPE65xHJQsdU1RS6xPSnK4qro3EWOuMo61Zj1JvBitkRKmGu3O/PhdV79nXX
UXE31EfmgliaNtYVjib8l8kP120Qppeb9B58+6FXXqJhPivf4R8ojp5M8y2j4Bw6YhwFOtNGiiNG
Rcm5Y3n+yNz/NSZQ2i2bGzM51bal7Fvrk1kwLy/BBGgdZ6cL96cnajKI3IuiZj9v51yMh/ANWrIL
d0JMbONz0fWyDeRxy5GwJPLQJpeEIIO0KKbh1RQhw80HH1EUCUX+4V2DwozgdrdC0LkYMdFLXVUn
WynPYBWo5SO8NmicxhondVd+z/+I8zbK9/E3k/XyiIoHs3k64tRs802NRTLgbodMoGzEUX1DDDPo
XgSUM0I4Cihii7B1kJpa3Gomg6qGo9TSDL3L4xFVB2XPjmFZ6VXWfX8V06gzCZroHw7lzKwu6q4/
y8obZPxHYTKkbn7MzSzFY6OK+spdWmi5tQ2LR/LCiyYGqGmsRNdRCK1hZohEJ0k8kHKFHMWOfQ93
TKTmPSsyu1clu8BRVV5Ymn7RKjYIKPBGhmgBOuri7xJh+lxvoHcx3jJTfoFlqkQB+7PZuI60Z333
tNhyDX9jLHzHJFMxuz57Q4VJxtTSfvygNGaOY56bezI6Zw2tdfII9SUxdvhIi7Sx/rH1m9sdi8mZ
Pn+pVVwxddsjXbm48xbmvQv3r0/Iv9yvjFL1uIsmSl1/rZtNclrVBoZGUoMDzMtFEm4qanMwaFgO
+sPYPLMBUjGEE24PV0fhH6UylvMEO8rJGOCsDPCk/b+5jSmbv6ApFZTIoS699v/c2Y/vfxkmwN/G
b9HcZaX59MSv289/fdRJJ1uNWfGRDxhrwd1K8w+I55Du6EDgiiCtEi7y7lvuRdHR71xT05gutJgo
pfQhWlQpJNva9kel3ewhxEkZl+QDjZLo3Cy/3d9Iqj40MHelpD+GSJGqGNXFbvWuxTcOHUw+aBoS
khho4/J0TeSsUlcqh/PrvZXNu5VDudS4Xx5KYYYd/DCBTuCqCSvTkrODwaluN/pzmDQIbdkYHE4T
YjbXszA26OKvbgxkhTrQqMDiGD11RnKLW1K/hwAToborF5Nrb6Fr2a9kOvtYToJH/rCwfqPesAct
OkgkoJW9jiRUCFmFIyf3PUoFTV0YHXai41vmXFTEMU5hh49ppXsX0jSfEgjCUA8J00nNQY0rkny9
gDjvXZig2WPP9dzGwwRdfOPAeEk1Xc1yxRsuiXtQOQwMpyWX4sv88QdRxkGCsmuHLDigU9Iy4C5e
mfp7yC8eZSrvGONr4y3ujJllqzs4zQ0Ga6b+nBu4xjDmy9UKOnmLaXb9E3tLdKtgKpY6SB9Lo65s
ebwmUIJYU+r6mEpYfsA4WT5durIRwGQFyryuaflDlSq2CABE8s0VLFI5iVDjL5QS7InRsOFfkteg
XvtwlYFRL7gzZDs65CIfKPFlJqmyj+lU83ijsZhojyhHNmIPL49UBwO0wUMA9lHov0JXb0+iLgGU
wYujLCLmXSoVggDzqbjsGE0iD9ePyouU56G0sfmTkyu/O/FOieFz+jp1h6B8Y962uVRqgk8lw3lj
pXYEYeBi78U6wIgelJp2Uv8q7agkzvXTl89hLCfKsXS3+aLfAp3/ba2xjKESXWfBLMhmBJTKVokA
4OxM5srizdvCd2ZYU0PdNKrfIHgPQXNJqttd+hLaagdcaacNXWVFNkX+3IQyPKyHMjevOcp9x6HS
vp83hJkzmOLG75BkWKk+aE3iyDHQkh7pJ/LWvtCgMzX9S0JbO2NOjWciu3SgSgtmPQG6tN+wWc97
fuhHzJRIqTSiXpbCaNXeF3h+rfRugIwsSPjLNFD3l0sNe9Zp+V5Z/lOFR/K0vDzHQrWhzd6wqKhu
SAADx2S4WEkYilc0KQUI9jH/jeR28biaUXW+jEEi98JfjH+bJBRK76nd5YA88MasJhSPSz8/Hyw0
yEqpQgsryolQ79X9OdS/v67wu0bDLjQx1Us9/WIxHR5GFKphsbxJaojJEMicj1al+AXGn0OHE9Ts
RtPAaUpDzldP/Sqk87F9Lss5Fcbj1S6qFUWaz2fCy7zVId7TPPq3kqx3g07igKqd+r45aPlgrIeF
Fp71je/QyIqdtlGyXLRBRtkecWSvecFHDyDzTi4zO8Zax0fTDbwkFxIvBwr3PzucDkCbcW4Nvlnf
zSeXaulxTEpnwTDbOLrZtTybrgZisWnUNVuBtXG3rXG+ve1tX3PCw/rp54Cr2uPH1MGSswmO5YC4
hbdFLWpZzqJzWpbuk7BUu4DbMK0ewYTIHKpjv0egz44Jvve/G+QJB7K3zbAH0kVdAq03iWor+CWZ
fmZHp69RNXBAc/mMkI/wZgcMkof3Syl2K7AD8hg4pYJa38dyCmd68f0vqy3wd4cNBMrdnmPFeBBM
sb7PcFDcB664Pvvvcgtl1MQJPxU7ltMNPLHjTo0c5AzqUsa7q3sZw/1I9TKEyrssRLlDAf7HJ5wu
OUFBajsSiR3uOLe54Ai/WkbMZJWrTHy5fefCfJPXxdlmG4phveVdnzUVziPv6j+fKnZtNzA0A0LY
bU4KTv17WkVZ9Hn2iF7/3thluyitlbSLlvzMGQsCzkPII7Vfng0jTIjh1D1aGkSICQyKkJeXl0hX
fHngp+BPgzQbqYHfoEmtfKRwpl9Ip0AesguVkzSCP6LjfAO4u8Q4KBwtZlXtjZqjdS07qIC7QAp+
ORciWpAVpJRBgaTVDPY6c2tpYCnsLQRMSL+0x+2qE8lmxD4uLdASaOtMp5zjRc1kS4FfW9IizQ8m
/ocrbp0hNEPttjogP7BgIJpJKElrm4KoUtLdEoq4/E5saLJ2EgfR00fRseV9woTh24DH2ZCTsvzI
wmV2gDRTU+Tl7+Pb44jG6CPUD4dLjOFD70K26FY0+ZtmrKyuSQBL4STBGXB9xIepNa124TslIA+S
fJ2ivbhFyP//Llrqd2fT2m4JLMKxTY7G6Emf6r3Q6YbbstlRg+4EoKim1yKjwyD03UJ5faqkxLYF
kQT/eUJELI0FSWAiodTDDWFTOuF4c+AnXDhmTfqRNllpM+i/G54NisvPxi685H2IA6YIHIk/Jf/9
G+yh85mJuX4PZ4Z9e2JmG5u66p+mYtbjjlxamRFOmoc+jW/BkHQEjm7aqiSAMA076RPRzyuqFSbb
ncMb7eN32Op5DAZVsW5Tal//APj2vODj+1WAmKgtxCikJF8nhMdoxfaYgIYCkMBMpxNQ4eNATYaZ
D0qzXpKN93SPLa7DpRljDeTHSI4Uy30bDB5T3lUpMVeHpUTS0FFB5VF+xB8QcZXavyZqszFgO5Mw
BUJD+Ch24WhogZRBLKlofd9IreuH9yyAH454I1ScYCGHwpSzamNt8uZC1u8hVLise5ekBJWMyVn6
FAn9YJcselPX7VQBK4Z+tHN+sGkpnoelRNmtEocR87e5PjDdKu3b1IQyfIZ0S4V+AulGME6Hzb8U
hhd7OpqU6BPGaSM5kA+qV9D7AZCdDamgZAJP3LPYD/OeV+zOsnpsg+JEJyLEXAwgmrSkUEs4nc7w
l00U7wx+kTgZos0D7QCS6jqd9ohmcPk2CN6NX9+ihwDhxfdTGDjLEKKsNvfFjnJ0wGW0QpWgM5kn
u2zLf0YgwpSzohenOk+BhkEmqzgc6y1q8X3kZDopplW4C7W3qCs0u30eD8RKMUxz+qipBnNOaEBc
tgqJJHubaiWoNEypkhKTTlB3Cch6bF19c324+J6JLmYxtn/tWo3XezspVu3WM3c5xwZusbj1T4sA
Na1HsVazD2FZaGjIxKJI0TReV7D9g98jXARc6XH2iU0jb+peVvflgW2WX61Bb/ZWm6cVZwRdk7/k
abplt2dP1YvIZZxrituAwHi/fX8X1Chp85KOR2Ov3jrnFpl0w9qaEwc7UsEo26OBHfvC2FxbZHw+
HclKQu18gDEky+9sDMjuuY6aUk3PgU3Tnq/7vOqemvMsmFll3x+65iyvHiWxKOlYo1+c6rDeMfea
6bvHL4+VgmMgfMzg+ms0HFAekWXPgcJihbiCGRvcZgCUGAE9Im2Skv/hVvCt5ff2UW+CaBew82w9
cKAyCd6Dpq9bS7wmTtxarRcGI/dzk/q5WH+i1Dh0N0DMppghbMrjJkONvLKIWHI+fF6S8/yDP7KQ
i2wwd9hROQ/zkHNHcqlqobDn5bttan8Ym9QEN0No8v9VfQYRDUvl/V1h3313gMZyxWNQyQ781REk
6NX9fEcueUzYc0t+IfpN3QNN1ucmoce6EIxM8yfluA0paD4mQ8N7Ew/VAYeTIv58zTeDMyy655Tt
HSyUPQBFwOwut1g5uEnsRjQee5c3FUFNGErXS5VUfQBfzb4eXLYq4xRDHK1NCi0FZQm4fsGOkzH1
8x0R3+BUm2h027Ou4fO8shVnetryMdHw1/R8IQWsmc02vzmtUCtukkltQZjX+l3VUelVhGLA53wZ
ldw1+z1dY+nAHy/EkA/Kk50nad/7NrHC8c+x6QFqs0nD42VsquKcKRzNPk64pi4CkhG26ouqxJMs
9Cdqv3isjuSoKy+nGYRiEm/vud5kAsLi6T20baxedxoHhfJYGVycybZ9WJLKHw/x3GxehfOjAlBY
8G0hnQ4oWXJ1l7C1f3IfYhSgh2n3htIq02FGpUL+gp1jSjSuFMG0IhzfaGC5aefbzKqtxcfnFoQQ
d/Qp97NmQ8WZAQTZtzMKpjU0b8DxP1vd4NqSZ7FdVS4wslkhgBNwhGsW/zEpknLe7topuYts+kH/
yK90r2mYwe56GqWiRefqw0SKuz9qcK4O/J04p/ypsOS7TMwys/gXmV3aidwIt6eEfdsJa67SSArw
NP45Uph9EF/F7LZxZiJeqMQGhrfoWqngjfIG7x7VEzpX9/FP9gxKU71nleJy8XzN4t0ibeo4klYG
11eXCrKvo1YY6aeyYYLi6mde8S9F23lceNPHXCx3B1O2y8D4fH8/kzHoXLx7Ph/HEXNtKg0nglCm
9SBKVYiJfXJTQtuVrDziBeIqgI9QO5rMyLiy96QvsiyGSz2CY5IDd3L8lsRplYwKNEtehQ/Nu2C8
QTIRnMKgYqSnkeXgEsqd7rAyIwSMyj1J4wEFE7sbYuLnBTjxw7gBGlfeFStU4ZHp13M8UZBA4N8G
JwGtkqJb0nJYIlOc0SotjTnyJYOZnOyizE9oXRJLO2vJimQPd+ju9OKLiFwZU1ygDZKziAz9OqAL
rrJ00oAmah/W8yiPN7gelQ5a3UQS9TEKNQ2UHSHIFaSsZgXKugksIkn6+F6UoppBEJmClhcG5Bm7
jpdjmUNnB8WFmBt80n5nF7rhrTI9X5/9zCAG+JR5z3RlMIA6YkaT1kx1ra6V0JLZPHXfF1GzheCp
EQHvWee6TINMWH995OGQduvt5ELsLhCiw1F7qC3eFn1GyQXwWi1k7KFDlLT313YJBIqXgjLgPcAY
5+0LDXIisgdgIFqV4lY3KPzanu0xPv21vJzRnG6bhwvEnveyDA1ZwGEmVJRlOEVfIsu+93L/MHJA
Ft9gFXIjGcTaBnKoasJsGDsb4/TmuuJnBikx1hg91yTIWdKSOiVQVAffRgHBSTNBHCY4ZBhwoWtx
JKREzkPcBuwfwpIZ39jEIFhF/Qik9mog64iQhKC/IoKJVoTaEeKk8lDupmFTEZps/qpwv+Piyp7F
yJYZCtyL85CwWC1m6MSCRgLYqcgTnyjCQk6Ll32cKrkphTrMGeXBM7zjLSC7kDV91yf4BlPkX08l
7ocz5fStEC/w4g0+VQe/hkbI21G4VmBy/9h7q3fjPpNpPE3Y+F79dy+oibSDNG0wAPYNm8tW4TuN
OE2AhW0ScFg7KRodwOhmNtCP/zhkPUqBO3Uxh6dJVgImaiAw8oP9x67hKASto6CShvayWJvJqXP0
EFhF2UMdVxzoHQfVg5PpzBdUh9msx3KJ8Itt3+dtPENkGVBNZsQhITUmA4cR6AwLsEwnggQJn9RN
1rfN9+CuL8TCoQr1chUn/16My5UfdQ96Phb44Qau16OiU9/esrE/TkALCCfyX4FZjPFzvGf3GHu3
rohmSM6LqrIOKYDaXdJ0kkR1PNoRnmVxO47Y5Q4SDvKbmTUiMbFVuEZFIG3ipbiQiMZEZ5jIcpX+
Rw5dcLKrtuh8mirTVYnCXp1dv13MwXAWBoboFXDUdUZ3nSKNAGY4cTd/6+9CzcWVAChS+Y2iYGFU
Z2xXz32qxNkc3mL6ZFRs4uT+VdRvUE13DBRkXkdEd4uxevlPI37lY/3e5+w5cmMoSumHiRNAgaYv
LcQWClKaVQwzLd9BDz2IuilOhC4yoQlfvE7O3b3UFljDL57vz4sMPKEm5QoUkT6un4rtc+iJ3jvH
aNwf8U9hPmTmFGB1oJZrsoWfRDcgIYZZR9qXbBi6i2VGvJJJ/O+6VHNE9pS4BuC1gGV1s6A0Vp3i
l9X2pN5/rx87wpsq5f4Mq00aw3pu1b3keaYQCfRi0DFP6qOzFYcFzYhJfzf/EYZClHC1lJ5usvto
gMxbA2mUJaZ+E3HEsNArdR2DDARSwEyPB4k3B4dUcoJDwFnTpDnv9PW8Oq2wENvmXmKlSAdoiRam
Ws3VMuO1jCoNeA8MxvofHA7PJ7hiwR5AqjXagyIcQ4AWMNZvD+2Z54tMMrviByB2yTpxZCLPhCqv
rZNN1LMSAdANpOKdX3ZCsF9ai3o4qtnBE8M49biAdvr+NSFp12WabOSy/bgUzRA0dSWc1kcSvDF9
MvXOx2LiR5I4nrHBAgKwv4ruzt+tMegNIieHsnwGt/WwrmHCLwHNZ40DSzAUSClcTSJ/oKw8ZoxQ
OCEbwfCdPfXDFxtM0KIU/ZdRhgkAEIOQFQkrOC5NjDGRTPS9aJ+TZGdi/XkOIVj40ZRbvfPOEh3c
ri+7LXaiN69oUfSTRMaN9WS2Bpp0Z2RZUnisSL1wst+EvkdbSQmMBGgzg7wiDNL+rXsondQjbbmu
2Mf6GYvDoVEeimfASgVBbPnGphk5M6U5jTZG9lvR/uB2QXMHgTU6sPZAALqB6ZNwhQ6R9gnVaUke
wghfl4xp0lVeDyqg01/cuT8jQh8b3PNVRkRNofmUlsxYYKMMEHE+r2uQ/20C9XvBo6H52P3rUx7p
ymfavM6l3tqvKhnozyaRjwRVZqbLCKKBajprZfUeQND6kTuoxroPP8LYHclumoSAsArlx0HRB+YF
yeC4vbjFqE5NJTdvo6RB10gehjcM1MI41T2/adhySaJkzzpLR/5l5puc09k+ho+yrMyf+/crGjd4
hpYDLcfF2/QljH1ZmSx9Qq43BILB8Dl8sxEIzqbHIcxlQJgFifkL+TNRVvcEAlfbQjNWuuArNuxJ
zQs9Vzn9Be8OWdxDk0eOihFbJoC4Pi5qV0VDNaDCOTWeD4sgkzbCXu+f6qK8cB+QTOZ6KWWb0r3R
g7tq4bWYCOhtQ6r7qcglfbfQOw+5qo+meAdZprIsBCAreOTLYF6PelJvDEUU6jOYRlEAnTjAy1k4
Cn6IyKHLroQypu1ZQDYojNG91lVUpSLp7oyYawEjD3z2Fr+HXcoxctwU7dIUBIULCvPZ79XhGCrF
FiBmLd8+lAUz4yjW3r4glsERjUOvjXTWziutl+kDlX2Y5zOmT0vleyz8fQOxHM4bVoB85miBVBoP
HotHoLe6GWJnd4dFNYvqaPEw4dkuZNFOyP8ZcdJivgcjVpvyB9H9yROSYLNyTtmi/zf0ILVEDLE4
Dgqi9+RgHzAhBnKB/4HoE5I/wO8fE4vtOlNgcep/WR/raZVALGvYrSNYU0S8H/td6/hosnRMWoz1
GWN5NuLeMURdTEDdy8/tz9rD8dOJAnLnZbsYBROkN6MNjG6p3qsbVGO3ZVk5z82T71KKL4seKPiD
Ld6qfwoIwGEh9mJYHxLgjPloo7iK3/1zV+O0Cw+Hfct54J0WzrFtwDjBxqV7sxTdv4TA2Gv4cMGi
3CVgvTnP4zE35GXrTWVtunuS1+g7Vi8cndvxJ/mG8gbdVOr9MnupRTHzFcy0nmnRneir1Xhihveq
U4Xhb33BV3mXLj7170UFhNAWkFjnjxaiQqRkUQM6NIiBnOUWHoV42jah3f9eW2qaTBmsJ0MV9S8J
sGEIJMPQH2Fz+qEYALwjaspw0mpmITiCQviSxyu78aAy3CqNHNLCstTjU167PrR3RtQ4wpm9eX0g
AVsyAzu5Q5vzM5Zi6as4nWZOyEg9QL9KqOfVs5ReM1boi0XE7PmOniCMjM0nsvjE/1/zOzbrLqx0
TPFmQ8D6JS1C/5Ltu/6/TwDPjKR7yDv1MpYKstcnOllenPX0cqYTbVZkr6L2QsrEkXNAXme2FR4u
tPNyU2UOEvDoB5ii6ovMQvwQl0jWGruiutGRVIrdG9S9nwHHqkBiWX2iPy5TNM310r+zhS/rn6zH
RQpy+CaL0igI0PTIcLR4y0mpnDSmoX4o9pwXlQcoSPYKqlDwQ3TMApv7CbVReSQl0MlmJRWgh9qd
7KqpdkaszpsMlvKBOw7yPFhIaONGMhuKtfnrhUyA9EgnYvmbnb84iurPAbW9sXZK2kBp/xMCBYvJ
LH1BPk29VkFK5jgj9aUddJr5BwOy1JGbhdiYFv3lRXei59DJu1A4BrBU7bQ1fuLdy8m7bjJkzs+d
W0Yt4Zh0Xgwqu2A193lBVm3zIZUAbkluZroqEy4UjNcnP8Unx3KnBbgGFX0eFXfC359Jx7GoT+WU
uz+ivdH0VlbtqtoE1OFply+4GjQCT3cJIRbAW0mTz9y7KMr9UmCHfAuCX9kEJSmfev9vRgN+iTYd
9ncYeAySmchdXXz/cFBIsbqs5sVLWqneZyoxnV9sBxhHM3ccBa7f745+/71t4ZJr6mEnFAMwH8Q3
wGzb9RCNpnAWMRoQR/OHg50BJ2a8uzBIe8s1hvMXdfC6dJ1qStFkZJasghrlqQpSRNuY9JKwVUvj
4lwtu5/a65IBI5uRxLgMfjAO0zh5rGZXbUec6h8R414uAlmNOSmHdir2reOzEkebvCThUMkN3zkJ
FGw58xck7tsNh5Arn58XCQVVIsCNPgkAmDRPsyv5IwfYmUXYcexOI1sGEDiUQwFBZ+WembrLU5Jl
buipemFgy7ALjnd9nZ4xx8/3Bl5/PaKuUCEKukSFHBDF1B2iC3bjzCut538MOAA8dkrIO2LfsKiN
hOuXs9rKWauz7TTSfY2o0QL7AQ8Xt2vN34ngcnLQZGFm5C69hnMYP5EV6bhJwlYihvcJJ7rNcxsr
AJetkkXqUqogD1a7O5XsTP9rswqcnLSNoHGE9c0x3LFOJld2drisLECoK06GBdK5Lx1zS8d8WtBf
S8ISfLKx307AromwAVRECYfW1CApqseoY8GFE+IvNfqQ16rwYPUoh9HJbuhdwkUyNmXvOpYSZJHC
ZIwbMw+I95YkjM6/M9r89gOY8QwKMVJPXuQbq0X/TiRLNU3dZDjAbaFt5qUkBfxTn85Y0AexzAZu
Cvo/NKCwiV4x2VnnhiP3voj8QAmwbDCvsCAy5E7e4r0JzjEHI9EiTCwXcJtqTLuDZKA1HDzmupQD
71WwAnpTFi4mbqX1w2jKKLqu2HPIRJC/9P8kjn0KuGEofX5YAa/DOd+lYSpIR5fECWXTBp33zdXZ
jtBxschAAg1HTaG2xMyxkhtcPA0D+QkiGOpM4iW6swbdR7K/Adp5cjVYHGnvRWLMP67DjQYXzf6U
GgGM0JyEw0PsAFRxZZEHbUm2kIPiICAUtkVyNeQyXRCcKjWki/WRsQvBHULM2Jo/7R9AihVAl66K
6AkddAjuiDs9iq19xFOy8JcaHm4J2sjgArR5Ni9FqMteLegmzA3C+nTfmG6oG9iflCgJnjJg/V6a
CK7yxRqLrEVDUBH77OpY/17ZkP2gxfrZhEyFVHjbBt8lNO8kGnjP6cILSBA0yMUTPFTP3B5AwtN7
UjN61ASo2ZZt2aKJ3GsXGf8GYJYS65zxc3KNuuN+dv4YkhZbK+FaAV0Rl7NfDh9OcNplErSy5JUb
NBGj1qCt4K5PRl7UZfHjP+v4lQHvlIWaEfL0qa2VX8j2Hw25pfT0HeRpl8oTWR0BWCmiwdfnxus3
AVXR4J8HrnnOQd3pnrYujVUDKpEAWjMgbWEz69ghO0yB68k20sQC+E7/E7o/JGf+4BOwRK5JsvLy
zc1GqINDKmmQlRWNjZFp/N7Rmxy+z3r/MKZyBpzftO4qKD1wGbsSLANGncarbQHGxVD4RgJe2Oj4
CxrCcwdpweXGQ7q9gcV13nmAuvQPniVB7yLfAV/TiKcvN3wEApBTKp7kt3JgysFOToLQgcpte26X
ZtwnhzOfLtMLs97KJk5WBgPZXCyQA2HhsIu03vpLu0K/NWQM3BaJar5XF+PehdLdddpmvSsAZD32
Lbm8R0Sxw6+UPEjJywXYdy19ir+AS4txyiyx0m9Vr21Pjov+kkSGCy+Us42tMFU9bJLlZzFj24xh
+TFefIVCLYXuhpvEp3o11cWMSbB8YFvzsMT2kDs3tti1IRWByCHRY4v6PUqkptafAeOBuRKmSsoR
EJkSZEwjbGfzDEYxQSjx+yA+rMODJEkd7CF8mGtZpnLBwjOwCPbVz0a3CeW8WLjCsBI+xcuqL/69
6cW1EW25mrOc/QGvivtLFnQ4BjZ/UHbkeyltEdTCKRwlwWFAR78xbm5DnbipJIXu6Ywgw057XKpi
HU6NsMjKCYjN6eAnRe9bo28IuDAIzP+V45VX4iZxhJjia7AcW8Mw8eMWx0Wsx2nCfL8M4vlCQfTO
NDshi3S2DFxtL5XuykJCwzjt2rDdFQLQs1I5ikLqDA0GVh+ebDRKLnEzF5Zbv/ltAd+JbZIauT41
shRXVx24C1NiO1/CBUkIQL7ONhSl2JNacDNElxDv0J0QY443HQt1MAMHXS32a9OTssc272fT3UTR
KRVtnNTwH5ECPhwdtefV1rCu2/QIuXj4jjXXkD7t6urcFVte2NCCfm9/3vyxK5fBVwHm2cRMOfs9
1LIT/D/RIGQ452OfjVWZ0Qs5tQctLCd0ZW2KqcFEzhIvUSRJZq0OzvA2ABEwlSu78rWqYIbYDfhl
+hOfuUyeoW0uSY2kvBk67mEkl/TkNjv76olLaEOFqIj9yOk4m/HShqCo6nkiuKl+yS4mMs8nrxBa
XDJAcclSaOruFpt3Eb5TjSP6tqO8Dk/oJME6QkqhkKZAmYCUS+iAOvtuPiYYWxTRdwK37eiHdpKp
1AtyeBk325un6i+2btpiFPhI6aG9x6+bL1sxgkR5MSX/xFV4rNUKZLt/axsAZ4fFBLCqhsl8cNQ/
oG/pl1FfH9BVqKKVVckyfFxNuI+TgVe7hMpP0VZx+wwjii3U2+hV9AqZk9ep3NIYSJ0nr5deCr0d
FKoYvACashQ+ZB3FtvF4nkVDkLGksdwT5Q75zt8folf7+AcPV+BR4L0h/uQ+KSK7m7JGpGwgipkn
YHH7g0xrreCmqgT+58j95nznSa6i+5KF8Mz62WvOOcufmYclDxnC1RT1g+sXaGFg/ZMr26XHnV3A
oSSNzzRY7GnKUf0WKaG0pXUNYMJlOCxb1gix/y/2PznuazWIeaqt22RmGvgElcCrOZq30SBzF0W4
psRgWmrbxi4hQ8WVYDJ30ge3G6O99QMBBnTr/7w4pX6+yweMf+ViO1KT50FtYLXqOCPU/L2Og5df
3NA1QVrZCJA9AiLyrtdART3kVbVEVBD33BaN7zgJAoFhIUDEKVLLV4/AIsd+svo0YV3PPFFUQOlb
u3WBtbFFrQrwOAMhMyKVgc40LVqrtRfKJwCoLbQ3AmBgXGvfHCYW5piA7izEoTwEg+2rARH+ycwm
01gYA8B1xzM83kyfSwfPlSnz34lowvK1DEnPNM7gwq+EdFsu9o/OfGrcXDP1ZTuLkKrCuZp4wJpr
bo44XpPUzeB1FofhFBM0W6qf1okdIHceZNt/3lm1t7Un9T1zHzYsTwdyAdGbUmQbsz4JGzQ+zLJG
4o2QVYFgJsGvgbls7lJLKC2dHMJ2nFjG98RYWiLn3XMpPsjbwvZKDTCfLZmKa87HmpYKymHfPlRX
9aTrruFbdCCeBvdfax0kid7/Lg7XjJDKke/4IxfcR05nudKSxjtjTClnE8OEMFtB8mkxCgMnzsUi
wJGiJ/RjdQJrsgMcEFoG47DI4qBMpQMdcOJDznMC9N7A3NncsvmQ6ssPkJH1pKC1LlEpRbnjM40c
k6lSrOhpaJVDeyxz/sYeye33mntPC8fz9YPd0s1qhsCQaWAbiYq3E/SVHfK7EkRFhqcjr/V2Ljpg
ykOBAAMh5KSF0XYFNHb0jYadyvVKLH/km/0fuP8Bz7lJF6+n9itRCMOgRPWYPra1YUzj8yTJKsA5
UX0oI5MYXZSiO9DNwjfFj12iR2QpGdK9g1EgZe9eG33K3MIs3XVkVwB0asgZuJdA96SzOVXbBu+4
5qVpntrwkdLAw2k+3yBIW4j9PECXjheorvi1xGtXJbYqLs+G9Wuo/WB5bAfnB2Efv+GoNr/Jpl6e
SLHXGiu08kZk0sbTLBUW+uRBCXioIOY+sXtSvk7TomiaHjelqCroZXedrNPfG3mdEKr0Rc/l41/R
2HNlrCbM1Yd98AqoBolsGuYc6Dme4zq4AnaZSUT/REM1NwI3yARdsYtDTguzhOFLCP0+2mDDosfV
7udXpSiedKMsv9l4mSvLU4+bXsFSugJxzovK0nXN3Em+/+tBGKNRkrymWhwimBsGxmsGHbSDzEqH
NZyoemUSHTJgxVpZwYJ4Pqsj68B083V+uRVV9uUdzAQLkC9w1xZ370lRmiZm3iWQw454f2wbAsG/
tTpWJy+S8Upyo/7AjHnfNZq1ZokXxLL9fmmuJOqF6/nK9/G+jTUatQotgN2rKIJTIW6eHNPrjqQT
LijO04Q3/odZom94SSBNRwUHpCPJvFvGd55Dkl4hDM4scO5anr3emuOa7bcZ4OPQUutvMtFfTbaD
K9p0XT6rCva9ZcTG0O6yTesZwSEqjUwXNB899QQBmoTKOZ5TX1G2fsAj4joVJPOVmNUbw1+G9o4O
vcmDc9HBijHtsl1ir5i/FbfS9ij7A/01lDK8yuJEHIS5t3jR//a4oraDnyf3cmOpqQsGbRxBoSPd
e0prveiXYfJskJnwzD8hr+Osz522fggjHiMWzgH+JFe0Conkyb/NYXGeGxeHnceC46VYsT9sIaEw
aCNEf4Rz4IMImxgW/ladpOV+bXmfsCxYW4ITFyWvd9wvrKiNVmAYuBSPKkj51TTxmSUaz/1+fEa9
7PgI6LgakGTCtGa/NaN4pVpxVieOOXJqZnFgMbCIfLTmcHKthw7NUdQFyqQyI7Qm35T+8tXhX4f2
6SqxQua00EIyxkC7Vyujq4H7NJ8bdOLGJYy3ySp8Tj72ohGH26JW/YPQt3laJQjKqbim8yWFMdJr
fg1Qi5L6p7Jm5v/ezYZpdOWquRYLy7UNGbJy5rhLV7zvF+JCehc9938Ux2lYcPDriWULkEtvERfs
j4kfPydPtTwYL1FE+G7XoXXVA+9TtAHhN5q+gn5ryU1yEkELv41lU6+wnxms9F1kl4aCH6QGvTMK
OvfU8Aw8Q4drRh/V76fc1Osub1Uww7cmH7nQRv7p/46Tdabxx6h394IIYDoWQ9TZ3fplEOznJ3a5
apkXWitWSkgPvgtHbVbUjphoFzidCHpG4eRegbl6O8A+lAKf83vKv9oLqVSxOX9RrMrrueOlc6ib
QHtyIjoDp79uvGJgCHolLYrk7oySjxcnbZJzpUyu2m1Ew9Xi0NCWcs2kGfqQSnBJZKxLoJVHRepq
Au2ekdU2fRfgS6crOdcdrDsjm3JsVi+sW1gbwFmzON1P5Y1ndt6T2dcf6wf2+JiJS+WCiIUsQeao
6+93Nz+bpQGgsojVnmCXJ9JyuTNOKeUiOC6o5H+yxyKLuFdQiWSLX5rj7AdxGAMp64w2dtJoJuVj
Kh00Hjc9zl+vMx6GooTdEuksFVOP5uKroVjzaa37cYuDZE87WWHhJkb6/9RJqVuTj5UpoqinrCuM
TYixwJzVZkzUW6tehCmd3ba78xfRI8mLc80NIJxOcoWKI0w/pPkkmNC+dOJMLVQJX/VALth117Qn
2RKN1ReoacszjA879Ea6tUJoIw8hm33dZ1yUZsg5himlS6X3V4GXc9Y6j9CxymFDpu+x0zWoo+D8
TeKiFQE89HYp1BY1lxI5x6VIRF/WJo6xpsm3QaSddKOldtO073r99uzGDNJjRmjbiIqi2Gdus9jI
UZc6WKonO8txBPUkF+E71w7gQe7YdfjCzmQ2ykg0ksmIZo6jTb6rCPLxGeOYzHCAid6Cxb9wPRZl
J/Zs7KnN8vQNBOfrNAoOPBH755RZ7WLKCPRqI7pHcwCiiZ1x0DgMv1NUt/OkisFe3taAGJx02EXJ
druy6fx4XxavGFFv4xLdV8gdZ9fzplBTsEfjAXosrJDRu5LlNmC/mn3VV2ytv9uTn5/vRUs6N7Bj
jO1DcKctUF0BTmMO7/tm4yB2fy55DcGDEB7kFBVfGRJRA39Eh9WEtoGSbdqx1OcAWOA4JDha/HeC
4ntqD8//ZCqd59SU/UhoQ+8TNpLkz/m9nL+vsjUdSMTGg4WKSiTydsyXmZfhx+FJ4qyXg92BpXW2
A5RVQz0cruAMu2IDdXnbWhHON5S+VLbTuQ0h4fBzdED/yiNYVvqwO+CzQMdb+5f87/SzxaHqHG6H
6cxj85gWTlMeAvCPq5R03JxwYR5nWjrLukE90wT8QmHRhUwKkfTAMyz32qN9tGhCl/hliUuTT9xB
JOZksF7+kosOaTtN8zgEuPMDAJ2inJJkENRTEes3b1MPZI/jLJUn8LpAtbjAZqqbU0ylq41vCfgu
JDOdWhV5JL/Z44gDpNqyGf33KFrfL4jW70t1lh5UcI57wxqGPBQ41zWgbvLSxblZXE6aknZ1Wd/E
Eb1ol6b7OVG3adu5zeUVhZpucn6JEUWHcZ/TcMs0NIp43sKIVVrtXujccTkwM8WBx7VqklOtfAy9
+EvXMfeIqjc1PiedsmqGrJiCaxagTX8TiQanSkz0bURUA0P2+Umu5Q0PjJWKrX4S8xS1Ch5a6978
2rKgFPyl1ilT6J5D6ic0kW0G7YvqFHha+atKnk31jLkryR6LR7bQNuyLpqdbGPPac/WkmwMP1D8s
h0WVFtwuwLClR7doYVYeuMNXTnP+jiU89g699wwK2Y/PHM9ihb7uAOOWBE+/fs5NrN3FwoucE9dC
NzxmW9LV2XnLB9ZA44/lSTgumbr0grsA+e3robobH0XjmL6G7oA8fi2MF0ca2NC8zcEx5MNRzH5E
mPx27SJKsErZHfsJjODcKHp41Y+EfGERfUXQoSXSCM+JkTcSV3NgYokdkxU+nxBJZyA1UUtE5Zar
CYUwZgGqPKETWOSjMzKVmLzKaFLSt2imkVPKA0KozSVe7RZJFNzYnFY/3wPTlT5/eZBDQ0xt1LgZ
EcQBSdbSP1RAvNHDb+qkHYEdNILJwYYl+TNKI71YmwjTRtpkrt3jFNGFXYLXPikBhfec7q9WwKtN
Ntxce1UtZA8GugZVqA7L6nvchoL0ylOSBBDC3OKRxm+WzrcSfSFE5RonNuArIYzJRlGhhXKOiqEE
Oqn2c1Ug61lbAKLZA7vLO4zFM/8vkVhZlOxgu5jYZClrEo1oOMunnTHmOnXOU9ILjYm08Fcu0o0+
zdh1TmY1EZDlTSymjEc4vXi62l4MgT3C9noql6ubO75YjivbtAE31tZry+IQGdcB6xC1vkphS2aH
t1LVSqucCOX08mR3NywlpRxawngUyajNnHckRRM2x7SyKs87iZNBvcriI9W9bUKKWoFnFuFBxita
FIKIX3pzMJI8GXyCZ2Zltprl2qwzoeCJuj3F/mPNCjfXVBrUvBpV7MITFnhTlgxgpNfNkiauaMq2
J2m/5hLEuh+FFpPPKeoD66aWey7cijYExkHpsVireMF5RzEIq8pBaCSyqkf5Cr7wWVfexdWSJnAQ
cjq4TTfiwgQFszhtbJ62gkFd4+TDpnWxjaytHvgB6VRDLh8OTfiZ3Il7ZX0dmQCf59YXBS4Ys40V
w+aSEVc4i0UrZL28GmPw7UCO3wgN4c7BAKFleQVyBo7JspHZhRKedlN8KPgt2AvDYAIOfey/jVWQ
4fnIyCe0wcEqfMpdMuSL0RJdsZuE2Y4qhQF/JceZBlMFW3oLh7qPiWuQt0iPA4QkFZZRCi4NggJK
KzGDDasrwbD84rIUVsupOHskGhAcQbaij0wYJiklK1R5isA/Br1evSFP05U0oUAAFaT8ZBDmxXj9
YH8vV1j5NjkObhI0FQeEDcJ8Ka772/Q/ZD00W4mH+4FpZWoGy6bW0Eimt9QvV18Dskj4ClcAya+1
tjTEk3Dc5eSwvFzQIqLtoEpdLX4PeYCjIrVHadUh8AMMGiICy1h/9GPxsV01nQIVmtH8/XchUpCD
s+6UPKrEGnAErZh+79dqPlFtLBJOE7UIDx0RyBC7l6SRdtNTD2CLVAnwKq7fdQ23MVGdhCuyyp4w
4BOjQNHyAjAPBV5wAQmg5M+Y77VYRaxvqAZ2h4fazd58wWyxM96U6kJNkAqpykwm6YrHnjTcLnRU
1at/1nwztN2td3SNSYABjMT8LwFSO0yvctzyIFEi3ycmLHvIQU1Zc9K/j9eISlDpwd5QTunUFkLu
eimaqRyi36ljhDyws+LCf/g1mPj/56s2MGdB+N+cyYtGH98ZESccSYp9eceRKB54ZUV6wirdHFR9
4DXKm/q7VtFy8n8QIIJTqTT3KPOH1TEtB1PQjF1fhaGLaSqjOoPZXlzBSjuT6WJ9cYdVKJjXs4TF
sFe9PpG2OE7DdIMRWD0GVN717NK/6kk/LELJ2GfD7rKuKCvIXT7GnvSxgeWxmQa8I94XXMJJTLYO
Q4e7z2/M4RjxqbITsDLfXJrEfOJJAKt3oA2qJYZr8Gj01vr5fsbzwHf3G3V01hGal724dGIzmzoF
L0MU+sM+M7bn0khYV9Xj5II6UjWkIwr8kiIpyL569VL7teiEDzTkpvUOEY0fHVyZ7PsK+nW2hrWq
ZAaBEZ0YCZH8tHn6aUmTtKMwNQA3qPVBt+mTrpvGwjjqJEoDOgvCniAalC2zHPJDx5BBAtFayOp+
+lgpryN++G4zOEb/cFHRktwXL5t5RAFDp3fzdy/NdgxRFacFWHZ8xR8L/8o7vFbTxt+6PAnNLWLC
bxhQfAuiF9iWT4t3oplYtjxm1+u/8y8t62o0oeYFtrsnRQWc7U2+uS4Ws7eQMaberYM5LZ+nUkqN
/w9yTu4DEba1oiCaV+MVD7AHT/suOH0cWvOkJkaKcDPlrceY2kt3J2BEJrVXtZB7VLkWfcyPEwG1
8fKQzHuCkSTokhdWUyCC4LbFjG47wotBk9bc4KOWImG6ipaobPUXJoeiyOk4vPY3Pb5Pyb6Jh6gz
YOfHvzdjfSzIPW87zW2z0uCc8aZkCjg/d2/KHvghLtpmnaijIsQT0cT60FC054PcPHzDgk5YwtEH
s3iCP0mL5LLLSpJOTQNe2gxvtOyqtB04L0fB5sqTDoGtRK986PU06yhRMsNX2gLUYoogfDwQ3LEq
hH7hf+Ec8VL8HOHGCO8jPJGUzaeG5pt7dEd0k2ImfwuOEJnzGl2V40TgPG0WiL/W6KKUKjdiJ8Pq
ZGFWJyjfUjNR/GxiFb9Wnxwbtda4KYJCLd5RC6KiexWCAelWXnS/sztVKYpZqARSib+P4HOLTHJG
OIiUlFxabLNSE7dO1baD7U2bf8U75KUmZF5b60HsduF+IcIN7UlM7/EkVNFr2LMN32tLaE8OvcOL
o+lR2muW0+VS46K0hTcjP+JYFpVQ5uQ5ftmuwaZGG2/MC0NOsdGzFjcIkJQpmkG6nEm3dDdrIh2m
9WloGD5D8joA0u+Q/1C/1tc7B8CYhDncOBlSP4NCoTrX3oNp0+UMvziIBfj24xqRXNlEz/UHC3Zx
6S5zmoxd63QEZS1zFnhVxRS+LznEQpQFzKqaHugZGlOrkHKzQXc/1oXnFCtyMABwiLKbu63Evcfh
xoEz2FGuCrgGE0BYEXFGpIRnCZG/bXloZs1nBREjgk8eyU4X18JybyOHucYe5OnmpzJUjpgMid3a
FVw1ls3vTRYYOBzsr/s2ZGIEl8y2m8r9f3K3loetfYIT20U122mCC8vn21FyUz8SXHwoDfGhIPD1
8cmcgP55Lfww9PaWEzLDj/jdbPD6/H4c1LLraTDvv/6AOR01jnx3h9nHu2vk8hFS0MohUKs74QGs
jpWKQZNb7zdt3Tjw/X3/BKS0UvBP/0HgOM6z58m8sfjDpYcXLYhGxVflO4TIirMl0Vl5fA8oZm6h
4R3jJcb2Zx1+wnPOdccM+qaXICh20kfoP3/Bvw/8AspHkDWMZjkxRS+qOE4aDptTrlhvvuhOLYJY
wF22W7QujNd5j1nC4SYDXIE0qF/vAUFkhcUHkBWTlvLTnpU8s6T92CKqo96VzqbXMZI/ML/r2Uee
G1n+HI8lagSe78t2dJRRSqLpN9YmkwsPK9hjZk6w8igcmqZyjZygPXEZvfdevH3hIZvNJBXwrRBr
+d631s7I21k8p0+wkUfcqmO8CFbIRm2OPmSnyTHmqxp2ZX526O2CUSF7GmesTsRRl3ssqxVgAgIw
c7JoFpJFNtJuUy9yhzu5FEJmbkiLeDpwn6vqSbai3pg/U2o9cpoy5tLGUnuJv4swkpjKvX4GAI8k
xbmqyiuoT0vzYazfzCALx6QMw8+jMlrCdoU1jJAcKRC80LQ8qGZP4+Twj+kRsk8f2gue/HZpmGVp
yaY1YP3cgvcdjVVgNOH5sUoeGKTkXR5ZqfN8J/z4iAYQGZ1S49c9J2j1L+6Jy6LoEOZtikqEOFW+
3NlBpuJv2vqTsa9Tnp61C2ypUsFCNSZER+RK2K6dhp+cPNemF8jXYN46C2QIYlGOLbykz0wzb8CY
m9inw+DfW9bIMoWI9PDeTcZzGTEEd3vbIKO8zjR71MUBwn0wjU6BHia1TtOu46uoVtu2cm61vvCw
HawmDofhS3avrLvnns+IxpfQeVzoJ0CMQnE5ysUHjQilDC9K7fiZmMhlTbzT3TRr99hyQ5vyieMX
hNL2KSBwYDb8IG7fs8aINosH6Tp//moxXY60c7mdNz4DvaSma6E8CWbc8IteUnDsXva8M1h/eT8h
YJRryY1+RuLTCflexRIfYcXAc43wsJf4kszXHgV2CL0Bsac+8NZ1FGUAtt/k2xmpAttLeDCR6FhZ
vRvxkAuecV1NycS0TixK6xiixJxfN6cOuH6enZefz4vnZ/6mN5i6qGTTVulrU+mODy2Zmpx+CvVZ
jPOQ2ZVjXyuOxrIgj2wiELm25VtptpOtOSv6xOomn1BsGZgihpJu0fUCbXQt/eLTjrcwQQQE2f2z
i7JA7K2obFIVVKWuZ7LFtaT7aTRaOpG+P4eOQ41xslpjDfnhI0832gYTDhY5rNaNYeJYe1aWTvBb
78HJ1eJjCiRVZhf6w5+fCXpuVXpMQd8IxPYpBkuBOQRUG0MTPEmAGmbfxDyB1mxIA53eQn+9Dbqh
5359z5D9elwoHB1eJ4GV9G+gr9kwVbwRjds3JyCcw6run7wiNLY/Xu59kRy59sbGEjFzAm/ZBWgS
1IAt2UQHxsfwJIhz/IQGmrMwd9/NXe6OKagQYbxg1WAIwPT+4gMhtLbqTx/LnAbow0GebGtKmswP
rum+CMmgLw+mf9GxAImxNdo2ioE9LW6b8N6lqFX6k6DHSIt8rsGBsRU83fKXNOMdvZ83ABZjnDd5
JEcx1hKnPq3KwDuYVYgqhsPRpyptlukAtF8/QaowWm0P74Wqy+WhuDj9xG5vEvjZS5xbdGy21ncq
zSn54TWvvleJJ8NVHbnLFGH+EjBeudVw6OrWKlMu47YfHruZLpaU3caFj9bChoA5TN64gYdZYEhA
vFKnATaz2tDu5n+fSqyZiTapCixCbyeIN6pmqiOiXaoxYjtgvXPPB8AFhMAjPYT8E4QgCq5MdMI0
Vs11qWQPOpi/ZaVJGNEo1D4hTGgTUcRGCMORODiEmoV4AkaHdLHdVRD4f3Ui7RiQA32kuSIACtzQ
p20B6ArQ5sMADiWPQdKmcxXlcAgaURT7EWGtXl1UZsuo0jN/Kg32KvZqf43Gomb3Uz1r7B7R1Llz
yJVvJ/MhbX4kGNc+eJ1XLO/aacueKSyGTIkBPLbHkSLu9GOLRq20c78sMktEqxH+ijzw7moXDMwZ
t7TkpoCHhnjmNq5feGWDX6KuFriNjKQTMQUzCVut7eJcqfqO27aSS/sg2Adyal8hg4ZXQwFkYMiu
P+dnnBLsrcRnQUt08c5YtUP0pynRnhIS8uMS97c03wq4YpMfpdqB2gfyuxvBdUT9OSrsBHkIcKpm
VWq2/szEMvF/7xYtWnSERfZOCKPT5BS3hsuadYQKVCzWmuUKfvW7JnMaBgcJ/ANgAsUlwZXpIHWL
4RgpVVal98ZqvPKlvPN8MzsACKbFOiMcDUEhPMj5B1TH/tPlPNCnD4zye0bhwVuS+F5j6JNGVNwN
HP+F0w9X5R/maKmpxsBSKHhNYpAa+otYY4hB7r9wyMeLKlO+Xh11DxHtL8j6fP2wTRlcSEPzHT3n
ii0q3/xamBuUYWJkGxWHnfSVL42Uohbvxf0dN4lTN2MaWikc3OvcKdQTwsozqu0Ht6Bk6Thdlfqg
jddWmFHmpLYvs7FJcs3IQ/yRaOUGLIZ3+X5D+fU8BNAH7nQfkr5kB3PmBhIG3SDidoWD0dIRroq7
ebzm4wkJK6WFlkvNuR/ViCarBqELC92PqsWL89b1gCpZ/ayGMjJ0eQVC751a/arYwRVw/+k5oF2e
mi86Vdz5R5y4DespQ7PXpj/nLv0bdYGeHwB9WxBhRYcrkWOMbjjZJDSqUoyaODdMzt+1eA0p1tdh
AcRihDSXROg6nL+VjgI/RdWbiVPFRIbeFARC0NcFGyjsGcLT8mmr15yDH2ZtUzcPgWrfUBFszXXe
xru9F3ItGXLZvYj2LDTFsP16ZLUDKqojvcEDzI8YQ19jVmdH+wfWgPIKM4GaWeRJLY5UKjN8sYYv
5HyQLGp8gd/KWunPfco7OGG8mdMPVPFPhDtetI66fWF7vjMHqGUWorqMOsacSvxK9pj0Ue9DoDtH
33JcVqApJJOXEc7aTGVLLN8ba5CwC1YvHP3fgDIenO696SF40NJJlHA1nTU/RmLLyzYtMk5nTys3
pbdbO+/LmLMyR9nW2JZefLJ6mfXM/HcRGov64chlI8cF1dvbf00XDyape8Mbn1Bk6e1ZTAx4uHlq
YAMz7ZPsLy6wRJYVbp+MN0m/Z/XhOmZOiUHW4IeSXlbtrbZnKgxkhIPp7yjudZok648PvMvVrJt8
ySFH5bDRhxAH0VQCcKYxVQclwUu6vB8RWNVx2Zg+YBhQuVH+1WaTSRprGulOHRCIYziNLHtYwfRI
78NYTkNST5DtdnV8/gTQ+NExFtFafr6K1TJ1p+lPVlk7Qzqv+lPHnwRKt/qA28/iulCt1A5ozJjz
WG8gkntasltcf9EZhuVE9C7027fbZgnGdW9pWVkr6niUihRfbWn4gK17eYTfzbZGbBXDESoRKj98
h4+CJkSx3apqPN8OqWn8SCMz3h068UXA7in7h+sTbwCfSDl4qSmIyvtXvuqO6ULI1Bv6obadjTNw
1dL68EIPtju1SV9QpzjuFwlKAJmYR1CN8To/XpvnneHQ0+UIclOOPTIlg/KPI8vWT65gKcHcHIHw
3bNqcimFS14QW8onEslHqsaQu/Uul3eJl42d/6bbzXSchAwPJjK6LekaRZxaeMzTBnmYdoBCMNY9
o/fZ4DyfNzxIa8rG5mPibO97RI+B3uugS76W8FKNMMB/I2dg0EjioPmtpXXyWcyaVL7ZF62R4BwA
haWcmcwY3VxQUWVPGGJ3aOoY4V0r27yjYuSPuOSnmX+RFdG/K5JU6uESuuZ7Yl+DhHmOvczrWtgi
UIZ+7o2b/WUsTZpOgsZY9iyOH9i7iROoZQWD+U/6ugMrtN7MWbst/hc6QDttTnTUUK9o+B7kaDr+
VQVGHmNi4id8P6lU8kAev8qWQ/V2h0Z+0XHBbkGR2Sd4wQO7To2gaVFPGgjSEjldjJlM19mtbX8H
3Q67lgC1gNW5B7ey0KuA+dG3hSs70jh8NxSs1XBYr1CANOPr5rvcdmITaQNOcum3gJPS85pX+GCE
ph4ciKPPSQoOnPgojmX+79gLKGgH2s9iGFtCbdAykbdB/lOEeSqe+m2VZUnkYDRuR3kzI/rkM05i
hm1w9gGO8ZpCR9feaAHetdnRZGfA8kkb2fdfiuxQe6sEhWo1WuNxDkqgympTMcvfLy3uXW1avp9/
ZKD2Wd6fWPkXKF8IWi3NX/QZZoc4nB1cj4ps8vU0aOKFJIav7AzXLtvZKYbrx5HQ+taSv4BRMvYc
6eSmHcZogJlJDHXCYwKfRMdBchI+DM8LbyNj9UqmEMMlBSy5Ilg0IEzvLHc+jCjh0OnYDLcInFnD
+g/9YVyQ0OnSf8WOqDF5+isSl3testXGNs302/164JmeJZR6i4Meel1x7p6fA9/rorZAp4MgDKmS
qhKubxulrEGCwBAgBPzeP3QxhADz/J2aY4ieGH9vb/bWNxXpNl1kag22aBiE5PTuc9SMuHLDvwXE
wa4tuwc9AZHQiy/0q2Ck8RnA9cOso+t2cfWzM5Q1h0YdXBjeFxJdtSA/CpxzOukCSFrbKVYWrqeJ
Vy0xVmgChnEIs/4UFFIVwF3y34cNHLC/fW1DrZVJarywweyP2azMAeZuCcV7dn9mTYrddujZduet
veChpODpKaZuaFde7DCrTZJUzTnyciTmAvkR4OkB0BbDpiOXCsCaQjOmx9PGzDRerh+VAFJEObCd
s9+JUT2Q6XR33GWZkTnYDiDDM1Pqzl9FNd4glsB2vcAd+oQ6xjD6kx7to1aUHd1bm7309DLzKpRb
LXavkk+KRM/ldnsIHQK/Z2ijeVtKKmwg5GmqBIp5DC/tjqcfdNl/xPXtClHxUbNUClMIIaOevOEr
gBt1kXjJ/dQyv/h5TqBWr55sZItwCUIpXhe9Qx9sSLJ5O85VrwzCiHbuo1KFb2BOQfQtorOWQtQC
OUWZwhhG5RUzuYSqE3LuYs7fNL4ojPl2j3q2+1L4mTmnqT8qTvACtvUb5FTG8J/HJdKIpOuezlsI
jjulL1basCkkMauLPK1UZ8KHKw3oRyf86S4AH5UOeYdEyOuJIrSxMqGWsuJCvc6d2pTQnj7hai8z
XD/c+pL+hth0GQl0EMQ8fBYcDmiUU3d1m5qggyMysckNjwMro4fOT69CJyP2D0RrCFkrVA3qL0Cd
mNlI8SECAPhcVi8VdX+qHmsCEXX3JrkVv+L1u9J/IzaEAPTHIFCy/pAWcJN3EsfeuKuMwQKt/M+K
AO2pqLoaTTq8TWcccJogHI6ePfW+mXGbR029MJ2o/8q88qS8T/OMo9g+KDWThF1IaPwORKvRZpRo
HpWez0rsZ7o7BHF6saXc89lYUnEJNrVSXwO4T6Wuq3iDgbkacRL6KcIGWmR9vwOy+gRaGm6MVWTQ
j27SVrDjs5yCDy2uJPZhhq6SEymFV9opIngjBNIoRMg0sBdIV6GV10/nRhBDmrDMlSAHugNSul6v
xRUaPkQkCHnrEFz18r6D9cMq5IMss+euPXnMUpcHEgVpCd5h2pCQ1lvM8DYEZhded6VnnIFTX6r1
VPBAiy9Bhhy5XlAAIq4oCng4QhPzXipopAiO+qklsfg/9iCi/AFsEsNoYr7rCYqCQzp9oqip6rB2
6qCrWcyFsolAqU3ZsAXr2EbN6cwHdtYeYGYyUB9WQRk6NbLnqmzjg+nMT1Gd2cpt1VAKxVIl2jzu
uYJpF04ToKlRLvzibWV2psYlJoIC8RyOBF9TL4dLdHFA6zxFHD887gM+X8PkJEgG1S6YmqCo9djp
TDOexKUYcoGA7e+6y94eO+2pfLrQ/zV8fbMyAdqoxH+CaijW4kNeL4pjAWQzn6EXfauqb9lkeEsd
nsKXzmTjOdkquLGSDVKbs7ffbMUvoZphnIn3MuMGaHVVF795Ed7wiEi6MQLlwaEsxZ8OaSQxpg4b
hbUl/SNW7lktwsjh3hpqXpFQqJSQ6aRNJsDUqey+ESTK8RTjhOQ/UaOe9c2+KwOSq8E+Lx7Fk0Rh
XbCeRHDelkYIMCcLoGsD7fVVhsFBKeUYXgvu/Gg3I5C06Azeqc3X+2Pbd69sGBrqqXVxKtDFBbDc
ZNZPcor6OtfRSVYIskzK8LsOS8nMG6DaLlmmkcd3kg8QWGD+dD+G66CQFh2hnTleXHaHVu2O5Cf7
2uVQ77u/fAYFIg/GxbQN0Wv4EjmDc88q/Ml3yjq26x3AYd3Z2lh/yw3LMTsQatRnhqhOcMObrydC
1rYxP4LakHe9Co8gNdE29ml29o/MNZx0Nvw2+/HazWcDCOBG/DMJvJQeS1/RkFptj/ifQlkx2RKW
TKsK8B+mk8H/3nisgcY24u4XomKnISSSnx+F3vSeRz0TEXy5by7tSRGNhzG+WeEIoutRcsA5nSC2
o8RUTCkP21FGm0t6PvZZO3VgCNYd3Ed49l4wkNyJCMccAAkZ+wSW0GaMA+xYr8rLBwOks/+O2K/2
BZdbzqfBtkyfYIAGNWb6LNKwv/1FplVbSnck1gz42coWzteIUkQLF6hsto+ZCVcRNnkycRJ5l6Yj
91FXIFRFo91HAixOsfduq3BaK2cd/a1HIyLh3GcwSIPjEHM5Dg9XvDGD9XsDpy55CsPFql3PnfvI
jbxPJ07t5m0Q9hV9Ffz1RMMDkMx4+W9ZWSY7DsxpB+Ys+1G7iKraHJuwEPWZnq6Q6N1X15065g3A
XuZ7/Sr7Pl897AWc5Qi/FA46xrIMBvIcaANBgiZnb5XFanPXTCWNrhSUifta2rMMiti8Q7Cub0q+
tQizyzYkdxkK+Zef0hQhYtJ/p9lZ7PHOTLYvKRjk0YEC8SQJ/8Z3tDBUapZ7g9tv02dF+Mu2OAr0
tSPtnbkpsqBs/Vpp8mu/JeEYxF1EuAQtV9yUmulI6gezFOl8ntURoO7aNalWeJ9LTbmx/rOVmMlh
8x9G6ZKPwegF/VEXcWKMEKAnemvrMnn2TqFFXBqM3GQNIIqfzGnnujjtm78U1kbjvFKLWFwbsM+T
q5St2zVsu/3jr/y7RlpmpJ+iXLmQ8xWQKa7Crvmlm/Thsc1WEit7zZMUIuC8pORwDXYfod4A93EZ
8MM7a8fK6vwE4s/NF9iY592R/cUMndbm3kbsFzkyoUKwnUUs4C6XEMbEo+TmJwOHBx8dOxyEEJCJ
1y5cd8U7DE1o0Yrwr/02Gbbi3qux1jCz3E9BtR8s44lBQWPpiWWKdnKm8fxOj8kl0VN0OoITz63g
zZm36kIQtVPsA8eAuXijvdZqgLzZ1PYn+7N+8/7fMdsxNSvX+P9KOBxrYgsqjz/oOBg+SDEliy2+
5F2IHxLCT/9LBESIMFvv6GdoOn6d82EfwtWtGNlGuPaWZ0hmk1P2qN4MgvgwrBX3kG8Y6qIgBPXS
kHJJpOYg+wE+i8rnthPflJhFuS21oqmbd8HOQddVorAmEBV5pKjYBGGJxybORI1OkIctWO9EQbO/
6phhbcQgQe3isbcBFVr6rWUhUIE8NBRBPjTTnNWjgvBPlCVrFheKnqCrBkeRmyGLZOpj/XT7XC9/
og3EBmEOApAFzfbn9glQqdoA0KEVBdTqcBNi8hO3C3vj5VOsBP9d84Urwne+arxShI5oov68BrLY
LRkpFiQiIts5tX3ETj6AEYDwaujuiBpTw6tApWM7thRg4d8K8N5xrdJEQY+IZSyhk8bPuehWO7a7
Rb5CW0hlLSVMWX4ym2fqdGMjrBvuqp9dQxbO7gXwMTsPtCjwCCQhieNBa2NyncXSRMqApsnEkErf
+U1wrWj3qZl+boGBv7LO/kL15DmUIJe8waAm4MKw/DqO0NrLpXOkC+yFqn2SlyEIFZWKVg3HAbzv
yWRyNtgFSW7laDW0puVHDrjGqE+OiIIWOA7S0rhfzqt6+fVwMm53IgatKJdLJ3U4+xm6HsDam8Ug
uuiORQXX8NHA8lxdB04NlUCSIq5hAq0AvJpuFVlhMRkwTBgT1S6jsxvRCKplXsMIgddXg6+oXwKs
6O8l0Uea0UxqgfXwMC1papXIQ+xX+IH/HuNj/hrRd/ijonqV6aeJhnoFZvEs0E+5OtQfZ+ACVrP+
FYETszuYgbXO2tnpqImzPKoB1AfZw1fazuf5dXiWuZutgkOFGMC58TYSzfT/wnElcZOn1nWYRhjv
xMEX4AA8J1fSjg1Ncc/810CJT3DYLUpSZbcKkJuQSjDXSd5RoN4X59+R5J7PBIq1oFmA8UlJRLjC
nLyp27uQimWtpIuKOQrS7MCkATAhepjQ3DUhLKa3xi/NGBYlrR5DQvQID0eRCd6X+Bry1Y1RLotX
kwIhoXWybT5XyKByY5gBjtQmiJQFGecHBa2lGVhkFBDCNSdS2kfepq1wrHTJNcM+DlaNf6+I8tNN
Wl52ugiqVoFHS5NWIYrlF2rokQEFkGKCwAOPn18Hpb7I3Im5us4xDnA6iRymcHTVx0Lngwn1xqwn
OhwpY+Vfeo37TjylfOhjblo+VqCb7vS/VZVVCcYsD6mmmlRT4bTXkwk3dJaZfwjeIF0COPYzQpTg
TOrqlakoMqANFxaua3hyAAZxhUngtiV4niFkhf580lQ50gF8IUoqfptDG2lEBBgdz5NyyxKaVVKe
qSTTzOU4hC54/gq/vz925d0DuXnMjnpc97hXED3o8pTIffo1AkjA9xDMoHbxA/Ouj+jVJdDkxn6s
I30nDJfgcjrCvWQB0arUWGC2Jh+gzTIBgJy1RKbRV5L5y48KRJLezmSckIH8YTd56Y1wm+1KqGU8
Vw6EfyQcKmmuIilHYhFGk5IkC/V6LQVAuZN0rao82mjuYsmIuZQ7q3Ixr9YpSOT7KaX2TzbqqAsG
mmDxA0OHpVUQjyRfheq7CXrAklzdbwUUTRx846BOfvCzWpN3saeoceON/cbHeV8OfS2D+/SGZ5+T
AF2JCFe/eqrAWrtEZDWMr/0ULvyo3oAwCPhEpT+zbgY3nv/sHW442+nXs6gcMiRIRLmUgff3MWfE
DTfApp3dAzU1WTe9KBRmjVA6fTH5gs9wDeEq72iAUZGH5GyM3H3oYNg3AjGoAhZnLC5rEmux6ZZz
Cm+xkvQ/q0ktiLHMmMTn1oTyxNfVUR76XmeLRucTiQq1M+TJLf3BWuuZWqY3wWp1rvBz5Gja9u8v
a5KEAGKK4/dr7lzLLOgK0dnKu+pK/Z2F/kWuyTfPsXPLclCOGFmuO7QIE8KkARfjnE6xk1lAJjQ6
wLeIlNXiMnp6YW+IcynNROn2PHplClvSWnzP7PmG0yPSbLoXvdXD4kBuzb8r7R4/brQnF82gnbxW
Oa1zHC9k5kRcqbwafx8xLfhm55LJXhB0tWKJmCz0cOhe7q9R0ltBrLqKbrnIXeIWOBIeCB4DkwC7
mveOK+C68/jKZQfzmP3zTxQimFk7ONczhYjoihq9lKJ1N3gSeKn5T55U5s5kEEdngRNWsXJwpXgD
Z4+fQaJQVrj/nhnG7x0lKSTceX9Esb+qnOqcFRmHIPU5N10MLhQ4QcahTxHDrILJzjIyfQ/B+zbS
ELwrVIvYDZgIPi+Dzd5l7bKKc5F8FqANKxFCd4oK2nO8uNuATr8JwSFG3h1dTvpf5Fl62n99UDbY
F2p6Amwv+W+K026OpscZyF9CSTYY8u2MZ6uubaIcFGhD7lvKgdBzBsQbal+gUEO2tRpEa1h2Y+4y
wt1o6/ylWK+rG8YjbdA0qMfHTvqrR71f0gj43mwszsREzedWN71dJehwD2RKv6BAM1toM4HIJayO
waTQ2jBaM51x2tbblSl8h2RJ94CDKFTu8QqSyJADNh/dHUcdH8npMlJkv++Gc76qGIHylhfZ9I3R
7FcQEgTGr385xg/3RNygImXHo2XR62gJptON73Z2zxFECZRjhX8IvxpZc6GD0L0sMdxWITOOdYNB
apw2YyMUwXXXovamRlHDWO3nprCvQiVDKrabvV5sGIkXjqT4fJUcR9vHJpllVFUyXw0wuD4ayMcV
BpdpWQijHd988G8JS0AaGAAQZt71wuwHdagrVEDbh+wvukJzILJP8g+nbk8dsx4GH4Je+BIwO339
P/Z4skoIXPU305sPzGzl5AHRH+UZV04XbDDAMkAWaQdO21OR6BuJ7yosAbg+J1W28bu6kCU/5EjC
nkf1NPVyHiOSPIhIFkeZHLMGnbQtfm3oW/w6GnBueV00vqHUed/cQEA0oKL/E0tR57FE6YZGBn9i
jQP4x1o/YiA92SurlOtHmwf0MLBBwKYCNHnHPN4kQBRYbZPxldEVDsPajYAzzMAzL+EqOaNPKiIl
7SapkIze0p9tHsP2jrbdVHF6dd2egQHvkAOE7yVfW+v86+uxiHwFrghg6UmEVsG+qfTNakdL7+3m
q+IkWGl0vqBY/48sBMQffLudIo1GBrx+NiSlE54pE0anokUB27tTu2I7L+hTqyTO32yHsaZVouJq
IIeYRJXbRP5eg3+OgoisNXEXoPI02sGJEGnIoFn9OfChlNSus+JC9n1N/zBgR3Hfw3BTpSawnj1t
aAN3SSAM3Q1WMyXh7AZDuGHeTD1gf5GiNMgpHM+ABXKNz+6ac5wvmHfkeuKDReJ8jtfusIJFQySn
vmAD+zIkZ9Mk1UQ5qzxEUfgxBnlcqmnv/Nqr27sBL8J2N7culC+JRuMgLB/+wpBa6IngiVGW6qB0
BWOAbudQgDAD8L9cJ6LVnI8KPFzVr2naxSde36B2pOD0bwbrnkrd/INCT3kkb3xCoIBWtBbY7vYq
5e01Tp6DZaDKKPYVBIi67FeB3R7P9LxRqC8y+NWeVG9/GJ/M9tDHnVryL83BmvJZp9xoCcVcIT2F
j2r2yr61PhoGwDzBhNitHgcfbbcDxKaZIgKIcTkGrFNnu6QCm4ZrITfXmLhhXRhqHygKPA0SNfYq
FYcRQw5yj/eDIwaSdICSDCUMxDob0YI5Fd0DV121OzhYhPm3+pVuPS5a3pgElnDggTHKAj2KaCpd
rMPw+BcxsJ1agyy1xwjoobTQN+prhZpxTbDbD9PzXlno4TCzfYJLfVtlOewKfu18l+XZdzGcpx0n
5Av2xnBbcJ3v6QurjB5080fmwasob3GCsbstbCvzl2/UI5JBdf/vAgjLsxK1dpGKXwYQIqXxsOJz
t4AWKfuB7qYIAYxyFESgwl5HFjF/vRHfnGygN7bTYJsGjj1Rqu9Ozh7r6qEM6Y9yFXsiuPPGObmz
yhkDMm6+9vC1ZJWusJSh9usxIkNTmYyfXBIydaoS/5QRjTLu6W/Xl24SjvGihU+YG5x8Dva93F/H
oqR0n8aHFL0aUDjB8vcvZWt9016kPEayMiCX1WRa5cyjLLsBwxFhRSzEbQNWT7zkdk7Ea8An8CkA
GOIS5gk5lxspLOLT0wPqF3BZtepb4oi41o4JvSt8Ph2wse74I5+m2nAV91D8iBxKWLPF1D8Zq29C
eP5mKrsVeLjMOi7cVJxQazGx5mWuxHEqO4Gpq9qe41LIJy+2VZU5qKQFw0L00XM1UR6Jn9e16E7Y
HFcNbgcKv4s1niuVPmfkRrK/DpbkiYhbF+HOTCJtlXAJDCwyH1dJlN9MGojTboavWpyytH5uLrZp
pRGQk8nBbKvgzm4ltstIuMUdtJz7PmlPqc6IGgmfsYaI9OS2vwOmU6QVgMYAO0R6hKJdKap4tcKV
jAj4vDSZsysEj7REmr5qSteexIsapdx+GL7d1WTAXUa+ZvbNgk0G1quLKhwxm2B1G7t1naItnelK
+TCX0DXA+LXwrZiYrxrKFfrIJ/t4htGI6Xmgshbpk1slAdRXxBv930RMh4lA9gUBPS+AYLZrqg8/
O7Ne54/sXJavKcA6K8sHWNw9DwIHZi70Lg8klTMSotkpdHHNT6nXEFSvj1lylPakiHO1vdBLczpQ
u2wOxOdNuCewRN025yonEpH/CKv+4FmAQZHZ4oNcGX1wIE9M7Jk5uaHB1RNaWvV+oNzGfe/u9K+f
jJ9c31kBcmzNUASYD9Q32J9PfWVJ7mDBdBqKnoH2QtKGgW97nxdZsz3Gd2H+iMwdT9sLPGLSAJne
w1vcQRBC+RdUisXwGsgRv46uQo1acXSu+n6lGUfj/JHhe87YxD2MZ5crzXZd2kY/vOvxfhRYBefF
DT+DPJ4G/qJlqnjTFejLKabgAdHlM2vKEzzdrwibwW8mRgzrzQ6finMQ+18lBodf7vKKqiAhWVKF
IPc1qwz7oA+K0V13MqCE3Vl9jeM6WAS0Sh6t6gSFxkucf5rQlGSN/ghwKr26Y4pvhW/ALA1KHjWh
UTJKoS1JKwD6AgFfTrYg6f2nePkPT9NwqWRdIbEOsfyqU4uBA4GgLW+7hr69PtUFD7sntP11+X7S
ySV6f/xo2sHNMTnw24VSj9nxTPy/4pLvT/TRySOV9W14n+xvnpQ0oUq0AeJCL8IM9oB+TPH1bUUe
7e49xWXpteLyUKntV9IMvO41lvjLAMGhZBOL0TJEC4tf9SyhRUTw2smC2gJAfOxo7YgE1S5RzXOs
Jikh2de6OjfeFLkffobDAE3NHjtqtZ1Jkfrd44SOr/igcicq+wCGWBubUn5BYIUepuXM1UifALZc
p8qXm+QAGA+zCEEE05OYOMUpU7NLnuYWGnCHviDZE9MyqN7vPZ9QnPhfLvA0C9FL1SPk+oGET4ct
p6pRrvlUL9tUBsFVQcZscCH7gr7SmBlFqlrKimOxGzV+H/aRfbMPUqhWlOCFGQxv9LgoXicfLopS
0TJfO/XRyTN52nvXMu0pd7TJJ83KUtGGz8Jau3DXqfGLzaunnkQ3Gl/U8F+pAvtDV1CrpwYMixv0
dfb1y78aMEE+1NjGaU1y7pytd8dXN/y/bd48tWvErt2kfDWjM4FrI2A4BQTP8rDqWB3cUpVqrQMD
rQE4fJ3M1y7kwq1fsdE3iu7WUVe/b73Xaqh6sdYoCYWhB95rKngAw7xNDf/NuhBMYzLc4+D0w5Qb
VtmefgC7EJ4X4OV1OEYh1YQzI06+mt2QZEUhnJQiDlodAzVGu+0jRXR23nPnyXxYCmIg4dGI8PaZ
x5rL69jwLzhnM4IML15am6XDdQFBHA9OhM0tRV63FG6L/bb8VuPkeiC+HQhH3cl1reLBVhR0qsHQ
ndZ8R43jj9w+2ZxbfimRYLM7ZUGmbf+kRGc6JakEig/VEPKoV/asgF7VNClfve8W2WKrPMrPOZhG
pxAoUxclbDe7W/3391QHEteynCl3nbRw6DZdjFWGx9vTEGCHcWkPPBF/Si+cNt6iCxRaCXhjPTK0
Y2cMYPXKdXtka2+Ht3dsnmu+HaEoLXCXKe69vA90bsw3zAt9EiDhCof8De9A3n4ko5nJx2O/AEcO
c3ZOch3KQbU2TtCRI8QIG9kD+6pwASM4IYTmmQdsIlGHV+SA62nZuDW2keUrPuQlx7Ixc6JQlSPl
OndujGk5F4a40hO61MyW43tlLwRDJ69rdNi7wC5yPzDUorIOFLf/GHlQq+UupXMmB104aeoHphps
qAiBK0rN4H19g8igaqnp5+/23yWqapL6cC/12dixk8WCplrn72adr4FWTVpohx25MxqHbE/HEI+V
0TIdCrb3P58U/IfNXhoXbotMM4t/aP239bRVuXGc3r2iHYYdXhPHpRuGjpJKLJUQHUOPRR4b3MlI
Aiy3+69JdS+MAOjr4iFT1ks3VT64OBRjZkqyosQ66swA6i/RdU/vNxo4OGk9H8vW+mL5/Qdgvg3C
UwK2T0xllT+AegvBgrRNFzRi/6EZGrcH2+v8PcoXabRZzVZ8meXVhJX1C9nQRU7HXCQG/1O7/JpB
I0BL8JNpOrYt/JKAQDmQ582HEiEXsc7LtP7zQKfqkhsYOhxND9O/ukc0COXDGeeB+EsStyl4Rg8a
rZM6k0QTkinOBToiY+iqRG8lMbzcfloCQNjFK+QqebUVw7fUX0U34kza8twsXeCkVwZu+olHBX4c
lQd0L5madByrC9yJLWXmTZzIuyuiGjJcE3O0QTNWu/DlHnlR1sPmN8wyTN8NV4+jhTE4O1rIMBA9
RFvmc6nFOpy1XGs6T9v1f/3VL9cwgaP+y8ScX12V2LgphvLabOBOggCOBRZGcejfMxC39TVI3oNy
NgXk26mMJxTeKBdwhvTwiNK8WUtQlmJ5w0htvC3s9jVoPdrEv8Io7TRJu+majdo0qgt2shqK9tbO
aIMN+y/ctlGCD3Fm5DBa/u+isVNLBQEIPlIMjwmNXbH8o1BXyy6LTo/OXB8xslnjs98YNfO6J02w
sVr4YffrmPwfFwGREU0Fddi/hNUR0mxTEAHJqILANLrCSQm9SqZICRZlruZfehnwG3/ksJ7Ts+8B
rOC6m9PerW7IXaB6Gc8inTUD+OFgMHjwdKD1EoIuefcOTNAjWo1xiARzX4yvs082F0J6ZTFg28eL
7TrDcxQiQEUcfZ4F08LENuWvRpiz6uaak9f7czvTJwdi7WX7ByZSXlFnJfoZuiWQEwKMzdNlCAzA
AovSfcGrgr2i1QyP953k+6ak0R16eOLhOBX2/1Zh53gEKm3ZfBN6GMuBouu6C/veAX+VTUe4XdHO
rwwmrtHYavR80LAo3StScbabVf8Y3O7Xs37JcUmr5dhhDNYzmfDTDYftWaS21uWbmfLVEXo9Xn3m
lq2jrkewWwwHLuvz/VBAX7ZVJL0RZRRKKu0nhG7m0do/whwiOXVizYKyY8Tdrz7/pDyCSKPzDo/o
ny4rlzkOIXlRIDQj8WoZtDP+AGKcbfMZ9Z/tTiP9Eso1bM90ZXW8bDAKr7zODgpJqXi4RSouG8+9
j5LFkDxz5XY/3bM/2Xs+Z+Q5g/9hofMocugr/fYVgFV05e8kWzZgL3B1dC0R+ukJKYkUCA2ohAEC
4ol9tTFVQV0acSzo5U/S6TKzDZbIPWwE3WQkFkH8nnfm9+0F8gWDRu23L+iZQ2S2GK2LdhT3JWUR
5KsXFPySZmmdanR6E3xUC+i/Y78647gyRV0cUi+TjSnvjqmLNdsZSslIZMWC+EfBKIiv8poIT+4a
1wBtKKx9GPeT4b9g2/FkbWsN6qlTh5U5+Y+wlbPy6fKx2HHQo4Elzso7PHfZNGtTCY4jZhTKDKfF
JrKdR3Edb1hwZFAzRlM2OyrfFEH0DXgfqp95zbb+puCKDffU/XZUC8xouqrLLuI9Lj8vPh1ezJfl
Ar8gme3WvUWlYNAVrBARMdkv8CpNmFPK1nrtUP0sDLqbfOm9ikyMV+Ff86C1dU2dcB+nWaT2CQnJ
3kY3eJbzph061dxne1uebkvpovrS6l4uroBJqvjg2FgkyvpW158A5M2tiVUfyRjK7Lvg4H6yiGW5
Jtg52A7gII8spbg8gtGs3xpYXkzqbx2W6rPhGE9QXR49Ir6cgKDkZyQN+6vMCMF4IdejghBPCD0y
/csDS6iVOCljLICdwKYUzWA5B6T6tPJc9QTBLRXkou2uZJq6/aUjlnZPDpA39NG88TnTCgG/AhmR
xTQP/UFfktn+rICuphqsgM3RebLG4U6WPHnxcrQmscM7CotFtBuYmq1hCkC/bQJIuODpNKJToLrl
bGf5qXAwqovC0PaRdL4OG2xjHzRiAjOAxV+qaF4ZhtE6djvOVgNe7+LpyNi2G3GtGghXccTEARhD
eGALriYUcvUPOBaOoImMOpBUyE//Mbk3rCt4fCESe9uU8IT/goSQ+nBCS059KELuX+y05hVvf1V1
AbMe6eurSRbFDQ8/SFr8VgK0QjS+F+x48ymtRyAutxxO3MbPueqIFY1lKp2iI9u9yaRM0RBOKam9
AqBsCWGlqZYCI1wUlHRzhJZDrj+Y6EWmFfhbPkN5xVDSrBvoBBT+BRfK6PWnCWfNpDNsN2Wj+ksX
kzjiaW93Egha4gGWSss88fjQqcFYlYcsfN1+zxsCYPCe/3raDUyzGALX8zBLqkj/3d1lchKjdp3G
aInRMU6BfMLb2c7EV24S1/C/2UscVD94aw0yYSzZ1Xg9okero5FtAKBfjE3ViPQFz9eP53QEKRsE
FwocO7UBZ1kLuqjeupYozSAm54nZdNOhrYv4dJrFSWBMKrK+vPvaGva+OceAOwNDU/vSqbNvBKHo
705Dymte9sPR6b+QZIfURnlGADtRdNccqhifd3ZxrpsEnD5ZMYH/I1BUKlIaQ/IrpfHPI70lSn8a
cwJyZyCJN/Rkru3x9hk+zDrc2z/s5Obgq+fLSbBObup5831qCLzp41rHn4WldLEU8+hyb5bx6Pcm
RjAhcmF+hpCVKtX+hS+jRun6+JpqiCAunXz+Tc0eBY2sMIyNo7ahLDmqk8GEadK1s2ncQ96ebSKg
kEyRPw/K/22bI/AVOBvYcJzLvleG1B6Vn3/MlfgLvkbKV2anN8OYRinOz1b3jNx6E1CXpAbvklSa
51KxQNO0TtvGz7LIvJrQUf1EKTJEneW9+O9yEOX5MlU6o8Zw4gy4//CHYTzGv/vaUaGLKvpl/OlA
tV7W01SGiGOtx06VPONxKWKT3GZBwxQNSsNVVekug3alxSttci01bF/6UFIpT2cNTC4XDqEQO+Ml
vtsUbgM2dJdLDqglYPwiZzlgWNkPJoucdf71RZPupoZjNMqqCLuryqDM5oQPCLBA+PbpJosQwDi/
e5WZtBgyJakplD1P2DkupeSPRPEgDjCsewLjJBQYmkbjySxcI93RkFiBznvtJa3E3vMh4WLf9Nxn
34p5Jd5LGejD67hcADWaZVHBHS3PLcdvg9dzl0KeNJdhG6b2DuR3gfzmz5ZlJPXAmX9ky7UZpoKT
aGVCuSwQF7eYPPsBhv71tU9SEyhioqE8dF2OGhkp6aW7bHCRWk/FRaovQiProqDwRGUONBmUkNGg
FeesMmQBsIKTc7FcmC4GfcLtQixgZQcHwP3vkjaNhmNcZzSxixKtOpvdlh+6cXmzqqh9aTdbcj/P
7IT21WWltbABkLD+wrDbIhlL1RQvZdloCqPQp8XixuSKYOFEDt8RCsITNAVOPnwzkoDs2UtGMgLb
hotqIdjOvPVCoO/qynOos+1Osfv45HANSJ0OllFsURf574dxuK2VQfDgElxIzNJSoYvDQZDdrpca
uAHCj0RIv8kZoM0tWa4FIPpzL8QY9rXKwryF+1PJuhgxfG+l9/MCgMnUTrQvjf/bONXJFjDHOibN
/MKk9HX1ZQ5huizqI4i5CAJk8mOW4bY2WYq6g4TFV4IAXZZ4obdceaf2Mlhz7GzyYGNp2cx9X8U+
3uwSEGj58TnQXp4L8gpKbhjOidda1uOvlm40RtYPS676NHGvu6OvF8jEw9XkXdQKavCvZA4/lXjq
jdMV0ONqVIOS7EHEd4ZJXUi+aYukNDzbfMVdnytNW5xabuReMyOl3YV8oo2ic6ytBflvYdhg/mKQ
7AeUgO4pxq1daCUaXIXScQnZY+xmYH0PqA7I9YiKL/NAe4VRkXX6Br5enDqxXnPUEPqZ4ieioPbK
wWGfi2ReqPIMW5vshUf4V+7STHrjO4rGFj/4KgBKCI1IJYkz5pCWc+ZtNrMxpu8iImLLNfhKt4pi
cjKF9dXboqps8sbq7Zv0yf787AQPCkVELq1buVpCm5m3NEDiasDBSi2HlAi+T0Ano//iVGuWwJKn
FLDb0oDwF+eeML6AGW8JxB9ccU02oKUs2wNIekycHqbZbAHbX5LgNpRmN93npRgzkoamFEA1kUpR
AyZSncqAdYYuab4USRmlwGiRC2Vd/8qyw5HDqbmzJ24E+/kLLE8CBrinrdSGCC/xax8SQ2mioV1f
DCc8JsZuZuuVwtihLA1Onj6zI1BaoAvOk+p01v0PBxQVvTlwNLQpNGJ2NCHNlCT3CMgO201FLqB+
JUpHoj5BWc3EJecOvZF2mxDLy17rvXN3x59PtrhDEbZGhX6WfC+0mNqOXnKCB1a6/pbGLvvweX3T
9PMBkPPsMmoGTBYNO8LfVUOU+k+Dw7ydKpgr6qGuKUZy72r3/AOYm8WPkC67bTSJfFCh7UcY4vZY
c2D0dTHzHk7DCH8fzySCqQykNkCuilAfX1bj3GV3rwpvdZAYfzJ01Qu6Ekn/DqgbkU7a0Hnz7SHU
3pQYKrxUW87UmuSqEscNOSDutHrGDn/7nEEW95+oEO0kl+juaI02WzAcEVgqoeBYyYrxBiMHoghO
qju2nGT77W7rSf0DDDp4N2OjtGT89fwMsDumP7wLfoWEntV4kKk7Cm0bDRXMPPKDzRy3PYGu+urS
r0HObOfssrFlG+3n7My9TriBRFAI5BtCntzmNHS78PwR6/XjQP9SJhk8rWLVQkVD/6JKf+lL4AsZ
wkjicpeALLAMHmrr7Fufkm07O6eu5qiJBDfmdfqjrfEy2YSQXOXyAQaCGCUeMOZP6Yqxwex2j1q9
nuhXIsZwwW/CrmyDSQJaxQgdcsQ4X3lVnWBfTCcWgppH0OfXBOU6QertSnP8XAckpBRNSmIwUezF
W38m7qUkEzbwwzkLe4sabNNxFX3aKByJwipXQ9TA3rUbiSNYnqovE0hjYpFAmSnldH2mf1YTxBvm
+crFiUmpstsM8PEODOJ5zX9z5euZttbGFOEVGAnXkgIYNck11iR1hNbaQK59Ym41wnl/qWhyZzxH
JLuiM9c3nPuneTYHVhI48sXeFPkGty1e5fnKGkO9HFKZm66Q3nW890qRQ38j7Qi/3u5Z5cWiE598
OdcoQLvO9Rp3KEqtirQc4qXbdEPQMhnsUXC0QOIow2qAvC8s4vM1wIWDHsJDj0HWNGh1tPQC6cNm
LKEHXuFB/FV2QTsn/40G9Y8/rWBfYi2zXZYe555etrF86TyV+BPRUfc08eGOPhCsWKRMfugep+3n
MOYrrILbHxTOmUsX2fF26B7681EWNM3zCbNvyg2oRXOxYQQWLqPDsmWCRyRK89HrKTk69Q4IRDR9
mnx1NJLKq3yNw8R+wdRUM93QQEJKd+hfCsezPjJi9cvpyBQwdaqabaGC6USCe53K2cOVfpk1WMHW
fVik1U71oTpEPHqpZKFMypBuwkmpnPeVXPuKNg1EW/qaZzeiAifRv1EMZSO0jjOIroISmiI/KoHK
gGXlBBD+/ctrAoVhq89zK2V8e1TL2s9KxWar324gxSz76nipFf132idV+pJYtXOSeO8Dwo7Ya4Rw
Kkgd7c0rn0K9FM9YDJQAYrlKXzkHl9xb4YlO0ODdrFHkssTyCjnJ7cTCsufI8HVUsmadBmwWcoK0
Qh+AyRu9wJl27XUC+N15KKuUJxaDWjKWD9KqTMy3wiQwQagvM1toaWtDWldwbe+o0RmZ4+0NZb8h
kjubMJ1gSx6VqjxzqYizis4IYXPOXSmGxEmBiySSwycEACHroSclvCrhDtIiJtlt2LqEZVZ8OGvm
PFUfP9zcvHiOtr14U4R/CHJfPT7tXUe3ca3+Jzbr52CqagQLlnfAaZo6mlGjvKi0gWBo+uawRfq4
BJWEFarqwghW+sdFwz0xIlQZ5qfCeuQZ8diThfXb8QUjj6BVkH3QwzbPXBDmi9ENiVVWxCo6uRhI
PfKF0VdwU+ZlpIboi6kLRYtOpI+xOG20iiSVItFG0Cc2+Bo/wuznCpJNVIZNcfOprS5+Hefo3aIc
Bpg+Mb5kQNistSBeL0LoB/dkoO6546p8+yeFVQXev1OAFvuyi1iPcdk2soMpdlZU/R/Y3FscJ19E
cMGVJS333RtMnxOQa9yml5HqtSJ9m0jhSYzDRjjJT7Iw42hH4isPtLRcIYRwUCRV9QhNw8v+kclA
6ui5pSkBWDnZSUs+jaRMbBRIPccvRt3h7uhzndaUktHLJHRkhOhDtv+DOJxA+J9xLIp0LbgdDx/u
dw9LyHYDpA6i4/6lz8qlRDZjWv1GeV1ROXpLpPGQwQkcOdeYFMaTk+N1MRehrsJyn4UoacwpMpK7
nqCDJEfuh5dROr1J+y5S9FaMjvS5OcyzFve9HmZL2P+eM5xRS3YMZpbGs30jmtTUipx3zwbYFV7e
1xlZ/QbL7WHGBBG24x4izTchuBeFMfQ7BxDFb59yg/P+ChxgCbfzLN2o/bW72JZhDywcq0eBnjY/
q9sgRpipBdf/CsECJjOw3iHXhvISD4RkTLD9s2uasC46V1VI9+LpKtT6bPKi1xtL0VFV/7YRS9b9
awNPn3t8VZwQOF0NfY3zvLnzxaVylNqGpmSQUvqak07+qmNGvIYw+lmJy9Ylbw2jfwQ62iTFiDHc
2coOfec4iK2jz/N686U6RSX4YQOUZfoUtRX1dwPX1nblwBrieg9Yut+9fTIXzujSlTF5/6FLcIOQ
FwiagD12anr039NSvSGEZwhcHlrvjxBK0S/M75iWONpb5Yv8E6baKb+cUK8dDymZHQu7AGwB7tWu
bE5sujQ1NzV4nu7DLm+X8WdMW1SbB5imWOZbwfmq8CldZtok1X1MCf4ssZkcSctBJh7ZzzgwV2wW
7bMKZxKOfZDbhMFu2KGImaRiV9kiHu70b79lkzGVDDmNDJZpoX+Or7VbvB3v4Hc7v6v9xvjUeS1r
19+A9DIT0uNwvpjAxdZqd1/jyN8CXx3p6OJctjEwLvTlKyEsWhEDarHgslp4rfS7xmDhp6EIxn+f
Yj13yZLF359ucGHRmENxS3bLEAVftBJlpYetEKO8BKXfd4Afa5wpQfulpJnGcvp663vvaPo2Enhs
LbO0gd+qjmOhKPMo3yPUx/tdbWMPPIEN6CrKpgNtKXmT/U84llCBahaJApq5izoTOU+t9Z5A4Yd4
AkMfIf12ViPBReeWlCU4jcBHGwtBd1pWsSdqUbI9tEeCEvL9EW5XvBRsavbpUfQm8ZN/LocykYso
iqWTN09TwHGY9aQC+09TSWDmnhyMPGK4mLLQ1E0azJDCnxyT8O4QQKFvYn57la2C/CxBtnKyP3A/
Tga7LcWiMG2CyZw1EHIWBOslMPbCSLnLI1HJ2c7XxsOTjZMZtOVAjGlxRLxwQxrs4fKfDIA7z4/E
mliqgnbpvDFzOU3Q33Cs+hi8ap8KL4jU48WIKQ1LDxkRKYiK5npreX8+MleSeBULvVcxezw7nwYI
mGnW7eli5LEGt2Hf9nK3vP8xWEollWChQIkmTm9fbuD+pn4307HvRS7rTpzlX69345PdIZSRfAyE
l3ZD+IlRph5Uz0ySjxlnlwChIPDdI0mCmaHYo3gWUp6xzXk7RjMBFlimdNEoTdYZawdQwENgjbyn
oAvee/CUSJk83wWBXOAQ5E/S7HxjEFRTt/9XmRFRTGp8qqzGcKohb8hPs/maDF8ginAAhpV7Iefv
IQAx9PhaW2w0ePHp0OYD1i/HdLneNQCDI3D+/KAPCobtiFEKsSGsPL6s4DUSSxZQa26TtrZTk57W
5zYem3L6n28t1JgoujP6/mXiiXuaNib3TVAU30bxWA9xyjWCpe4ATLR48rCGlFqwJ/xUsq3kgs8R
xABcG97FqOSUbVL3Y7p3dXTKLHUiFKddsqTnatPYcNgjJvnWiQDXw4kZyKTyEvivFRVkuSSDBoKs
shW6ily2VaWaatgIpp6Voiu2xgb28830fcXuqy48OeUWdIP4CxL1XmU52CdcsAzoy1vG14Ebl3p/
rNlLI8iLPZTJgNSbraYKnSi+jLlM9qBahzXh0064a9L6hpsdyiH88wmW0Ka/xfxjbQ8TroWRpO2m
x5YZhQY8zrCvc1tlMwu3dCulayndWQQHN58iflpncc3vYRIqpjX8ElidBZyyY3B7QA1CgxV6mVyy
NrHMqaoEybHfz3VZpuKyrBaZZHawmM2sWNXyka2CkZ3CQQi0WjUdqJFSi4soPDp6juscg7lmcQRd
Yt4i+pgSiJmTIuewidl713S8wyAwNBF1yPheTqorey4NzRchFlo6Px3LhzMZMvJtnGKgMVxuNOVN
UIwGfQJ45mhBTRXeQjrntdTdO9HLrHkuWCbD2AdAubDUz7wcA4MYfg5T6kiB9vL84SL3i8mUol/G
lGTBJkWf/kmBP8kB0DqlF5AmxaOluc94Bny8wOGmJ050aW2guJi/h4n/TMX+k9lkfMXA90wFUT9C
QBqd+j8DP05CIW/SUjItH6c9Hkx1ym59ZvCI5U8TTUk7nlkaAmHd6HHRRUsWAeNOzRUFaSg+y/VK
ZjoKQHhLu9BoPHF+a2apn7a/4DQeZvbKYmyKHx3stPo+NRF3QXfi0sKJuTKNNCnHgCLrL4z4f+ME
9tWxAM0+8PAEgDTNDR0JaQ8h2WEO/k6045a+8jUH9BZSjOF7G/QpHnl6iDGa+6FEm+FKb9OkSIN8
GgMLZvmg2GiiBJw63N308Ean/mIfS3M6RHQ8hjnG6GF66oGwgXUehxI8DGCbceBfZdIn09ihwAQp
TL+0Z1blisQ3NQQgu1zPHRx09EhBoByIRm1UsjrAbu6/MisZiPZVeRO3iRGOCj21rDYB4Fzct7X1
mwOz7VXf9kJeu5+0L+rcvBAk19hxaiBTtfuCXbdc3bx/tAzYeuDp2lIqGouPSU7C4QCkwaOykA+Z
znwFmyKMgjmgFgUqdZtqW+jGv5lj+xHVTWj5bzR9rOIDmx91hWXxmg3vX26e0vBlpbmp2XYNob5E
NWMGdg4RCMZvsL21q8BiNHEI3tryX39H4W/efg7tKxy60EA/pIVs+6+tccrHgroPWcmHgAGli0+D
1QoWJAFsCG2Hmak3KkmoWKuV303Sx/S3RafX2p/0uVm2KvC7O9UnFrWL1LoD73UrdDivBL9N4fa2
0bVZb+0C6RKAeAUun2wsjUsIdPkINjms/OV2EuM5+N08T2qMKIwQjTsG8DAOGR0pQB/beaGZlJUV
vz6oZN6JxLDZ207VLfu6XRa8dF2HiuFMPCRTHTz0zKMKNRnFDZ2DFJemAkJIjvN7xeY9Y/rE3tgz
cjnWRfIPL5D+SGGu5gaEvhxxlFJ4eEX2HW0F39SKaYxsZqNYaapbistyeUv5F/MUSXUkY8n2Yg8B
ZtSIBMP8lju9jj/3yT7OSAsqsoxyir1ajYGTSJmQXN1j107Fhx+eCUCOtnckf3GmfHOLSN16mu5M
PNb7MWS88lKtA1PB++Z5Cc497ZOKkEJd6/HqOIvu+dv1DsogCAThaZjyzWVCSy88qOtzvjmTGCyc
Qgt7cNF/W/y5eSe/0QcMRDnA6y4Pnv4LWIzxpfmbIIzIsuHmf1KlIetwlIVBrzTrEK9McqgbjQOs
llbgWONJZizQ8vBV1CnMy+kdptAolD1dEsJ9peJrJFYBTM7d5jI85XwFh0TOwkG95EaffghARVe5
PFkGxb4FIRGwtVJ25uSVgwtGhkKXmi1BtMLjNnQMgOwbUa0iYTRnxcvZEZNd6iTX0HK1HqF0yrNd
Yump/4/CfeHr54CsHHxtc79oytuFCVigV9RnQ+zevkMGNQGftgkpuyNQhbDitZxdc4RMp/5JO9qu
78ZCYdBYD1bys0HidtbZ6xJaeqVk2O3leG+myek6ecTnMX+um18ClcpczRPSN99z7kPqizX0AlVC
bP3oV1VzMw3JYFKiFHWJBGOo9AcyzhMYmkEHeMSqwA48nfnnkQHYzTC80mSlvwWGeFiOME7knNiy
fWvo9XIao2bI/PPxZGEYaS0P/J733GMVFgRkOJW7MMkY15lHYnBnKEONf7Yj/iAULoxVPE7dB+FY
udpea/jNs5nQqWo2VUlvOP8e32N+EQBCLBATAlACThp3ocDrChaRh2U5kCf0C2PBOzD7OIJsn+zw
7aWwpAZYoGSLR78p/AiRE9pEJCr72E9oBLTElcVJIhm8FDd75PLnhFFe7RIXbjhKW72RyaQhFJH0
hhjj0BwQ7vKSBaS163nHdLgcEooRCssYZwvFtGQLxKEzotTQmWasBRuyne4MfGAF8n5obC/4chcr
WfGs79f7brhPgmQ+9kqKLs+Cg1i4xXm8xn/GXQVHaC8AXl/R5Cv13UKVgOKS/gwcgSROlr80THVd
h34J09uMiWwjgj5MjSDdBax6TpTtsyICXY9BYQNLuxVAxd/RQTlZt6+dpgQz04B6HOWb05yYD30i
MGFiS5mZGbrpuO7U6m3Gt/07rZrOxxVisvNavQ6hXhypiY3FGN7oc2VqTovyIbL+Arb4+mhfOWO6
Hp4/GgMjAAqh5WK+wfOmXsxjPsRs8zWNPjDfoxJmWy7TwvpYio4EpTaH2VWdpIxFxy/Sl/uPO/CL
vWaLBZNowDgv+/vnb6jqNaw9jAOPJ5k9KKi36gf2c9TZ24k5kLmTnEgHL6TGR/xjAAh3jQYk+UlE
Qs407OAHkZjtNy6crKnS1s8jlDnwXl6VrP2EwJz1J/VlZp14pj7r5YrOIJ+G2zKdS8YeypORY2I1
asfXnPOFFsTPuTTmEeK8CQNyWmmTLHtMxCf3b29SgPSHdGRr1b8iK3xN8qbxJhA0XaWKty/L1VQC
QHQOte1A2hmhxIcd8kdkdlTkM0MzjEoGuEq+GdGQ1PEBCkUlPuotPi7KwaNIjGOYzrA65W8/KVBT
VjrZ7QFUy7LyZIIv8h+JqNS8SVmJeweLB2qLNHscxO7MZmHXVxxWTuXcLe5t805ngA43ZQgmBYN6
nhbnDk7QoN7JlVIklsk9CwKbFz45oSVllgJX/M3cIBlUWO4FhbS73Q0C8tm+vTXct1497cIYzXOO
VNOqzKFNw3+PQrfSNlYJBBPGaZNdMFa+8iKm37aDSCRXg9RW0Ip4O3WJL5TOeUGxg+/avDfWxT3F
TfW9lcKy+HVXCOeBj5lGa14UBCiWM2Sm3DlMfkhUy09xHrh6IDLJoVoYBcs3HWwMadmLFbj0oZyj
ykzWudc4RwfD+rvZ7Bs2ItAJXiJIU1LiVvPhGUxCBJ7j6khfNfgd6Xs6McFwLg2UeclKlFkQI9GC
lU3FEWulFD4i6fPcD2rvO6QjTO0dxKOIu4EiNo+upCSLFCwsjMDgH+u+rbv4cFvYFruEdA0CnOTK
6RdjaZf45VpBI0QcrjykhUVNHhs6/sDVOZfDl1Z6A5xFL9txV+nhxXPwe5oF1kBQGCnmCGixU3MD
XYQaqWE75jusM4mK9+Z+5wn9ArV/1qu5QeQk4Pli+5+9KeT/cQduLnRdDkYZD028aW757o6nSaGv
/b2/bxncNzuIcdEGKkMdeyGb3G5/WPfLpBWuZKMtmNNjav6jDSA8Krt9dcTTB6G5XJNyRw1oCspi
2a739OoNSK73LzhNY0Ky1cpew9stk7JlYhnYE2OXrhPYRdaT+16Yd0tVBnhJnL3377rtHaWwnuV8
F6SP8tnfXhrnDZZ+YRi207NkeCV0Xt6KWV/fRsTQbtk20/iABn0QvHVMjzo2pCqbD0/LTGXTYykE
7hg2Xmx8NPJLMEFTXn+14dCk06FDuNc4rsmxUR9O3PbXlvg1tfa85ESz2dOB9pwykoSPHil4MJ8e
6snZyqQSIgC07XJSm7In7YUYk2tuPMT6gOHHN1vjKWPEYpbAVpwoLV7/dpwRZmG0f9wNowJ/0ckV
Ob5yVW5uVCcBjBrpYUBgch8idOXjazfHsDq9ERltAR+c6hPsMNp9n/zscUn/2he2Z2Aisavo5/1h
WjK4NY+zstjHoo0mvqpL6iaJWu58uBicak/gP6h1JED3IlAWps/agCKbIHI1EVfTwOEiMusLAlgb
8G+YyNyoUlx7CREW4p8LPHeDgkY/HHZJJZPS56W4ACPwEFQ8cC0MsRPBGwCmSjy0NLLoQuwZib2s
pHUnJwIQvS6GMxkDbcg29zGWsZs/59+L78es7jUy32k489+CJDTVFRYfDItaZwlOhlHiTcGRWCwk
woIOqGpkO1LzLbhyPCK/HgaJ8R0Lspxrq5cf0aAKrt2XMVJvhOQ8Ao/6EE/hEOV3dx6FUnBYBCZf
cNnhAvCeCqRpCrFy+vBFLkiYqhPUKpZ6SvG81qbPpu/g1EEmkKhgyag795gH9iViCSD9TPE+//pL
YCogCAQYx64gZD0nrCsp7KTxnwwIidvlWxP1qr8flkGkiG5iQeCg79qpc4Yh0FwIbXoG6Gmax59X
Ao8pIckYiJUW7UQwZ0Y+guDS7FAa/ma8QX2DT8flCeA22+7hhaI7W1XZoPOCMADtw9SfODQrCMp3
LeQFQaymXxoQ8X/hzEYP657nAjRN38874OT73ikls1t81L+HyoBNa8VK4sr8TxsatR4yN1JDhSQS
IrHPKb6AiVHKvJ4xd57N1ZGNX5s0Hz13oFrYAfgSeWpYvCveAp0h9CRXxz611zl++vi4mHOCA50i
jc1HpqKvGsyMDK8XLW1Gc0dtzNZOrIt9026M2N4g3Dv8MygX6oyP82f5fRFHq3BJGn9UDinRlqGd
Dvz+zK5jwbDCpGpYi3LeDsHJt17du31cDMe9hwYukzUHC94ROJgOcpHo1StXT57jmcHl3kQNXPwB
rIUuZ3PAe+lwKcUk94eKtGXEfvMDJeJivg1J93sUCIi359CPkw6q87QQ6Cx/3txzjb3EzX3+9q2Y
gvGdYEavAeFsESyjnfyfsl4BuRygTbmS8RnyMxwyXgKUizoU9Maeod1jBm0zdA0icDVpzfu4+zve
r+Py9AZlxkQpKKJtj8DxHv8NmrV1qiMw8LFTsD55uScgX24ahN4xNajVsRHC/qbnrUErO37SSUCF
70nKV6YRMtdP0fgy7OksemJASZ6YDVvoOkpZmtFySyCHyodIMVDEFa6PTBuHVU6h9uxOr/ja1XQ1
mJsJmt+EZ3uqXvyl7VkDCEarvbur/d8pIJzCP5dvNt0EvYgi7G6yrtxNkHNj8zdjqeGi3wOoREOX
lvWPPrlJNlGHui2Of0VtAusqglGCzj3dxLUoTmIKaEMVvYox+TapePAxl+fDmsO9qMmyZKhLOjok
WBQv9L3NQIhusznlHCGsJGi6y/MncceCjcLSeuylmcpvoCk87zIOTRAZbuNCtfOq+oM9t1nAt448
mi/ZZ0Bo6yowB57FA7cqBRar3/mYZBG9MhQRGDNgC/d9LbqLGqvQEISYk7bHJ3SSvlez1oOZAWhW
cchbwre/oqNp0zMacm+rPKBAsPjGNqSKvnj71jy0zx7ly7tDq0j7/BwiijKSeLNCs8kXKE39f1cG
ZQNtddi4IjUJWboHyesxdV0jhrRvtvC/1QRQr4CFsoiMjxEk2DDFtl9DVV1eSrirbnfXSTZwieY1
vz5QdIfMCELUXbry9HgazLtm2C2yJMSONcip0l8+7PFDRtuAezoRMy58PcmM60vUgm5MVlPL68Gz
FV50WPO2ZuiovZYh0JrOjnS4Mp65m2Uy74tQDXII1JVvMEnq6eH7dFtRYBnHzbqsrutkEgdvA+v/
LblLPMV3pI9fXrakfaAFMkv7zhIh6/5itbrDzL2LuBaK9avyLohq9nn32DO3BFr+S/wxq/RhNw39
BvMGWC0Kgpz6ImhrCv8NgXcofLFI+IAKvZix0q+FCrN4QXw3wzKtH0XBfLl9iTaMDxrz9C/9p79J
12mzj7jLJKddqIJ6etIrn2CyS/xem/9VEmBEQyusm/dVeXcgiMGpnH81xFXJfawFSpFdbMKvSo1R
56KIry3KNTIZvQnBRIi6VnPxLh1HXts/7D1HGwFS7BYrsZde+KIBUMj7gL57x60cgASueunVwEgb
x9en9D00K0Lu5mUhM8Xm/80nRGah9ypqVuquhBXUb977GyrHU2PWvGcwjLtjCJ8OO/2yUM6k4XSt
7o6h9JpPDxg4oabvMW6AVh4adS/TWk38HFNqlgkhiRKhmposLyG510y2I15HdI1ibVXSNwjpdk9Q
T5VfAZm8fYROzvAti/+8X8kCUK/zvir35pxB7azKYzxNm4fgFpgVKWGyt0h9HswNigntN7NLmbcM
TYjXZTGXbQfLo2vyZIDGGMkjMGN5qRK/FbuEYbMMnzS6oLvG6q4zCGZiXGrWplNbPUYVpfMICT27
FkIMJG9pjRyMwcyPpTQ5ptwWqoMpOTpdYO27G+sogDT9obj3qBhbpmwK4TWIkYeiiA+/H2XcPRyu
Sa6CGex78nbttqB9toplAtUz5qCtX3gz4mWVKjZk79Urtp0Dm4PWf9Wnmi3g75f4ye+2TznQ8rsn
s9OV5u16WJLq3huI48eumFbFxJjkWK6h593nlplggA2XlgXrnc9tMXndJKZKaHhgndAE1aJ/7tDa
Ca8CImLTL+yykcS64UoDCeOKILv8gImr5WDNA/mXhxMpwoQHFD2N3FpB99sstCoL5WMuQwnPvxZn
gN00RZYXXkIj35HXn36ylbxUTl1La7tNcqh+x3KXq2k19Bb1yzBhka94s93v8sZF1TA4QhbPf2tP
H21be3S48ZB1TPJRvYq36Ervil4sCnvu+5RWb+tOyUmQVgwPeMRWIBfIg1FOiISFtSMzIPTNyN05
sl34V1P2rQEQ4f7qu/XbrIVqlbXcfPG/OFxBpqu6A4Nm+UzldJj9+yMs0tB3o9f037N2YdP/mB+p
VvdvNW3JfWSdMKHnkODABCbYtn422oWb83MqGMtwTp+jw9RT/sT2MS5D/vtVX8BhrNTiwqnKITZN
sPBYjkLkEPsbCxAyg4qm8xLhhbq7daKFOEEtAWYwSqo2fIh8NZEvzdPMigYVamVZhxfrOZv5WMdc
1mK9dBPHd39iq0I75x7GqpfS8jXuisZ7vByeu3HdOvuUarsOH7owk1+Rg8F7eWkiC9qPqIwwhgZZ
D0SDbaF0cc9unsxr+AtJtGKs84/ndKd1uOe3jTZZtmTwDipiOZOUpwPPny6MpraNYk2rOwqO93Jg
FLsj+5nC8uHxpYVUs4fJJcdNpJrkOTbr52Dncgnla54Ng1J+edBYSe4aTCQk99N2tHJKt5JaOE9N
2l3wb/1wfN5pbkjXwXQTC2GGh8mIeGTDetArO1jBWA5USPdGhCaZZkmRNILpF9t6W+ju2VDpcdx8
udzKwcdXzu3q4vkcVbS/plwByDvSgkPBSv5iEjGHif5H9wq5xlBESQnzREngfbDLwG0mFY/wfXCG
dpDBgFIV+XrxL5zwh4TDgwmnkeAn5ByQ2xah5Yhh14oJBzePrryYHLN/rPl30hUGzGyLCNfYzx4z
IXirbfIbRJ1GPLZnGBTS5bjc3pmTa9fweyI0JGVgBsS8/VvYgftiVoBTZGX1GJxuy1mdyrdYtrFX
5UbeF5ljCDNPyYM35p83BveljKlf0Lyu+oV3iuLOObCF4sNXXyRQI+oPPMByMEsgfyEKicXzYBw5
tv388m5ww2Ys4uRG7UT8k2lYviburhHV4obRn5TOlmkp8wgDmtLVQz1VlF0UfnqSxsyF8yroMG3+
FS0YyB0zVLoIxQbc+cbuzrfe1TSmS5ublsBxf30UIdXmtEhTSm+zNRZUvbMbOhPxsLkkg6240xcg
jYjvxOxtNeCJlzxdcYSWBzn8TIFU1/hYSShkKJN2ckXBLgN2+R5HGwcmKbmkoJRaf0FQZiQ1JMsE
5C9weEpepIjjd5TQLLZhnTYAxfwZ6a63IZX7abAeFuLMeTlP6xLA3JGSNe9U2e39nJ7ooTLnfgAy
DoSvUH1pyNOBTYgOIaZwvJrYbv32JZzUg44KAnLhksKXMys2FuHPaxWljlsU/21AhpucEeFAiSuQ
HtVglO0GfsIZSnx4L/3caLOYE6ntrb6tUfOqppfLDZNjYdC5sJ6fC8e4E4CTrzfrK+XyYauF5F6o
M37QcWGbvnqBtTVAHusNzws7jxp6kVzdfOH5wJArxMYgh0F5CvJUM0Md10JJP5RTv2H6JBkJrgab
2qfoJdgLTGAgyikoeUJqpzu7v6hCwdANfsm48olzrkMZAzpPxrghzJ2lFvdNT3DICjRbCdK6/o50
2rVqaT9UHI4HLMZtY05rv2mmMkpyFBd3LLv3pj96HcOAq6Cbu/BP0PC6TpzgAJuFDxAQWL9cDEw7
lSFEB80Us7grHb5OxVgJ8notB32nk+PWnEzI6ZTPjsJAvD46Yzae5pOY8H1XJc16PPqA23+MLbYf
kgUzgMAcDxH17vEFVYCGHiu3F9mzq0d2V5ZKL9QaAKH9iUBjF5h+OT++G3OB5NnE6uvMHZTv2lCa
x1ZzFqYCt5nzU2Ht0BdzfG808mDttF0B2GbZtPRquWN0Lo6M9prj0eENOIv3L2Dfsm2UzItp2xgC
dCuRWBMot+xllREVUU1XUUb7Il6q8/tZtHBiHQtw53Grsozh6dM3KJghwgFW/mjEdRCfxnC6CPcL
8aSsQY3oOdDvola9miCl66ExfS4rtsJzzQARncvgg+7OaxTa50pkUb7fzJXSXaIYJ/vRU+utZrks
TybmoTNbNCr0GtxaQ9dcQQ5MAmOq3nR4D4UKpI5DTlr2ebmd6F0dbcOf9L9K5nvMdVqgjfVxPsIr
NVX2cQcaccJAZL8feXP/TvIWQOF6RRo8Ej62mgepJbf44NCm/tBNWg19Epw4A3I10xWdXl3VJSlq
kWj4ft18IBYmpqhcRYa7V0yMYAFft2vtDxItXyt24CfRewuxyxw9fpFJN7CPhRiTeSzw83Gjk3Ar
JU4B8F1UUve6a5YaOFrOdiTRw8RE2obrHPAgLJPZxlAiwpFSuDvO23z1RRE7E+K43zX2YIL+uP3o
KEf2wzK3wApEQWVgN6K4VmblAkhXYCfjxJhafwgWGdN1Dz4mQK5qufnNr93OvrZzdCOI8GYhkhP0
bIa7dYLYcgWxSX0mke9adoAfHmqfefC6PV6Wzo7z0DZIy5Si2kr3zLx2fM7eN3tg+0x0rbIos0vc
ad8B1AfhowwcVPoUei7xUf68ACtb9F9xuP8aWQd+YPAicX8d5Zu3V85auQ9xd7q6cT6osty0OQnr
b93bgTd31ImFWAvNi1H2KprWASffEAFWnbqGsyS5/64o0ki1wq/N9C9jboTD82mDuPZg8Zbplc3F
cpOHqJgf8iIhmzpcbZuHnvUWWIDZvplSgPt3p98ZkTqR9j6B1ZzZ/QELi/idXl1GfE7jr6AFMt58
FqpfYc+4mwYafEKT9qcve6AdrpvhV+ZsyCqeVVHzfG6d3NVu9POcVbek4CjEZ9Y6S9VrFrCa2ok1
t+3FCNvOCC6KCHKuA1a6ugK5qtwRTKpBHaWN10W+8HzC4lVypsZNnKTmulWHemkz7yaXBzmrUJ4U
//vUy0xZdpgMHvzSBxG/dMrGpZR5ZIz0keGDPxS1MPuaA2Zbj8QMK2pCvPSX62XksSdC8HWkF/oK
s5RdO4PjMKd9Rh0T624sDfIBTzmNIwC+UASNsjNA+0pdp8sRJuby2q/ZvFVnwUQkhgtrsoni7d3E
BfZWFC0p9QjDH6H78fZCM3+aw5rJIL2XnPYejNNPQ6g7ImYdEh5cicv9+NG1/KbmCzaqqt3TOPNa
JhHn+NZCNbcGnfKpHg1QbbZ/Alcm7Ho3s3sVrbR8LycmFkcOOpAoyBGtUTpNJAfCBUETNxpplZRI
hO0+tpYmeJVdld0ccsbAcp60JjOfRf9VABXH39pdZrCiIs7bFR+p4SXCTe9ndlLbQYHZ0o2CBf8E
fOBKoiFGol5mfPiAsxgPSPVSwB/HBCOk+4YOJSs99Wt03DlocYnfeIO+bo8g9W8sxhlBn5ciRzXF
SZt3dskpT9E4KVqFCc4H2Y+fG2whu86fjA+gvzA//sB2+gt2det+n+iZpO/35gwHAZW/GP/FamjR
kVnVhqVvUNaaPu3RsfJbxy7jPyxLC0kSzQuxp6DD9+PYVEVC+0HX+M+flls6MG/BagXczqj3d/+U
w5flcrW9tYsfLxFgcwKatu6Dnsbhq5O0BveiWNWf5JczQyfEFZRUIfuV5l5oK3eEbLBoiKN4taCZ
kNnf+57yZXmE4IwBR76w+UF49WhBt023DIuAclXTh+DDrrdCCdQVWqJS11IRVkLi8lPA3BT49T4n
mf/7H2KbzsDfyeYzO1Ht+N3atThV1RQ0GaDGGSXJlZ2VPneUDIBAG/58JzfdL+GyE7AIp8ZeQ5/F
AqJPpPg1SCzpjlfQQZqwKFjwvuYwOw8ixY2gFtagNnMYrlMValwafREM5R2VNEilzsASREGFB9ND
zKT2MNoOZ+GeJRu/TryFAYwQ2TdkzQkPpX+etyUZoonfpbogRyXlzxNcc+F8NwjysIMgCK4mZSWo
TKHK9cocv0sgd5cD+ZpIV5ZpEg3V9ptkearuCZL6+hESPbJ+3ioAq0RYFSDPqqGe6+OiZxAfAhee
A14mx0Fo82NsYDLGzJKCgGscKqLRG8VKQehNdUjJsiz9eoi/96xp8cX39YA4crK6d5Tq0eJ+1jo2
qQCWs9708/dAewVM4Y378kR8r8MSSz7LIKa+vakM9ijtRrbxzOn9o7ts7LtSNXT811EfhDu68mm8
Fh/VIptzLS3bJoKl3lmfbj9Wbh2e2Xh7LwwdYNrIJs/f6Ib1A49wbrAT7iROHkmL15GPcoHf+ogx
IUhAua76ht+vjj84CvfPyRhyrCFBhGLxXNtenvHalKnFZU+f3EaELuGHGUqvHVz/f736kBKOWFKa
csqpfldNUuBKLgmQkPPUcodHZfuyGCFqAwalboCpJyXalbL9aFtPzSQQsxs7t9nkKckM9jXErur1
wXneMshQ/TQ6gZ85N473b4z298OPggMDbACs0OxIWrqJ4/Ea9TUYY7/MOEvOpgHf40GTMvZeHDaP
wcyekwL7N245uyH/ZAoyYW9P60YDJbZh2yaSdvjCUMPT2nFkNYp7ANk677AiGDu8dVfISWKX33gx
WF4bxSRQFPQwFz20+15sHHBVdcLjaeG2EASCF6KURZURh8v8rdbeXOETYZkljnJirZzlg8aQqyaL
5MhrjtdHGnyGz4LJqsvo9OXQZ7K1pL0akhGjSvCPAW4EevDa0Z5a5HqAT42o7MoQ4f8baQXgL6Sy
CesucKK/IQPNPC59LPSuEaUzTgBTR1eyeUcV/da8wAdBDe8EOIjgVOAX4iXhnM0eLfxof/vjy1NM
2XVnnKlxKwMkenzql0L0Gb5AR/57NBK8H6NrjqV1MNWJhTXG3bR/M8nqbSO2TXdN39IpW2WFZADX
orzmrJZ+pQ8/4frYrqSRMU5ZrkAFIXlI+3MvQQl7NrKRi61rIPanj6SG8BuKcmkw+yj57VgEZFYI
+vtwrLXVeuBljm33H6LST2u4xyr3AkwfhKwr6MqfRB3DwyYWIQ4gaKMwHg5SyguN7u+Exj5hray7
lRM7E5XDstivteDYoPWIaHDlEaoKH2rml0HcgT6J/6YwzIIGnrr1C1FIMYq1wTAdRUgbh4SMwVOg
AGr0+56pE7LJXu4sfTaRQQRbGEZ2/0LJpyfIlNp5xBteaOT7EP7QFt0pWaX4gnX/C8zkXDnWOAQy
b7XCgYCo4tDELVYEM4crF1u0vFZ3TPI4c69/QPGHX16Dzhm98EHRnHV2x8Z4X0QyotT86+0gdks2
q3+AZkD814hPrKPNC5mE0q6xzXac/rtpvo3mYJRfwQcBHzCNbgqub2jtqZ+xo9sYWUoPb9Ov+Sno
jwI51hIgC1k/0eTmZDVqSjcAejmEqbymmqvLozFf69joYk70Ru8WfDLn0gTUkK8y2d3dae1zCQlx
/Vq0YWLPtnMjFluKHOKkoTQ6ZehtIkhnvK4xkvETayQKo1/IVdYG1A7yVStsqnVWwj5lY9IRsn4K
DTfb0lk6SaWhUCHqXp+9l0/1I0rPSAERipx/5Q2GuU1dvuyqRMNjxTcKJzyLiSyWhv08ifaiQU1A
4vTkIwI7jjiZSVZKeeeLw6LS98hVnxqGQrMNx/0aKAtGqKgK9E2hy3RR5uKe8htPHXN0zPiLvQxX
lbRqMz6eJHpdat9OMsegXjjvjQ5Eveh0JseIf3qSswqJG7019URXozJFN+btAeOf2WKdatds+Rv6
qygSQr3+/mzpdCrHFaTcRBZ8LZSyUWwzzIspikXy39xw1zqG3mjXE5u5KIyhK1cTzY0sLiVNe+0r
i9Y2nh9ZiyCYf0F36z22609maYtzb4voRq8HPPMsee76raDgduqcQt64sBKLRQYj3jjgR3yXzIhl
q05CofJyhvCYAyM22cm53Ua5Q9W0b+TDsZm+avNQFFeL3LBc1yHILzMkH7Aw1P1if1cVRJzRp6xg
mZhGutZ+y/zGDzGo8EXlBOEG6Fco0EHhUGRC4ty1ipmNqzFP5Nf9A1Z5aW6Ay35zW1l+cdoyxo+K
iVBSUeGUb3+LKx8DqqdHLLlTXwTS4t/XVGp9MJkrfIVaJgT3TvJRebZjjc298dWF/NhuafoVrCis
u19CkKLt0a8F+ygZrBCv5tepelqdELYKaKfakweuKbB7d+y97+DSl9VviKcnfae1lOBvQKGTKH+C
x0zYkQJIwz4qyVjYLGQPfrgIyQC5Am9u9RLEaeDvX/11zPszQvX6aWs5uWY/XsDjm0DdU/iJA02b
LN1YtkEyHgifVr3IX5iuPSp4mXwzclw/xg1yOTLWor/HIklyOIV8oCYaIr07RHc7e7TUUv0r3Vyg
98kJHRz91PIpChMZkl8H+f3+UE8BGnWmjs+hirJvG76myxgw55OhI48QTXV/EyCNt30ufP8K5bnJ
mynNV7lxlxi7yKlax9yM1x4m1y5Rym1CG1QBl6t6tfhPWvSUeyHcYA9t5mcabO4rSqihi5Qo3G9Y
LpMaDfPTwhPnSr/gx7cqOMUONqPCsnxX0Y3CK0o64F1hHqlp2RZ5rc80yS6Q7sUq4Y65oW9U4Uo/
FyccmEZmUibUOA6xQghhpsb4e0aypo3hUb6328Jnzs8VaM3weCTVxv1+0ifggeuvZYOmehJkEG4Y
FO56Eo0pS+5nqNLt0MJmaayw67OCM0ZHklj6nWINRiEPUp4QKeZuV7fBW0ltq42Qwojltg0WjHeI
xkse6x76yF2U2ppRWYyoFmERtKqbXFNzcScPOtZ53GsnDwu97FOYPidrwMloxWAN75OVIv2htF/H
Ww2MBBK/v0nKfdWaMr86ElENHALM3XgsAzWYoSNZjspSKz6ZN5jvq28dS8xgNjbKWp/9SCVIIbdH
pmXcvQlnQ6mfs+1v8Rml5e0Eq+kyAOJ/OR+mkeoj23DD/M4IHjDXtMsu1JF6wa5McL3lGQJCCPxh
6r4cju/ewDukHOEe5kkxpWggzRk5J8lrzcxNLmY30DRTqA3SksM5zqpOuIQC0/EyD+ofIqNmbMJa
wGmhrlw/hRcu9ajRHzYMBSUwX6lPGkZrb1okwo9aUUtzw0AY5hotp5mFHoK1p9JysSMAN4wX2Om7
Wxl8/k8bi8/gU2803utJKYpe2AT2Elso0YLJ9fYirMrDwlM5H93uIJgCqXH0H3FjLD1Wcyzz7X0p
+5o34Z3MyLN0FTjy+YhpRYz6zS4aBIEy6d+/5RVHAkyWR0RQJ165837iqsj1I6Pvtxw+MdNqarfp
N4MXyVcqiI/mYC7xU58i4gLYc3lQxpRJR8ffaiW3i0ASciUyLUAOOX7GvXAaKVhymiCIMamD7Wif
HhppaTDRHRBY85eFbUKLxvdSwSjje4LtqV1Ql8HLPbk/vd8/4nEmWUFwd9S9y6o0/BewXiT9pqeK
SZmNpB/WIf8f4hZCPao3KJUFoboxcuY2WfOZ5mDCztnNwBbm2B4FDb+DN5za/UzEeftYPe/3VAiX
JX/6y6rwj2jCgc5fvJIy3kyOwX8qvnksVxnIPzEAjv6tViZhXlC+/Czw49Z8RVpaBepMJxGryhwx
2BIwnwGwpsoN00EFzMcrZvsifptEoSbn9YdKHA8SC9lSDdDWMBW13sc7QxHSc/jvIXtYrl7eym/g
05Izq545uXTgprHjwe9At+JSHLMhBBQ18WVmgfW1mlvv6RwjCcFN7NkLIeIxADtHLb3+DFcCxRWz
jV9f2Z4CZN+C6RkbiYF2uGKMZHTV6a8TQXbG1r9/oOJTeE/V1AFZ4lzulprqauGEUnmKXPm+TJtM
iQUDI06FAPox7pqiQwH/iimH4V1cp8VOMfp8ZQtTaYFfIQJK+LdijPMa7/fkKVS49fPlY1mudT3K
QScm2JXpj3Jpgr9CJxFnwxsdKmxF4ZP6zDmWCrqXfu19IeFBP5SbLReBtTI37p0/gL4SDcqxj0a4
9IRy5/QhtOVgiSY9C4X0lp4jEfc+MwjX8nae4Dkkq+LBgLJkMcIpTM2aG8IZ3fCQSQW2yVDUX12f
yW4e3Ea4oM0K1bzJ4hv07MH7zulNKbTyvm+nZRfYbaGIrBh0nmB4tS5sWuDSWi/yLIAviboRtKQn
0H106m7suq0RJs4qif2wdDMSFZiflZWuCFOpzsiRoH1KDBLe42LoWOXmNdAdWIKaEgC+0YXhmVA9
6rCKy+XsvVo4h0LcjiG8l93WuJBPGyfi9SctwXCZjkqze2gzp7hFsvaw/6Rb3m0ept5G5aVPjRry
NTow+i/se7zGvHujol03n8dt9ApqrPYuPNs/qUUN34/Ti8j2rluu8ST9i/tfW2kQ7GGXNMeWhVqw
IdtNL5hLMVqd2QyLJJUnvf0Az4nzzzIBYzXtdh/qx3VDdJ5FMyQfqKOkJoBwvgdI5KGjM7rEkBQ7
31OQ1WjcF5KuPq3vwnUuK8hUxwy9OJEaKnLb6vuysvtEo/RaQb2gD67WR6iApTDqx22OHoNsnT7K
TinkYxDYolmosVI3d4bdpMcV9JSDIJFe4yW29hazQAhGUOoV0jRQ8BrcC3Brn6jP3Rf+gkv9lqCZ
AOth6fA62q7uOnrRPFJOSrSt2KVFKB6LYb9PBjHtHAFh3sKtrAL19YxvpPXmfly77hMUHsl6IixO
AMRCkvRGrrymNFoCkXdOIDYIt5AVFVo3/DY9r6SX//FLxaeczL/QgaEIb1Qfvbg8B6EVyN/oLOgB
dlaVcqpo6ssmVrNnTE073b7Q7Bv55SwJQ/elf3TRmnmbaY5rttEqekM2AsJHjWu7+eDd9AfYtVu+
BtH3tceOs6yrrhn5iLDh5A3Lch67DHAPObYRwYNJFoBD0bWL007wQhjg6fxQKsmaIsibF1NW43Cm
MrwDTRIILV++3NJun/8cg13aOiv2NMc9/p2NjoZeHnE+bTbKeMZq6KSnak4gldPXGRKrxBwq2hi4
3Iyun//DyIoK3mps/5dbiULAW7O5BoMsRn2/JWx7jHDtXik372lYIbXI/7Hyt0OzmgbUNyfvoH8h
vKdl19Nl+NEsVSdELv87vn0HHUmq5NP+2kwzsL2AosBW2tCBC8bgJJgKa5kfVi2DQq3Gpscgwuwv
WgwsGuJDjwqNookm+VEsQZrR1HWoF82bTqcMCUmWUSzyLgZ10I9uw+UN+kn+H/9sYHNYET9gyp6X
Hej9jMjejeHTCg3QM61dwKgfPxo1EdYINF94ps/2WNJ6TjprSQHBgZOcYM1BZcaPq2ewCnQ/QAr9
w+tswFj39i2H2mHpSg719zgAMmX87Gw4Aisc0FFS3ocNITCzNSvrzHonGV7qeY1qtaPqTDvMyvwK
3fQ3iYN0FoUJPSwUc9UaavbB+wKJERd3jV5pUY6Qze8DMS1ANINPnZLPRrt5BkWszEzlIxhOxEUU
YOwbyW/ldXszxXTjm1GhztXsQMfCiMAjPJkM/b2j583O9fEaHe4k4IJUTPWAHz3jjHM2CowRsusY
GI+BKbuGC+iNjLFDNSXIWMm02tihqYvGhqMxP+CZMtrgvcIvsxnJCuVI9c2pd47d07/qh4HZhKf0
u3eCsbvV4RmQcQZoQXBV0zQW0uCjPj6Rc3y1fg4LBcIxSDkxq21RQwb7vmD5KJye7Q3Rn3U06V1w
BYYET8fhigZZ/Kzmv/fL/T+AHjrqpahtVoeFRbkTCAY2CQt7zAoL7UP8oS+GpW1c9tVUnval4bUI
xz1mC3oCU6wCM6xcb0IBD/+gXrFyyr87TEnnosQ/mODFJBE6ywcM9ndu8vbUgfVkYr9jpSEV/7Np
2hlA3J0DVwr8kxhCjUnmj5eDjqDtsHl0qPYDQkItEwmBx88gbto1B8K5uaG+qeyQ/rEQtdF9WaUy
awN5HVh+qy8bCsGjz/je/M3OaI/dw5UvsnhXO8t45t/zIbvRRMJsJ6NvEJTO0DOAHUPonqg+qp3m
jol7kuAzFerJe5RRmHdMMUmLa7loXWTdtwRkxFqK5G7+Vt+O/6l4PWaiVknk3GH4lro1qrOhw4sZ
ylAlCoeUT3yi5EUm9iaU58fa6I/+J07FfRSoFWNJLcNpTgaduC+M6LrQJs4DJHKO+vgbpxrbsgjN
+ExgxF63tCGG07Vj+E20PQa3VMZtEYj2I9sIKmqmwFihLvzfkaGAQwxq+9RTFXo87Xh4QXFMrHRH
igbpvdluqRGXrXv7/JT95o9N6F2gBqJGfiF6qL3z65j/VeBXMsu0EKGLeOYBxz+GJTMpiPO6t02/
y0Fpyo4k2+JA3Pn5GRwCkgI/VSKuTmF1/0FA3imyNj5+zcQEDtaxvtR8J10q1FnkkFvFudZb0bOk
wTkFH+CB0hrh9xisLKqmXQ3NT0nkLrNRZ0LWgYcI5LOK+caCW2VG8ZpTJPoX5Ev39QQPQrhzilDW
gDWiEetgVI/h4ThuleLAePdFcePMytfmJ1qxLKn9nJNGIn8q2h6KRdI4BiWDs/tqbK+hxJWTkyhr
fnVDFBgjfHhlk1XN733KJOKwLix8xzZRNQdprr5G/3fEtEhxKoDfd07eXOTH/lMKtW7tGO/rCU+v
M7fgXeBB/I4g9ei2HbRobSw0dJBt8raSjkzEVzdzCwZ6K3ai5cYrAzzRvbOIyC3M+rsMvgHDloKZ
5Mhg7zdPGDjZjDhRNPReMerizYvp8QtORpIqrKI7/F9D8jpkzr54TLKLklx7N1o816K36Gw9NC/g
y48xrsYpzBzC/DYwT+Y8Hyu2/qeiGDGlvUXWYQRbgjy3vlSghXl/VuLmD24wCpdwAm/hsXDWtuQI
+/5REUKMkY9QjJA+Rl8mP+QuICulDiRYPc1QYOttMQYUCIIQqfhaNlTmAJF3EI3ttVaODbynEQ9E
lA9RRTDjJIhOm/dq4snlqlDmcQtPBsDGD55ea/F0dn7jcbcmal1lXAnf2OEU4Jt8E4tYyv/VewNA
rQwPlIhBUFaoAc1eCg5GCJhSFgvtSXBnNWobPhvfawrUYVp7AyeAcX8oBtFLiAggOrMYNrJ5GVCj
9VoT+a6FXuUfwdBbw9IixjKLxxPvfpUKSsNq2eL9kDopeWAhJDdTKQ8zHv9r4kwMrQlsSg6D/LKo
rOS9vikw0Ax7yHy5T5wjjZaw6SFxXjY9m165fw32J6sQyh/x02nsr9EQuO89oK7KYxkgpxXl8mF6
F8S28YpZUAFDaBKZUhXVQ810XIBqY7pa4XbdI/tGY2f6f43bfc/7nzCxCDN5Nr9z4b3cIFyjq6Zh
p7ypLxmmbap4Md7oh6nG8DrcKQzn+mVzWn224ZLfI7DsRye8c8zIcX54XrhRRmiNHgMeivS0wxsi
X2yw6ty7Oi2DtfoZb9SP4eTTjVVzC08PKE/DUqoFkgcLs2+q9ema+xXNQ6PcZmjll912/153gyCW
iIXkgrI1TmtppGsuC0yRgfwxZhBiu0SMjvRvAbjR9OKveYUWmbhgY7O/4xML3DayBzQE1dGe+Tj2
zmb9QqH6nr6GxEqMIOmyVg2RiFTNW3B2QrEY3UaiGVQsd7O6r+sf0Bmzz75VwLVp23wVwzeLSkDq
5JCttzCmh5DTGvAgLf6HN93NfCSgxK85o8i1u5nILVGy+1kJ14ttuQJzA/5jkDYEjgUowRokg0sq
QONxeISPLsB9AnpuzsWdTlfFH77KHIOaNDZvT6YlHH24i5hX6RP0yUcIK+AgoBqpfr0vMVpxwLKf
3hqIhESSjtfFlj+CZedihtjugKYHhdbn+MBe2XtglUV6HB4cZrV84Uz3Mk1rwLNobDHqkn0374Ay
4ZWHAueRF9BsIuwaaSnbX9hcqfP5yv0ACEXQsP3T1kKUciwaYdukCnBJr4m2aPr0kYRTwslsPfmw
fGpfRCCGhoFoeR8o1n+Lg74TPVlGYacXnPDv0/39V/4/Q+UlRvUPLQKum372QDzcxKbNX/PNrzb+
zEJvVTPyn4NAZNdNhRTiX/ZVW4/LU+QhR9lI1p8nEnDuu1vWbyqftx163g0ewfVHmUkAOAETdm3T
JsBygs/z2snRUEzDoxaGAX9b7aZ/dqtxWL1DDeioEHE5p3lP3jpV+9XcudnSqtUAAnLSgCBtRR8q
0k83M7zGd2qipSbTvVdU6OeO9MXdhdzi3+1zGRGTVKYOdRWWsBwVAaQb39mDG4p2hdbPZgUvUbzk
HNjvWKH4KL5GPFihHHutgzoFy+slGMTPQoghAcnS01JAvNvgnZlBWvYfuy24zcCf44dR/UirDQO+
dasLFggAeV3PZzdzJYRGeBNUfAYMf8EKqI0GNrNESRL46O080x9IgHL9QoeTU/7rv4Ezsll0xytd
34DKoSvvbx/JeeEkMrDc5qT2Sz0w3/d9kyk5vc5d8QpHTK6a4BkRdaPmNBPAkXIkjYRUMRgL/9d0
RbSomcWZQIZV+Dlte2F+RQtbcgT/6VF5gtOlc51PXAuTvw9WMQn0HVulVG4oCDjjtebE196gFJpg
a2AplcfXrwbXWPvsLUNuWbO1PzR/JiMTRu5nQT6aFnFdKtS23id8fgfl9CS3fTkP97srOgk7CeGI
q3zX3+VRDfx63fHwx54ro+EgOMPMqxeWPxaSrP6td8kmphJ7Y5r0KCx0WFg7QZnPRT6Pe/Hp4bEu
NRTwy0Snscf1VgFbgLEPvaoqNhk8I2LVwuMtaQR5z4BwSv/XbSUqy0fURXs7ERb8SZG29LMe0QrH
sK8xtuIrWRKFRWRfyOG9hRXXlDhQEZzCZ6FAVT/EBE/3Qke53ZipDzTPbWeiHOf56245qZrcOJ9/
wPsI8nM3APtrPGd77yFaulJ+HujQVgRT3oUNBDM3y/xuciuvZM0YMhwTd2LfcL+IzDlPbdFMZ+QO
ID9E02/gx8a2+9UNbK8fJYHqfLMDtR9waMe0zAZ/G8hjVn37yg41ZjLMCqtxvLublRKUJlx+az4N
90KnqsgB7BevZtcUYSK45coIsCl0r5Tg11K1tHcqwKZNZYSLGDc7Le1LRRsrmiQdmLwLz7vdOOI7
U2oc0EblD5ri3mhL5nTJBSFXQAZUAZ9nHYl//xR+833gdTnpG9UovnbHhBGMEWM/SOe02/JZaco3
TCPAlCAACs+bpU2dQXsGlgnOfUCdluq1v7n/FEuOC8K3mzde1f+ToGxoLKy5agsNrNjwlF7qawdL
Q+wJhcJ74eeHu2NlhklYh/ABz1ff9PdUGpq/15+mNU84Eb2klzevVXTb4HH0swSVKwKi6GGtHDaF
EFg0U6IYMbshfhmpj/vFkTkblZBuMmaWmmh7JWt2H9G94F/d/cBcDSO3HQGYb8LxouyL2avu85k+
7AQy+G/H4ErUqN++ONOXpeomB6CJHCFuqMUiiZCsC/IRglU/GqglTA0Q6Nut2NPsjaM88gN1L8N6
whLZzo7xUO7AtbRFHC7uUFhjgkiH0Mp7Zhxs6111X/j2lSw+0UlC1Yrb9RBr4du5njp8hNWaToVR
0ZMOcPUYyuSWesGDEnBcwjUOrmXk99YljP7A7jbGKlZ+5nkonbYkZ34FQMjzjtpdaqGFtg9dJjpJ
bOF66mAtezTfQ09MJ9uzo20J5PoWA1lc5pPeMtJw+tcZbIV3Xi7qGcJEG/RrX1jwhVoEnNgSbduM
RhOZiYFvmvk1dtVPRxUvjBYWJPCbhPQVfRI6yfOkk3St4BQHzccYU1weuwr7/w9VMCOYJxAyN6bV
KwUnV+W8nthOMSaYF5gGyzY1m2mDsmb3+X4M8cTGt/zD82ky0lfWFUvOQNcFUFXUU7XIJGmQfuts
yosl90YTOvi9+sX5nYRlIvXfUcDIq9LIia2oqKy2+hViXJt647dS0ZFaWdbPylfGCL9kQ8trTRil
r/aCinqxnC+iP0sTqGwPmt9U4tzc5p41zzdU9j2Assi/WTChDZB9dYnKYgN3F87E0pdqxWlDKZ1y
2NodVKJi8dBJyK9hU5VKliPozcQcBYFFloSYeoM6STOMJ5Jopdg/x+gH2D2Cdzz+TV5YiKRXUVzj
332tTlCMv8LTJ18zatj0ldT8OD4U4v0pOrmX34c4HGmdvmf4XyF6+6eNr9aIEid+hMkpLe2cJxCh
JOxUBPLUwnc4jxFiInVJxt3fzC245jK7Ihe4+WrWhFo/zyiNFvUN5WN1lbfOQ20RnpFE+rPjOZn5
HivStxdtz8OeN4rwDG1qGMmIa1c7TNpkKzhnA285lf0dOTE9xhsl2jM0mj/JDK92KET/7PhNAXuL
+ILxVK0/6hRyEMc3Ta8vh5SX5SCpdg8py3pnP4/851vQfHiLg2wDuW9LYdjHqUqDYsIvcocjzcTt
z2kmQzNee+9ElE944JRDjLtDkOr0OKGp5zPKUzUYTAVDaWBKo2zRrqFSHzajl5If/ATkPshsYAY1
MKjmvcfW8SzIaIlbsrBwoX4qY/Bq4ne/Lvg0jgIWS7WIbSnkBszjai8Lcg9vs+0aPaCA4foYZVfi
opSCBYwdMr6WUQhVrnqVXizPNkOs8sSbvD31PM2qMLnwraF5ZEaSPMkYx9LY6lz4UqidB44l/UKF
a3b31DK/mey3/tv7RYGar9GOMlKQq/1dd/ze+t5xOiN1mkRGCZoS94SmaTCbvFtPPdiNAYnRJ8iG
cYbSQ3V6o8iWZ16XJVIlhEAjNUDdFLbEzzJ5fcGbGe9oBu0fYYPgtUH24sxd1JmtPe88F6FoKoOs
/oFDQ45gJWahuOiL8XLEuBeSnN7pp2wUoGmGaaO+8rs+vHmaPC3XimJxR0svX9vtMfwy1kUSn6Uw
fxMEl0aadf9dzC1T+45e5PHXsMoEuflOS+GRgG+ouN2uP4VtG3toUZQxHkXUihxAqYAh9btsnC6j
r0s1LzMfcKmBjV7Qmhlf0l+YnppHWy5fE2dwZ9VrwEjQhj3DrrmEApvtPLs4If8lxXhDfRJDFgKI
ZbrGG7wXwep5E0Rld+ff1JQjtdfLtU6lkBOkBRMGHODPHhQRsSscHmXbBAzYCNLZRauVaOfHpGAD
45EQmWpQlEY3jRqjyrXNorST4Yrlp0o8jEzyOTgy8CL5eUWX4jRZgaHDURqyEx4r5sZZz3WfWXLk
AzsPgIreB28t4gE3ZPwZCv/CvJJKLnQT7K/jFkuSKDHfok8Sy+avGBRgWNBXWquZihiZ8x+jZyUX
Ad/YthsWl045js7GPTO8oHjwrUpfEEcoUcYv4A2XdcsJh064QYJn5YQPv6jisAVruhnqH4vwJsuf
diFjOGt5JcvW/SNWdh9S+xH0xhXtX+XQmj7LdDaRyez9/RCKQCFPwMzc1NFaGpEuGqi0rXiPcGGi
84+elxS1Ixureuporu51pzB8YHPfRlDVausnnMBl5mOKKmsBMCQnTr6zq+F9DXfph+namRxzOKo6
0CP0gD0Umt4yVOaPu8RrS0FooUWJFIlhtkN40vEXpPRlWtTN6P/x4sTan+2evHS0U4UtxwpWSEv7
wFLqP3jy2eBZwaJn1E89rcXPBjMiDnw46cbpgRurcp2wJMk7ZFlfRzHG273YeFaA5yf66ze6Ps24
U76jE594GJgmvCdXs9zKAlD/gTJzYjDN983CdkqST1ueBAf25cLq3P0MM4QQPj5Knug25LsCA9Kk
+21Fah/u1QqnBYyhUUPUv/FZYsBkULnoLHmKy7BEpooFwz3k9+iHgnXq13zDJu0/UX5udg0hmzFr
7j/VhBCgQqRHPrBOvDbBnoC50OOm/P1zhNOZ84GAa01mIRl+fpFgAmBXhUGUtzUEcCz5YJg3M7fK
0xgV1ZGaxU+74N5/8i1cnDOHm4EdZdjUgW8QYsZU6nYqqSF01Bjr8POWa3oksayDOfCAlgUGBrtg
W20H0s9T4WWyBIEsw4QYbdbiPHq09MRku8kgGn61mLxI44W5zDpAXDA2eLZu4fU37ygv9kV9GvJU
2tSl+R6Jkndlp6V4BG6MIFgm7R9u4Faz67zEmyDa9c+Xk/SBrJYZu7PPMAVKUBWrIxrGLZl8fBRG
wUST1wuTeUufyUa5KcRpH5jG+oz7fEt2tfY9h0sYbYm98aOLLc0pVNvK6n4wjWdvfoTtwIWJaFpl
LXoDGkf414RgFYHZAZLf8+ohHOpW63hKSAdFX2J9fV8EKHsJfpk6aB9MWnewtQH/6oMZSwH/0pb8
hF3tKB47YZY0q+Vl1KYeVRZzUYCTY2Vf/EZ+GTvPSXc7e6UFU7f7WLdJPTpfhcDA4lk1/0WgqFZO
D5qeIYFdqsyYtQev+nwiGhvdiqfTjlT2j1P2iGsMR2wwBa3ELAHSX9E/KjUQN8+zXQg9nGBjzpuh
dtHH1BdC2hQgxZFlXR/fjQ0h7c1d+kAGqm+U6FSVG1QfymcnATLiECP5o3Zqu4E+rlkkowmMTm+2
xIZmDr1xow8A+GwL8da+MicAVfwEX1yGRGPFVRgv3TpuMrau7ggJ/hOzx6iSzZIKfHs46oLm5X1G
x3pZFpjGjdIUPaJLqw8zlG5gYdGIlrEXKx6hwr+b4xDUjkhFEWtDSgoFih4v9jU93vEyGBZGxAHQ
Ilj97HBi38yOwWNxQUAc/lArfpTZzaJ+MxeJn5aRbPjBDlZRVy/9M1uPbbquc2GT0sJWC3nAhQfJ
7H0vkiRr1vsqOwrSecxhd6ArYSLmL0Zk/ysSkX0eLsJk/aYrqfcJqvXh1Z+E4w342Qd12uTWN+bP
cqRlWHPeEoRUuFeSjF8ba90YJl6JLpHIIijGUIp4NWVR52MJCnNu92bBpNtxSLH8GXB+m+Sf0PkR
35ZwVXMCjpkaXlUR3Xzra4F7j3TVx7FwY1mDuY2UiK7Sq+UJLlME8fIh9ye6zVDmZISLs+NaUjZc
vAIeXvQrsEe7dswI35ay7aewJw9S9YUGUiBPJ1FFj1Qyp19lTS/wtnE7hDCT/dhYXS7sUo+zTn6b
qbxcjxpP3rB28KA/ycHhREc5gC28qtehWSBw2qqyFVFK/I81zTOrG4lrJHX3+jgFbIGpQPrOjWKh
ZXbCP3V2CLQvGV8v7ZhfHMBJT6vfmByGcoog1lHPjfrWDrgIQISqsKWkjzH8gi/t9Pdm4aFHusb0
nSf322UM2RYKnZqZ7fkMdhyLrDArMc3kyj5hv9ldmuTClR6wqyL1jK2DFTsqE7WKiH3ntjKCuMi+
59zQtfkq2RoNEXEo5y23rVCl3LnUeUUitgEuvZjHxYHOye0iHY+WN1E6UBz883+yXzjZSxdUYAha
EdyCIt3/N3I/JShZJMWWtqSseBoljnyKnic3UNZq2Iuky0OKsvywvkGd1Z4KYz84wkI0GNPJLBGk
SsHVwjlLB3N+kAewP1wqdTGUVXJ7u1EI2npn5vXDDs5Mqo5nUPo+bQgOOq1LDei7NPGbPSO2SNNK
+uMCupoWmB3VgvCnueTIQwznQWc6fqyE1LxXK9t8d94UAuAL0qqh/s9RNse5cv3NV/Q3bMJVCaSs
Z/KDjh2g/69PlJonkhfZaHDbVSd2eE/K4P17pXdo1/nh43M8Rdttc254vtM/voPAoTcDSmbJk2zS
VPKAgSDbukhNtFKprOflFapFlBvj+J/s+5/oa8cxg4i60DcDr3cS0jzepBr2AxuY/f+nEs60Irnp
JxJpF/BTBHC5TBiv8io2TPtxn0yNigJLxV0+MKIGehRPQoXUABojhE3VpIs2PV47RyJqycZPEeNf
lJL/Dys4Vf8O7iu3fJAlwl+UDqI+6C27NEek1Yoa4vD14DVqRxwI38PpMKFwLNot/YyVULgrwPXz
vrYfHfAnxS4xPGgCQN2q267JipL2tKLHPv5L+eKBPwl9z1T2JRNEF3C489poQaM3usWqF1HBnRHQ
oMtlu96KgeIuO9Hnzg63Qkz0ToPRp7rYiRIJuRzzB/XToxLxhBzWblG/N9cHyQYjNpolsaOW8/Ry
IElRymfStu/N9Z+aKhQJN9SEMPtdoarp5LJNUssHQ9gmsVq/mFdmRGvpC5bQGKn4hfteLWqPA2RQ
riV+RGR41Xe3wfLJWXTFHXW0TV3dYc7wdY1bOZnVHtJ1qZlql+P89sGl2kV7Iju8+h9hhdRfs79Q
yb+1qV7wwYOoIHuuS1ii3isQHkOJ++VWNA7dht7sl0qLLjpqHAUvRrRpKGBFtC3L37DQs9Z23wOV
pA1aKbMaSTsPaXSY0r3jMJ6klX2fmIibJyBGcNuLpdv1M8i1Qgbgac6o7fhG7+4Tz4iVbaiK3mXb
0+lgmg2lfp8YnGIJD190Vu6SUvB/jfxCuCUTTFXDwlMtBN2qD7XCRQ2kMv3vtmOlVmBkC/qNFJs0
lm9I52twAdQnPBgTtVR69lOeUKSCoOL70U0nJmwEYjLBWkrLKLjySb61llclSOiVgWl1zQXc3ky+
zC9emykGwEgomCt3mQCWUxxyQSyq5w2NbIqUCTJnhCnYAicP89p7DxR6kd6cVbxNrykz4tFH8iiN
4/t8979ee3UxBk4dcY1ywXBOq1NV+Z1drelwfcASzor2afEJj54PYOepu41Lo97JCCj8ZuTjYhUM
wg01NeZayC+BwN6kDdoOFUjizqD0GR/rIG45VSQE9unbEPUcCaZ5PZpzS8tlYEBMdFekKLukRRKi
ROWB0Y/QC+6jpYWGJWXnZBYevstQN5xtdagjYIdtkAx9mdacRuhaWT2pu6ifIKpVb/BI/KND8GVe
Qe4Tr/1iVOGdXoLBsYz16SUYtDAAoxPKSjFBU3r+ngdWhacKwDGTSaFCtzuun/LQp7UhEWk1e1Br
u+C1Xddnq2p27czDFqXF2/AzX+AeDpNbq6/pZb9Ol0c6KDuNfOJ4hWZm6VyelmPR7jaMZOHsm+4z
S1kwlKMFg8uR2FMkx8/dx4z4NS0FjSUZXoHsCg2fPVworv6BA2eGMugFrlb3+MIPXIB6yyyfs3CL
RExht5FBaEVCuSAoh7dsrhDbvea+9EwpBCxqH4203+NaxWqatU/ALVTCMgCHt/Yj9xneorWkHX9x
aX4BqDVx5B4mZsveKUGc+i4MgkfTqyS+E9L/Ydb56anpuhOocQ24vqhWzDFdE8MtHhO/RZwJNHba
an0Xxd2Drmnbv6xncvQkccysoa0lQmmVT9F/YwSKj+uOMPlG+3HR7CP43/IZNcZ/Vp0pY0dGgObV
yVvSnpe8EyXrsO2V5b7oc5p9W6XLbMZG2MmKCaOt+rYW71/3RLLp/961zJ/7q6lWRQ0fPAJdHutz
iITL+zKUfPR8KlFt1YfB/cV9SDKbpl4ox8OGX4Jhj31r9+vTr+PcvjhkLCRWHWK8/X1sZq0VREoL
ie7YqsdbidhzJUpooEkMWtc7grL4WIvhSoLm75AKgwIR/nInlfaxTB5u2HNvjKL3WJ+7PuwJJ556
+9BmjW5fAD6TznOQHs4O5EoidriucpUAjL0co0STacX4zMLouGJA1s4lZvvcqVVyP8BYb5ALIPIy
Ya9z0xD1W5uHYnkYpQQZRn5l8nXzjfD41WlpkjJIe3CUgxJAc/9Ur38EerLBU0UCK27zEgIsujpP
ifH6vFvFH/K+rEpsenvVl0Sa3aZivCxYMr97biaW4R3XMF/gV9YX1EPV9vpjlf+v9lLmjx415ZSf
KX6XS/KnXrjJZ9NVpRkXzNV+33j7mHtrqsNv9HUEHZzVP5zwsLXVExxZKWwdTBrb3PpGVZYES+JD
+OcEFTJRICWIPfkMO7lXiTed4kSNVL0DPqeqhselOBSaZWAVZx1MJZ9+UFaZrv7NIxxihSjWR0B6
6kAhbPaVWLzrqLrgSQzWTRSJLdsDLryK+XewRPYni3HL2HySxcwcFWcs3HyvNWh44eoyTtvhI9Gn
ualWqUChY5oTm1QT1ZPe9UP8iBVLpNSPuJaluRRQsz9ekb39SngzXolBIyKMucNWsLNQWNNuFOM6
Hak50+1Ugbmu25L0AqYSwa37Un9xcwnLCcABl2u5xC7hq2R4Os057RK/HHQFtgEIQ4Zl3zkUMLvo
w9iNtqqngYDGHt7d5SFfVNZQw2Q9e6Ltdc28yeLzJODuMFBwH3gvqDBA0TlgRP2V89Av1VGP0876
IJODmMxjCviY9p0PgkZGjv8YamGMNEcCiFmvou8dpaHlZc/fNfVXqqgcwOHl0oe43oOh4diOwR4N
1CJV79cJtT0RghXF3nZrdes8k6mKH9GBn8hKHs6HCsWqaMCud0JeTz91MDLXwXu5dwvx54dST/hj
hWjCuEC0Pl+ehmqNwumSwB18ABkYZK/AUMgufamCN6PoGoFiIgGQIQIGSfC+Ncp83B4wUjJzxPxv
R0X9BUrzhu97WrgQFcgs8Pg4bEXJbgT/uMEe6WIc9ZMBLXgnbiVi0KdaQQFMvaUq/Vgi85V+VLVq
scabMkJDMYyY8yy/7fP13PGcqA/wbQlJbibREcar7oN91+zt7miAMVLE/HHj++PB3VRfRInrmZCj
4YBpve9f+gz0foaoQgMfDumu8OY39ZS+LIfLeE8DEXTyXpj9bjBfwQTjCet5fhD5tuFbY/hRvr4E
3x2gG5SsmDmDYywrOJnfMNScrMrjY7JIiJvaesA7jDnNDj1onEJrvX3SMOiyxaNRTzjmwUG5kEjk
Q7rYSxW8KTpX+2XrNgPqjUgOKnwx9k520FJ7z7H84qQpBnKJRhDWRWFwSuzMVatwuw2rRkUbt/XD
Amgy29caxpnUH3IyQD0wyuJ9k7NYQ9wHusxJuY6jtk0yFeNWcWf9VB0WdP+yAIiE9eg+w46LRvyj
X2Hf2ycMWqNJXxfqOEJReGAoN0UnVc16q7l3YH3yd/VFExwWXIZzTb3u214ong0xXG86G8v0lZBr
EJwSRK9sk66x4P4m7drngOySQntPNSKfxxvPjsrQ72jaWUxUE3dcOEFAK5Bw0+GPKcIOpEYUD8Qt
ivveKtWrXXallSVKvmeD/9ZAku4pQiVbt3/znJ6VB3uQUS9zFxQhg4eZYbYhj3tW3dE81KO23vop
7YOryDH4eIHrXHBuK8p6+P3QRfs1clN6QR1Ql0eZz6xG4bmhLEZeC5Mf8Bh4DNfgyQxJxlINeLI5
/BoVg65CT5d70DdztkaQjiQMLQY/NZWo3xcWFHlEN5LTiAQS1l0Jgy58oiTM2S3AATUgzYsSolem
4Rw1qima5AWTwyNmdFesBsGrbFcdFJjb2yyLQ/MWT0wBxmnA/AksNNYTljfQJpD3OjK8TmS/XgVl
qj2FEfQtXwBHeQhgLIkfkF8+FtIcFSp3oBN7jbHDATRW1nLuDhg5jhb3ntGNpGXF74YbE+5KPHaQ
g2amn+ahpJyD6KOky1I2xVtwNp4EkYtXHR9EWTfq7qFoMRl7OfxfWeP4/tWoc2cGL6N7ZYQN5wTA
3nyz+allkAwT9Ml6v/iAOyoZw69pHVSlXYkNtvBSwBDMPhT/mw2bawXV5xXJvOhOgPCqw9YSNUk/
Qw8gQaiBodN5yCihSbrTLOaCrHNHtnY5dBh9e4zl9vv9ovLN6eVzN1VxYzO6l4vezkuHfh6v29Ap
3CO/bgKHtSxmeYe++Mr0xTjYNYI8UpwnJ6aeaRtsxkhUdBbWj2UAgWE1CHMm0TircP0RWQcQHvFL
Jkf5gi6XFwYWmw8WRpXQh4MZd41e6N8W3EOhl8i/QLI3ZP/YJSbSO38IhDvgVcU+hc5H1xwd8YPp
4V/YvblZk2yzRS4M505f4l9J3Gd8UHqYaPW912Agzh6x1wE2wm1avF+aOfGP7Cgkp2smdk3UeZ2J
pT5glKkZbdkIigPwouJBKgPOaPQohVVD4grXMQTxDIlI2VDpCqqzWLOUWURvO7tJrde9Z1Z4bmTg
BqvW1vRIecFJIUS0hKukmybwvmMlPRUgjFCDGY1YtIYGrPQi0yg5/iRng3eDqLYDzCWu26pA/Oj0
zIK4BjBuMLkDBd3CYp1x09EjObNrL48Vb07LKJU/J2u9ZobwX/X5dzSj34iSC6tF3+QvbjUXC9Ic
o5lc3elPfzE+5ZaQDNFjbtqb2ZM96lI/MR+ZN78CvICFz9YmAyuJtwcdNUNgSPaVnjXBytXPrwd1
otH8EhuYRZtIl9sIb1jmJCftwCREBt0jL9tkt1WGP08//lWQFLN5qEMwc5fc5/doocYanOvzTjGN
Td1bXO0UM2Jr8dSDZyabJKe2dfq8v5xTffoyFDAJP2qzzHv8gW5OK/MhJlSYFm1AEpxKLRkT0SNk
3O8hRcs05IVfJASpVesfSQ69svcRj5xbjgCqyBUxflZHQnC4dCxt43JmccorDmFhStIPe8bklpjq
nI/sAgXY4V194b4B29xFQmZs5no0aIZUchQvHNnOlWsRVAQ845abjWqIEGYPWWnz9OH1UM1tGszB
zasdBvUfJIAKUOR57zHIa4MkUC9Cy39x+Chv/oy0ircddvnaSDOrmbwHAwKf1iV174dF8VTwrujR
aDBK6535+4DM2iNxd9eaWmrVSYrqHvQnBVt7YJUbhx74SVe6ocZ15PZExJrhxbBDMhdZCq6DtVh1
S0cjAzi1PSo1aR4p2D/j849gjC5YnEpr3UEQtsxJFirtMOLuss6Xjwh5Lig3n0HRUP5LYTQwFnZy
dQvQPi4e9+8DEuWxoKEtU+4gzeeIzz+If7osGmOBfUbUmn1ciuWcIn0tX1aRpEvunmbFUtcMdv4x
bBqjFQDjzWnAy3IJF/Ho479uMVRLAI13ObZESpW7te/e/ZZgNqtieKBcMBB7M4nN1GCbJBNOdd01
abdI1g/C3UQekWdKbAvpzS73e0+u8qkacO9IugGXFxywaOXSZ3xZHoaL1bK/3QgWdF/mLZKom8R3
aymGLlt1Xky+k6PAvHR8pdONhg7kEY8mG/VISkcwqiSrR7SZVFy2Zw2HKPqxpBOwheZrJoboHlS5
mmAHcLXqJexb8PmsLItyrZ6PSnkilT8zx9rnKf6+83j73Z7yX9aoZuoc8O5Cd5QraRquLqpsQkST
Spr/e8MLkhVWt8nOS08alYrtY8nsgxGN522hyazwIi4cRlKkJnC0O1ASPWFWbKXS4T3Lu3VHVjp2
NnM2nk/DeOTCivwblmPS6EVVf0IbaCS9j+UPp3M2pjtWUZNW+f1tKxXpHfnsOAC12S3qIbHIPfwQ
VESfwVF0ziCg7YT734wrKJqXAZyi9bthI8w7Ofk4t3/gVEWe2p8vxbmd66OPj6Mt1Dm+1RkbumcO
DahCHl7YZZSjLD6zuMTQkpwKfbibZeU+pvsLXfFK8S4DbJUPn2O/eHyC91AxiEJVxgzJJW0QEFXJ
Zzp+/uuhIS3j1lB3bcDAPS+UhuzQ6RGN+A6FQiGJNtGHFTaZFY4HVQHdAaA+1rYr2uY8s9nE1HHo
RXfWJYZznyEljFA8HzCIUcuMHMRpml4RHCdwF5t+9KVFifaZEIL6fKWTxvcwrcCzqD0svYRgC8tA
Nul7Ikm4m42vnVvD2aVAty4NZDTQ0np2Zr05l3xTJ+HI+jEKSu5mlz0541gxw0yDfZRbMrzs5rbg
OFS1Fdpx//YJuLGUn5pvKKpa5TKP8s/qwsQ8C04dg+05IqsS1ArPsFWjgbAEY1Wg2wNyBdWZz6rC
MqUVVqFg1UmUcoU7mIyLmxwnlZ47P+R9z82Mszn8LPKoLTc4RbrkIY6sdzOB3/5V29Yk4l0N488B
MuS9hHKe5Z49dq05C0ccJ7tT7zM0NqsxsLt7mXvaQ6zA1DGb/fNLCaQH2crzFvXuFcdJoRCSjqbz
B9+bKYI7YevFREvi7TPKxTUmGg9bEfNX/j3AgSJoeHLyfXyXySaJgaWSLxA+QnNKTinZW9DAZ6mU
UB2OvRBz5HTm1mBW5w37SNz2Y3ioSXHfpAn9g0CexP4jWO76vThDCa/WiDe0RcY6XHTmfvoJAbI/
ShLatdH2pVW0r4yW83GLzQLNobCrACV/WOpOUxv+xvKHkZUkfoKuorzyrFJz8Ynak35oNOATOOvD
2J+bP4qnHsq6gArvTGFSDCx08YufN+v2/Z9xzN6IAxIBrVmU9zNz6i01tPRVOpu0XO3lXJgUI8MO
W6DmF0oX2ro1SMmcMMqKj2ogJFP+KqpNTDvF6K9TMF9zwjCZnPExYdc+U9td3PnHSmSIQU1UOk2s
4h96ew6IpNbRC384lT+SHOgFhZBslG6mOS7Nu0XsI1YujsL6G5kSQVTpJIpUPHNcx3n46j6BjU05
qvO0RoVWZUuTDazVEHVH9MI1nSF8QDGxVsLUt8dABtZnEdlP3nC77i0Xg/8n/+yeWjTboyuDQss2
/ToUMyxbwXgiZM4pp/516JHMb//URcPUJ1MvYipyxU8Zz1dUAL0D5F/yAablxvmwdGmIUU4bnNX2
uaJPBmF4RVl+3WLFezWfxl+1KnRXVqtCWeSKNBei08efpm7XtRWvnNomFjWFZbH4Zx8Okf0yoYOi
lgJl61fJrkIlYuKAg7XVqZ7kgTTWdxxZ40/fWN8RmZ7Ke9OVTfRV3ysdHnkHmf8sJ5DOyECfHQHt
ynfWxoSXN79jNbc9XnhqC/KDLJFkFDlVvfNA82XaHmqxnLRDP3NFzkb/D97stVIKFRZdNoO9r1Cf
uidcgyyDV7Vzijkt/YMPHUDLGsgDhwb7Yy0sTQDfhxIPl7f51Yjz6MsDIg4Xo6pZbHGyVo5ympup
YkKWIz/oyjwwRJu+E2BkHrJaaZQM67CHZYeZ4igcPTD0Y/mFIhxFPkH7HDoF3V/q7fReLA8qKADb
qZb3AbKK0AJr15vj0UPQQ3Po5caLC5PcWjK+Ftdjdsx+K6mFWL6ClUaUemJV+wyODwagRhcfSusM
MJuVSirFRaXfg+4RDc1B8TMhGh08d4E/4l7TfhLiwc0tH4125bJ22t1IJHiKasBu8UhsR9w/XrR+
Y59j8QWbMy3BsrGrvSGZdxIYH/LfW9anz91Bos4SOS/3mkjvAapKc0XKRcst+uIiubv8Gd0xADd/
0izIYsq48A3q0FoGg+zCR67K+lweHkquKtvwFjJ1ixSImwEjrD8DrbId7G8wfozMxux5YaatywZ5
FOA8qi+EPv8Jnuc/oBOUhir1lYnkQ6u6t1Ut9iXfaWzntKZBPq6NIXrCrGcaDtoIIPiK3Jw2FYOc
q3uvhjYa2w7rvltzPtCk0KaW6BJ4veeZIJWDC3De3ImmsO2C77m7h5MyvaRlctnXd45dnEeSTHLc
yAdoBl2Bnmg904AMWnvrqihzAvdVj/T4ITZjHuDWY10JhWDbtlj/9HLtgtSFguCXTV/2F9/h3RMp
Ap+GbwuRMizWH2W4wrx8j6K+1wAG7QGaqTQO4d6+CTteit/0/vpNLaPWO93d3Fs0R4/JLSRbzS8q
c+HldzK2ikR1tXL1JeDMW3lEepEvnlC8n8DWWUloB8pugSzPh84iE2dGaoi2qfOMLLMLAOdEa6+i
5i5pJ6BiQiNQIIYljVIxtpeTRI68NLpoD3nlHph4N5DppGIO9BZb604kguFhpPZ3WWz7j6KsdHvk
H9mcXrQxb4KJmvfRlcvqAFdDPlQ8rQml/bkAdYnU4IOL8GTdzJMmiIwT6P71/NiTi/g2Ybsx9Vu8
rHqMKvZ8g++kWnxu7YUEw7J+6ibuoXwgojgmVifnYLX7wBniEVQAOu4Q73ZzhJmpF5fCG1euwxUB
KEphVf/OK1zTo43gciCTRs/idalgz4SarVWCbDVAwXve6LyeNun0RUBHhUdgJhBGF9nkrFcDlWAs
GsrJuykXYpQBMKsNFEqM+bcvTfMVxsDsPazjN6ELXHJrbisKO/C3YAWZAsMQw3SVAkFAnRwDgxzE
wpg5I3iBBu5LPOulqGExNg2rvBrERKNDddMLtusd5Ro+VTJCc4HLbVC5qOrDKU+JK+qjfpc4BCGS
r8kPXvDLcQi/JV4jwP2dKPVHBZPEbRhH5QvAwibF1puTC6cP+dhVKql++NVAg3b3nlR8i41WIPHc
MbjDHONlk8NNO3W53AYXZbKvwiAx8vFrG3nfhc/2fzbAS/xpW+0c3MOZGwWEuigAucBtBibrW5Ew
JunandSbIOeOM5c2PTKakXIGa2LAGgeLE1O/KDdrLvorxFaI45uT4KeXY7AVQygQL+EKB5YGzrqS
CQNhOAmj1/3uVk3IIwP+VfDl7T4QuSShXukNUOvgt/2LYgUAaQckCO3YlMPa1LCcNf3fO+B38Yag
3UjD56WGq8F96xenNqSFv7L/AQZXtZftADTzvkHv9r3fsxM0u3HDkJyFU/L3qCN7juP3AcOc4v1I
51lqY54tBwOP/WG3CzLf0lJzuXYzBaYgQgtSAlWfxiYdNbSryE5Q2wpRB5o1mV0VdYLrTUzlkfse
Um4vsfbBtBWKoawDPRIYdM2FWErHVTo7EV1fVUJqoh5IjkzsdGsHLWIhnfjWfdkunUjvaoInpc15
lSxu7Nt9zBlB67+IQvKpFVddR8XaijY+gsChD0xMNoJ7p6P6oEtd4C2vKLr3VF61kVMoVU96fJxV
8NskhlvVEkTh8tvoJtElV+veuAekraBP21rsA8BG8keGWChZxWmQ/tM6vFCpTS3g8XYJ1xPC/XZP
LoX0mA2V52JVmQ09rFyC1MwRJfOfUbtBMQdsfVugwH4Hm4T1PVFPSF9F+bYWCnPN5qYq5f82+SJt
/TztrD0NL998LkuOTsoFaKRLQBq/5hrNGjSkrGN9acKGH+irTqvePDLGWLOU5O+MkyGqFrlVZDpt
vlTapJsIbvpGyRemh5f7lcC+W3NrOxOjz9wLDVsbLF/kMj2atGA3HAi8Lld1IqDUXG59s/plcw5e
mWvJqpJCIw21jmtcMenpGnsPVuLiR45b8XEgDcTcAoWBr96UO++Rehaa3jgMisu/dUlNDCzKAuRg
b/38wxEwMdQ+51fuYAZKwvU0LZH/Kuc/bG9k5ERVHlF0etdb7x9cq9pl1tpo8Q3Yex0H0LWVZus9
heOvo2gDcFX1MzYnWa8f05sGj+8uToIGKSYXsTGsewMg+AP8Dr2NnK8dez2Lvf6I9L+/x1/558Be
MKUr1JlazvEo6g6KauoEUEjIIP15WgTzmNNDf0DPbu26anwecR4c4LpgZFQIT+uUmFp9mO1f6guq
US1h4UaNh7Zl52JdVbxqpM5aNyk/SN58tNu788HWkLf/Cxr5zl39RCx/DyYuJyLQr1/Gy0JD0UZK
T18h6qkYRBLj2suciyudADSw7rvkpbTfC9Y/MGprmLBK8wbDqCRdmfvA2T/Whe7aLqKkKJ+K4F6G
yvlHFziwka631oaBUlYLp+GiEqwe1pZBDbRiDpceOtBuhPwbyRQwGgfhL5nF1CuU8FRvD7pmYhFu
BCTbQKosEsz+tac0ENsU+PyfTixez2Y33Ae0nN4MLUBNeengN0p2STGD4nyMMdqxJjjo0T4gRjHZ
z1hpbbMOSpjeJAkCvEH+nQGRud2q/OH0fAdM1lYxu8tiWhb5wW31u+XKU8dkhb7fzatja+gBwpHI
Mp+ZadM3onp0mC/Qf/7n0M0B4/eazJbQvelURMu8AHKCp31qsDWY7At5+1mkPMKPfFMnTE3FjCEP
3j1fPjeHUB3oltwUTayAfCF9Ul8iLLhpYiNGWc51iOTN22xkzCj3fTPKPU7in6dmtqAV+a4XaT4y
Id19T44ZcJIRaRihHwwhxHmupC0xrg0WmguWMKEVeDnvm+i4LQjaIMp1RYLdvceQA/20ku3Tt8sj
6sA32kZncBzqld+/pcs79uWrN+25RtsLjeZZpbywq/uGc+5zUUoidj1M3ISALzqXayPHi78t0oLa
lSLzRvKF47xRQPIKI2LBpOvRTmbugnY+R4ViUxgBp1w+P7kDaD+R/JcfYh7MzR5m7rl3A+gU5u3T
1yveFs0KebmK3eMNwEbfSyIt7AYuZsNf2p9EWHdFeAQqG6FrrEW/yU+oa1UcBvoWA8TkGXmiMPhx
JoApkwrM0489Xni7iZ7syg82MwrDw0XP+gjEDhjodUrVtq/TP+Ohg6qsazw138BIkQsLjJAIvg3f
WzFt1OMLcd+WAdU2JUMs4XTmrRzghnl3MvJCw2MsuqgAXhGz5nsHNgSGu8Ea7PbP4IY/TywRnkGo
2IBgHFHDjGZERTg8a0wtnrpCqfBKS+XBFSj17gyHciSplsEsKZ9nxEKumeelz5aLk57ZECaQ1Nb0
Rg/ifDA+L9XkC2NWR6dTbXb4lbaM0z1AwmCCBz+lLKPsMZhpV9sa5PC0+8REHX8fNfZIG42hP1ma
5kdR9iJXCSPiGS42zICk9+Nx1ZY0vWT9bV41Tsg78jDOBV+86enVZ1Ei6Z2hYVd2atrBIgX3NZtx
mU+PptSU5Bpzegpg0ctIzcn9MpF4v6zxLdX5prJvzhZbw1sxlWNXGaD3wlEve6TqorWKxnJZp0To
gWAL6gswAa1UHhriJ6l3ZlzQZQM8bRokm3jpGir9ZZmgANUFQQWQTW/4qbVeLpGEQD6cNsz4fmai
NP3/ebloLFgLj3iETJfo9IEqXPUq8L4Irb/ZZ0/OhelrZYQjdcDo5J1bA+wxgUuVbp3nn8jsDjs5
nFgp7avQWoGilXseEYfk+tLGpZLSsfptqgBxhCjFtRSWNz03S96nvLwsmgitxMIbmNy8wWeR2B56
8K50JMM6CHPx6wTTK9QxBtw3UAqGCzVOYAdtVTaEGutPCfzTVPEBXiF/QNDLuwFpKOVlG0l9aE3U
UECT8+nRreS9zQ3FfaPeJPA4rbPr54fRpk/RS67lCRfkBuA6CTDtKVDitP4QNCMZFGEVGICMRIN0
ZnwsJJdBO7Hv2lGlvIq9WM324vdXdxbyjGdtRnljuT++lFwd8E05Bs20eWi/hxxVTkJA2v3h0txd
ww7v/aks0iTFAshKL08vf5Mjod2QSNey0VpiPHMBxgQUNflxmKnax67MSD7Z5GFaGiX7YDn7qslB
6NOnbNmqBgBSQ+PJbFq1Std2y03BhlAtA+3VAfkFcbCNMGxWyt3MlgmVdyfUNwoV+nvatMu4zq5y
Zb7LP9euHnX9ADUh3d3p8I+xzOuev+p6Viw5OxV+AiZKL5dJzNUXbCS9Yz36iEtfvmOku86jX0+4
QBHw6zH9zOI9+zARllfrx/WtgsD6f8VMDj9lIUDB8YwCj8S93b+DWbbEtZdziXZhw0f4uL4TUTl8
AwfBJGOQfBWLOK+dnbHyaLMgTqnJlEtEp4X83wR97egyLlvykW0jrRuD1PJ1PIZuMwx07HRuM994
5bMPbOOIFXq9FIqKJAI8s6iExSu+CRedhwVLDL1CYBwign0uHU9+kze3UlCUKWo87uZD2YjK9viT
FfAWItYG1T/f59+de84qkH9KijFWcFIqFMRH/jrjoK/h34u9/FzW2AK7gSerWw61/Mxp/8xlSge0
PPA54WhlVKSxqjt7rgOWosmYY/r/IUv6ujEyr/MqyaCDjTp70SN9cU+ZAM0TmY91LZflrhJBA7X2
kxZcASZ9gUCndDvJgHJpJ2UJXhhGyVeJeeNJZsEaxNg/w70edROWkQw9a68Gav8M+C4w7jdWfgNw
zK1bBRSnXvzTiA+Hr9r83QSjptb+blkjFoig7WB9O6KLvJLkZhJXCxxGk3jzK7QtIE6qrh3RJo65
hDho0gTerpryziPHtehjJDZhc18lxK0j1mLOgefl1urTxLXP0XbsaRIP3tSZNXDJQiRY7G7fKLKe
4DzHH+kJxBelf8xVYC8iP8Eduv+vitKNE5TwiS33XhxBsDOgCWW4LF6pqhdaq21i7oJC5L0l/NC+
FyDHtOiOsmrP4uAIsRvjaDifnFR8Y5qkzZtkTTPt/6Q0tCg2FMV5cq9nIh3Suwd4Fw2FHLb+NLrE
oq1y4LmLZUnyImfNn5qbDTO86Ai5X9jE2auNoEvoiJjpg4rKSCvtLHWViWXRIWi/Gh0gmADX2U/6
QOGi6h/Mf92KwylY0+D7G4ZWo4LkbEFFA4z8fj462o177teGPi2Kl0byHettK7ad4Ag3o2Da7Q/L
qlsdTPz+ucd44GDwJBg50w6CBufknjHb2cSyaj4dl0sYU53ze4ywKFNoviBkuPBzF8oORl36nGC2
HByi9oBWrsvJGXZ7nlsv6yYGoY5C5Y60/EzE42X+hFwdJCr6R14SW4tct3gUyUy8lZbRnM9oczcn
VYpd+vhGX7HhWQqp8FhJ3tPqREBlK7MsXIjSwu+21bzFQcp4dUf/puwBxjCdoFHoXJp7B82PmyC0
Nh2eBPkNJVzU+HxiviAv43wmxLIeiOb6l8wiJmpLDVxNxN26cjNHbgeYwxahJvGqCxh/Wel2LfvM
T8ELxZA7/WlUT+SjpUM3Vc0pNGV3fa7eFy8R2eCrYKkv/oShDIJlTQsgH7YOt1l+oQuD3Rsa4TaQ
RsMNtZOy263HH5oEWM94z868dMgFrr6KAg31kfyoVuofZwQ3MQRfdwpkk8E87CtNYY60XHy3Y+bJ
qOGognnp/Zs9AukMzfCII1+skHDuSF52ATNv6smjbYevyDPl+P6qD5Enm985/COHLMR9s+Otb+Ug
HMP86kkXBugF/IKBm3MFxV28RNfQu3K+q3rhOX+jdHpjppHhmTvZ25DgGDJxFkf9m+M9zhwLmM5c
D2mn9ojanx5raul0E21X650tR06EqoDfcZk5TPOfKIYsqCrKvkRwxVlhUzd/13sJQGHM7UvR/0yG
f3zO93lWrBVOdmfaQx8wcofkvl7Bb4Y6bX3Rg+rgnzg2wq+2YkGZOONjtKARq+s2U+yOyn9vQxQe
g3y6asxmdVrWsBDSpPEUGL9kNN0XEp3K2y8eoXTnI6sQvqTUZcHKBhWVI/dxdBsgY1jGb269hCJX
9URwmEPYi5qjaaTXtsdKAMwNiF2DUc8xmdIwaRwLkWfsX+O9HyuG75DAFe0rlBIYWzt2agxxCPlK
JxpWca82wyh5u6zDpGUmI+/iUDkhjblRj2hRmT/OKjD25q8sG7KhODwVPmIhYFstHcy2XOR8oP6m
MMnyUkTCWWEnfxDJ+uTMUkXbR+bIWkiJIM6Dg07cdIfJpSInQ9eRkup/n7XR29t1qCNtkS+T+G3s
LMsq8dXUjhamv3B49S/uW6n5pm5PHbKdkWRLujeRze8K+otZ4U/75pTHrclOCbNLl9JO+P/eJ8ET
aXgvTypGRKHMlJEbgfdm0fzRT2b0LNl+Naw97sh/gJ7r3VcsE0Ly4GfcX1WqkI+jq9EkA25blPTH
IKhfSXb6FXupo9BkUMnZ5IGPzNLEDnSS+IYe0c0nJ22L3mjIywFHZEgh9TOj3kCG6KPboGMQwS2y
c8wY0V/3zQHNCt61pgGLB/2oHP9Fs3O6Sq1IVC5dfZEJDMgsoIMBHDyITanpHpZZp9Nx6UfvSByQ
xAB3lEN8Vu6npbK9UY55n7Pyz1rAZKbCdOsn6Q/P974wyH+Zt5ileXUr213glP0ydPrwmvHWJ8rU
wgw+6+jnWWuy+P1VuKgN2H26YUKiHproKcFBSeJ/lulfjRNRXVqMP5nwnMppdF/4hinFHp5j4yDZ
3PD5c/dRdi0ndzFAuZEUPuGpv4Tjdwr83MyNwcG25nYBNTAQvpBkYweBp5zhXhpDet8b4yeg2wpr
c0GlbbHnw3ZrQuwbs8nPynQMWLddcQYv2NYkRLPeFvjzjoxKbeMdQtgajCbsALGTXv7WKZYG6OfS
OMv7SxniplhA0v7CqwvW+CkjDQ9aMiPRLB11lWHt1cw0zfgHx9d0F8xCHUikP27Tz1HACOYV2JG0
fAWAUqxPnnTHbPA6kfOdYYKQcNEKrIrfXbPrwIm6wSv6y1d2fUnPahMAFKivacKidiZd0YrxDG5D
UPFCMq21BtduygDfoSlqXSlpVq/pUY1kTLdGuI0ZBNVaJG4UzC9DK5jwJnSshZfjnWZgGq2mB3EX
lVcdBkrNyUSVyoWzZ5PtyUH7ROs6xmnjVCVZ/y5vTlsa91lt+6ID5CxtYYS6F1t5+dndtaGqLule
zbY6fG0s++lyTrNI2o6hcXW6Q3E2YhShux9nSIhAJcK3qg+t+Lg3MUDGmAjCNFWu68BiCKzYdGxd
oxT1uN9izPzRygi6CxwInpCr+FqbCqwG3aE3HPu83QZcFpXgDHK4fj3hDdf9lM5oBowdSxVXKRa+
f8Q+Y9kTM9meUVZ9zBKaj4Oh5Gmz2B/fFdTFtdpXfy450kiWixgY9GtzKUX9yyrqFl5rjX0NNOXo
Gf3LSL8BVIQa4ALHw1oDe8A2c5/EJRAq0CYehz+CuvUBWtYPMFgdKMfgodgBhIfWDbBkrkMKywku
MabF1sThi90dfccB19/eTm/XukCxm2bz5wzaOqD+ZmoJMh9Ng1/Q25b0tR5m9+vAwqMsNXVYS9xA
k9C8Nz0+NCGSxi0E9INgPvKn4fC3Y29+/bHgzFeeIEyweujOvdx0TX0zB5e73oIXoYjJE217LiaH
6UePsnrfABtgeMgc87w/lxPicY1mFWqlW2COIh1LtSl3tNMPwPduaMjZdoC/e9sAjnhQH4AIUHR9
GnVMAVvlHyJiM3rDOib/YKd6R/efYlUehVDvXsP9oKCzacZo7amqAMJKFAQZcO5Bq8GSE0+CBKCW
aKp4DITPAuE9tcE3J7jhURBgAGTrIG190qkiSWggVlS7AxYqkTT4fSM2NAGrKIVkbUEYV6enBuUK
/BJlPU4KVwJ8pHalJ/Lks9SJXFSjJmDL0nhkRGTNRladrEU/JIqVF7HVWM09J+HC3pc7e9BZ8F+v
Q991IKLia2xk0xz+/RcxHvPtEqe7CLRNJrw4Zhoj0EmFetbZedTmMYB4GXP9ITsqNVb0KMEev5ZB
5idUPhGkC9/qj/EKYn5OHigN9maJHiXdBDtVT1WOKYSFkAnnpCWv4rdmMdi9ZEKk3PTESB+jbSzg
eQs9XrWZrFIU/yBeqGcJICPspRWCyfudma0QGaxEGLzsBCwU2xiVXVw27q3BiM1CagBQWfPMf+3K
IYNL0IHuxplmsM7lFbrVmo105Z8TDQ+Ofw8qzczvVwNxB3Es05lOROZTU5085IIyppSP6otuXX7X
XBBO1ISHQQIlzP9YFgfgvsmzjfhrkvtTk+7i5x3BUc52huSsF/Ybq+Uce9PSAfvhpVM0Y/XiF4Cm
P7u/mnS1wdDyCfruWVVNqIO/sqdffOJz8ZfqbxDOgdUZyUY0f5g05OzleD62RsSRsLJFlXpO0ErZ
DO2OSwnxraVXfW4ssKO9MYDbos943UUfLzVjCyVZYudA0ppY4RU+/hQd4YAGzr0u62krXGrmbS9Y
OsX6H4pjIKn3g6z/rOoazLA9k6teoraY4I7KlEch8sfOcFZLb9DxpNKnT4TElPU/C09mGzUv7qQi
AZb0DpA1GHEunMjPY5JGQJ6Sdhrml7tGShYcFen3naxOqMv297UEqhL1yTp4fXghdZ2HK/XUj0qM
hoOz1r5ZgoU0DSEDB4z3knnHpPBK8p5LtR0T/U3JjnK9uWVh5km1ARowtEt/4qL5/Y2B+cZhnidl
rv0Iv+shMDw1fhehvAFZz+2QBfiFlVZ3rH8bkYlv35lrkeIdhnpfUsHherRlgOlwrgyA9RKMbp/N
t9YJlHU+ILzLWPL9VAxJQ+4orHMQ2FZEM44RxdeGKkfn4SDwTZc/Weah3dIcE0JmZflnZU1ZUnt+
2ZctvIVpSXkdr/GLbTqaezfSoudvJKsJdjQJm62SQGJulN42SyXk35icWyl1XWHO9++u0/qYlQSe
ElUobbVpL3fqsoHhqzGEyEcDwGdnlL1UFkxnAsp6V0betmQ+D9OqheBuFniB2yDmtwfWsR1827hR
1+O/mvY3g05I9mcVrqrggkbsbwYZDgYPwkUpYcEkWZbtVANe1ccLNmbzlNZnZjrkPaWwL8w50ixs
iFTq4In0pHYCdssqLnkcRaoOtNfhD3wBJKx576Vfqwr49aqLk9aqGtkDx3JeIRt+KK0sVoLqDWZG
O65ztjFS3mW0RdE5gGCc9cFK3dfeZuaQKzgyMUstapRUlOdts21gd0XXajs9z5FErAfGbWhQYxme
tJ39EmjWskma8x+lYuXA/8J6pm18AqcncIk6OKZ2U3uUEDN+keM9w1K2/YdV6RATiX+yG/sg6BBi
YKA4Z6WP9E44zP7FsSQGkW6Kj1PcQFdT8q9JMj6KeUDQ0utoNHQkpdUM+l5b14WCPlViZuFrX0/U
7w5eVLn5EYWECOcaCaCNIx6f+s+r4bnngIvILUdZzTOYGD9LyZw5eWbvvlXakbtulq7WZbAoIZd3
vquU1XXdqrWV+MsarcmyMzliOi4P2Eo1+QE3hmpuFP3vC2dltEwJi8+kzVExtnqOzS4bUUQU21bJ
ouAazylOffpUbHpwUw77v72iTbMsAws7J2oKMxprLGMFR3+k/Yh6SFZXLGqcs/HIyNxg5bCQfmSb
rcMQZmdE4QUeAjZCRY9kykhcV9YWHVaAQm/o/k7IxUQJtz5ubxxzD6pYdRpTF+pF1b9yd6sgxpqV
jKyerCbp0Nwr7ex+dML41DbW+9IZ2slot1TZp6OQ2JhJGnFATQqDlDjUPL38G4BdbGP7rR17dAVD
8zQyAWhIcJIloLBd3B5VVM2dnG/oFV2wcKunwOQtCcLFAx+Qcyrhxd4PU1XZHwht/yZt2hiMbzkM
d3Kn30ztS+wiBvOIg8FwqvPiwWupGKdKDnj1is6Vxtc4rwxs6AffJYVn9uvZsl9t8A21QM3/4QH1
uQHmS1zr1hbNSEkESu0R3k/D9aToPeHneQcp8rO6LXuDKxeap1FnUs1E9SR+PTH0z+mVwujhXfVG
CD5UKjGiSRHyr+v3MrLue3zD+W1WZEnGzPWgGO/rL8p5R/N/GOx8DU7athAvzM/rQmXdwurnIaTx
BAOp25A9mj9BQbdMdyWEAib19H3FOH56uhGpAsak1Tk+b3dxQMRCY3sucXfv8BBHNzxtSITHub4j
zM+mU3sJx0asYKCm47U3+ZK0+IjshGI1bXlHaSvJJwdbN5y5OLHDRUp///eK0IvGXRynE0qa/TKP
KHbkV6sqTFjaj4C5OitLD31cXHKZa/BFD2D9q+eU4Kt6q/PtpZ6rVdSo6nOYHYTGmMRcMkxcGdNr
swWuKH1nbrafZoN72uFtA9R2zYz+Mz/QkzGXDCMF+iW5RvtnZhcTWF24eUhPKw+I7UFvsmRVQ1IY
HtXXO3qjpFtUVp2+2ekfLxpAQ0uaZJ5BbuIZO2+UT7dumLuSNji+jg0ydGVEnTelPWgY3+SAXza3
SzJHtFU/4C79a1otwtV/2+03J+ZFkbAT8/v3WNxHGQTKFoL5/qXEHUyJWCXeA9Vg0UD+vdItOuNT
W0WqcB0H4G468EeSdoeXnrUxdUCJbEBbmjWb+ErtG5nClIl0WvlAfhSpMTEj3xbi/zLR4TTD7cyn
WfhjHWI+fDEnccb2/ZxZ+HJdfs2PauW73Ly4dZvr0fC0V36PQcZVKum0CMi1a4oafqrwiItJTdeB
BcYfK8FWSKZfOJirE7rZWF4zpNF9NGzArQHtflmf8O6ZFijWgXpsu4R05EZhvFbJEVxgcgKhUMuG
4st+eZW9N2cWu5n5GoWJMmGUiGgWVjP2pCoNS7uREPzm/I2NhOfXvpQr3GVB8vfyA2Q1LzfiBpmt
Dtzz5uBOwVcA29xgbsWEbW1pdsFDTgBTuFm16LybkBJWQ/Z9oD2d3D3y7ZJIEz3yrXy/p4wzSWtw
FJ8HBOYwXSlch6ZA9p+7ZiQ7ekGpn90/itLrwDIwIyJ9uLg0BjI7GIkeNu9AuEZYYfADiwKWlehA
f4R19oaUbVCu+XYf7RYoJA5vNVBuZBJ7Y8hM9uOAw//o9LylvXcw2bNlgoJquchCzSMmcX5OAUpZ
nE+lqX1LkIudoyyaIiIh4rwKHRCPQdGv2VZYHUwgko/99hQ/qGsDnCFXi3SDBGwXQMaCHlPqe1uU
NvW2OveDKb5Opr7Qu8Ct1n+CYZsWtIp8vLiATHXxzEKQZhAuNOxqxKh9d6NBnsM1eua7exQ7Z42O
6SNSl3H2qM1DuytbSBpGqP35FW+TKDkX2jJmPni0z3V3OmYgb3Xo2L/0mt6wyQQXRutLwqiLSvtg
/2EMBtqR8LIowTeaYDytxi2iAUUmZLhbxTVpiyQCLNkDboCbG8JZ4/dheqKePEXQiaMgUo+1x+zZ
B3HP/pk7JexkEQ0InnOqkvzEzvyUo19YXPgygQpCkfychp9t4Eh59eWccnbXu3SrOTG1IsrVJZXs
rCCuTtaiV5617GOOLFvQhrS6ZudiqUh7eN58oCRRiUa6f/aqGY5qlGLb9VtENOXLpIRSAV2Yql9p
hVVBEIx4emfy8e63c26pf+klQhRzXQNma7QI0Rj7W1Y+mYniqo9LWWinqrk8ObHbal1uRkRc5l+1
YGyal1bfnqPC0zX1wZTkU5faB+cCHWaOUZwab1OWKWUchWa/1Up4EedPhzofvmsjf/h3QmGNDDDP
JhM4Afh396JSDpRxjOZTCtGLu7pUu+siHJ/BMmW4ny2/icTbRQB0yt8IY7lrTt0vBus4DvVy4pm2
XJHHDqrQvDTJTbkK4UQbSIzK3mJxJcv3J0U6TK5wxB9l694hMi8cd2PP0sj5M8lq5SM0e8wAVEzN
53IOEAW9AMwBkyubjTSNUZe4MJb+6uYogjmy8pMFPdoiNvkT9BCRk9dUKfIwehOZKFtovMVTJk++
hjhA7iItq7FKINwTSVbdOB3xu0q/OxoBWEkoiY4KqEDvpBwHqvHATcmoa5drZPRudwavYG3NK+RG
RpGsP5kNsNiv3dLiStywJqg3KPpMbuF0xEya7ftaHA1ydfgzQZiFY+RkEwyp84J3A7Mi0+AQ9xuG
n/olx2lV3Kh657ImDYys2Rj8uaMUDflrpPFVCxsyb5+tKm8y45nbd6kw4O5Mn2eG4scDBKHx3Led
1GhG31G6Yb8LneJr9bBUO2nXgCIuH6O4/3tASIxUhbrwL7kmmmOz55d9cgr/qTygNCJ6xkOa3UrN
CrJPlQvgC27IPHMRt8ppx6yR19pw5Vfqca3A7DMlBHGg+ky9jkDsCQzzjEk3q+EEiGRkp5F32J1E
Md/UVcRlZa2Yvaz+hyYRmilqmks+U2sUoEIcyBqZw2QPlgG4JQqnVxNCIoNkvWqNoBXWrFY4Recg
BNrxUYzNwD/EpKDpwhSMUQLNnV0lsXfVRRYkUaHYX0NdbKtjwNqb0BuQClghcI9O+E6+3O2AYQp9
lhJxiEVWKGdcvj2Ah8C3XiEu8FirmQFRAHfOQbSZZNT9NsShUYuiInSzex69qQWabPaX0tkS/rfo
m15lEKI9B9dQJBF0OM4SEOjXZ1zjwXiRbO6pQ0XgmpTKQw4h5vwlm4ZuKykDzyxP7L5QXFEvDSXx
sMq9IEDVeqAawsL4QiFA/CTRmFzJbWe5zgK2+wjsyRo9tI4NvB5gvg5fDrcEKF/ZNGYXF1U8v1lu
MmC751E53pcpY6JlyyqOJumVPUJZm1O/EInqMwPWF8tEP8+CdiaN4POp23nvHjh6h/l55Vx3xfQX
V3/oINni0joFhy5VD4ZBtER8IvDLwt/Clbj9gNN9+e7tDCT3WVhmEcjN5C8zEA6rSUlS3oe7dn7C
z1hFXRwqAGtXyHC63gjFX10lA7faGh8hWiXt2GHlhBLeKXa7VCC2q4IJAku4rQjl/48hL+bjP3z0
+70IvfTkdzaM/0l/2abRdXRPVVptd2la73/L068XrKncdEjhzjZnv0qgPrvfyrQWXFbwYnuxRU6q
wEzafssv98Zdti+7eZY5FYLGPBd2CpdSmympx0b1KBmxkzEd4sMvUHN7LnXldvQRQ0HkJs5vThIA
TakPwg0Q07wChkz/qD+69FBY0lSzvIM08b9MSMLq3VX3QJ7EZZOU4KiFdyrN7INq5JB1RYR5LM8M
P3+7lEljMa4BwS1ZzLz4n8jCJK7vG826SrpX6dRlAvgIlKljPrRMlm2n7sBjoEMr9RqUVheFbBwT
LMaJovWEGn+qPR4Jfg9expUdB7kt7DZdY+LZmMHjAa9fOsZ1/vMFVEqpBerQlsQ77xXN7Re3tBYj
0T0VtdGnayF6ojZUO1Qz/KZ3Dwfy60D7gYB9VKTVxKsEKeyksGKw6ItefdKIX/bNq1/T6AMwAscr
tuCCUbuq/YEEGI483hn/xguBlEz/iK6tqozq3TszxPE+Hv3dvBHO5BedmFL8xhFnh/jU9xSK6h61
zfAcLul1ZopupWVgPIT5NpSXFygHGPF98rsSPtjESWNWq56gSat+Y67rtldFoDyzMLCn71MEMedJ
XeBcHtTGcghF1CHv5iMiqWv/N3FAl9N2sOfjb2DEYdwM5DIUcWrRvqOGiXte9Yw4OYoiO7FDzw7d
0zX5eqdbmfGJDrJNmm+nY/upG1siFwjYWQ89LRc25UAejc8GxuO17DPupcjNuWjIbEo6kcJQ0FP4
prK5m5wYC7JcqhDsuTorkLVx8h+vml0UPuuUDZVl2hDlCvRwLu9FcjFBfGS/xa5ZzGWpFTmRGkLf
uKf6M8Ih2PuyCusYNEaC2ggTLSWtMl2dJ/C+1JswFk8r8BFwdaImfVDXGw68BBHembRFJUE/4TqD
5q6iKtafsCMkjm5e29P+QJjpCUoCd3/SQIWIAIUfJzGJaUtwc1F1fibgL5isEe73LtNx+4ljUCki
u45W2K3MsrDSDdz1s368dvUAFIssN+6TFj0lpPnuGy2aweFdzoN/vkdSrgCBKdNcNeUWOrp25J/K
q66owKlzyE33GsbLMRHJ0+q9EN9NXVF/px5ZJxcRq71UD/AgiiI60ZfoJwaZMf5pLc9YOr6+fBeO
NvgKmaLSFUDsv5XbGF33BTO6MoyypXYclrtBUpb968s4/l6As5jzR5ZAXndJ+a8yLgEIJQBaJRuP
OzXTsQqRSwGQDas3RX7MpO677jUOvRMxwoIOIQcGhd/L8HWKGT2841E9vIEsLhtMrtHzpLFJrTke
VWfj4A+jUnl4E2ElgcezX4KUc3n+66JPNB6X7zQWnw/lSD5QmDymxz31yOCSRBaprYTlK3uza832
2L9JOay+nR09tWYEDioTqGuaiDuyRz0OOOTQYe6X5RKT/ZRjt16qgAebyeFS8/4LItxnKfytHsdZ
ypd+9DXwE01K2xdGK9CwO20TRE1cjEyplLj1xiFqwQ97v/6QlbTde/yQhb5Ok63XAIyJd+gTTj0+
bjOpEsNPZ+qj7VsqBqTXlPijgaascN+/xJcQWwRBPaIWgmquDYDYjdlZpT7lAad2AJJ7/lcMOFvG
XWxZ4oDuVKQSc1uPSjQGwdbfxn+I6tzbCBOG9hPtYKPspqb9AuHuwEqPgi7f97YLPZz0np9QE/CH
xFRrlcNdWBn/Iz4WIhPdCJ914b/2YEvZ1PC+kgetZEfLRdT3OH1yVTknceU4VSkmaZI9mNnYonLX
mMlvugZIT2i4/Trb4qZUTXfs2Umby6wZT81B44oLEfG4DO7qGVd0dsRm4PwYwaMxjPhT1JRFBVg0
Xi6xE77wHiO3EeWOFvcpVHpqYaByVvdeMUHwraBKeewQ58bjH9W94VtNbwYV2n+ZeWPpIWrAMT0n
72FGaUsfcw6rZgzFA+bAgaHuV2yrce3r0P0lc8/nvElVU/tQAK8sKTxI7NagyvycWtU1240MxTIt
i3x/BgkbklSogeXCpWs/c+TOdLRX2JrTxdAadmH2NerTE7M+0/DEhVYSL/yaHrE+RPGPjUqacH8B
nofHpJFkSrfFahsV73z6BHe5dDk3q2ibNUv1MvdecyiQBwF/+KASZIZXsvrw7DGnB1gZ891m9P98
IksA5V3NygZjNu31Ow1GqlIRWiYA4PRoxHXmpKCsEn7SWaKIGJtkPiKkV09qZfKaS3J1uDGBG824
3hWudbeiDDJn4/vxwsgjuTGfrC+pabRdFw4Mo5QH1LufZJFnC0P/2aR0omPCOa2fv/7tKHJ9glsl
oCYdImtOzbnzsLFX6Xzq1yIjRC4wvScSD37FXb/tv1cMVQGwel14aNMNFvdE0tURyy2V/2H++dJ1
3dCLuT5i1K0FwRufS6f7XNm5Qj/LT7m1+580js76BKigluGZ6bOCUQYi0NCgz06tz1OJ/KbZ2erT
eUazhRV7VUuZvmPAz48IK647x4Id2tILq19XZu5PfkW6onKcLiLCid04Ex7LlA+c+P5JC8dnX255
GYR2lkG7Ns97+5WkiPZI/7XbH8+IQUGDOP2d5W3TULvzXUkpR6YGJbnMAbEyJm0JBRjQlLMR9naZ
oEiRcRp2zqf5Ab0IzhxTY4ZsM5RVR5Mb3RxmLD1FWyjtXHB0HW9yiJt0tSN8xokXBvZelwcP+n4K
UgVlMtqNetMpM/llCYFI0ggxSCoafjPY4MyOgBI3AZYvnHXKqeFrvaM101ErbgZg1VsUSuKBopP3
meDwu0P7WVeo/g8At5AdFVGmTQtskC0dEntWvWG4TkIJFSZq5BO3w051yIrsxxKAU1I47N2mB8ER
10qtT/4PXq3Vry1Th3lTfrkJhmOGGiYjEO03mWD+eRMheCaPFfE6qJ1aTP+spwQW4NfZ1iaJoS6/
dRdJ2DDjagkD6cmRMJ7ECU4clEzoAvqbDD54cSSAHEDnpMKAOlTdwPnJCKncxqC7pdQ4sE61mbu1
DO3b8nGcO+9cBe8e+v6rnBT/r6RHJl8EQn1lrand/Fo9RKDQmI2nEENO2rblE/3vCJlABHqNMuPq
eHftXHKrFQbTmCkskS3/bWY+GuBWz8ahM8cRXTnXsIXHBzij6PY/QvcUCaQvsH56jR5yiiRhn6wU
JEXTGMCakOeZEYeyyqq9a3E+lAxmj2vX2MCItFNMqardbfjUINEbEmoi88yRR/dyfdtglnrvwxVc
TIJfdX+JF+ZdqIQGh2Tr9kfzEhZWj308z/Jcd8m4b4R8ngGyC7Jcrmgc0LRRFvNPyBr4q+dnJE4K
mQ94tp2+ZaNtA0TwCKvFr8rsKFiEcr9JDnD/YcUPalmORMP2OVkOIipHMkoZxPl8ACVUpTTFEdWy
qWsNmZyEO3JcSBJ3PrVizJevQlPKVklw7ZI6PX7xpZ8ZbJaurgz0GDkmHzFJAx197pBdlj6vFTve
DLjLThsr67RIHzAkJPt4cpKuedFDtFhH648i8wm7RbX+clOZt4KOqpCdnSt5uFw6Ytxo9Rcje+D+
h+FfI0sNN2KuDA77/mGJoqE6XAn4jTW5+lfCXFN9TpxVC28RNz5DcC3jfVEA8QB8YNVkBurfApQa
w1sCBfZ3LCCC6Oi7PMTMFVcCa0oE7tjumcoNx9afRh+pjM0q9aS1C33ZdwXdVw7wEZwj8/t+BHaM
lXkumQoPtOkA33WtWIE/O0nKAMxNlhJ9t5i3egNCeKl51VDxqVJhLztPXfBIdS0j1O6AFsdfOx4Y
PPwwnXw8vR0+21MEldIxEibyYjzVFw0RqnW9cF64vz4dY2RS0t9hRkUAweZkGm47Z8qzBKwVFtbY
q9Wm0NYjMhzEFnhRKW/0A006Pj4OFRNSbrF2+WEzpyBnYh9MwDJUyhCFEr3D6iIqE1GId0eSKTsL
L3kPyJJudtwJkVWUdNm/S/OqT9YCB83RsjXFHwKRFfgi1NBF5XkurhzU+O+UUEphwgq3IiD72xKy
wUQX53A4HQWzk+CiGdOk1e7HLkZ20UMPpJJQZq/bvHvFWfkUWg1kFqZdAiyj9Dc/wgwpMPSmGMI0
SN98om3TMkV7yp1NQwy7z4zvhUubCgC2OaXjNWYV3PYtPBeM7TlXcXVjc0D10027LAO0dFUiWfDD
DQeStn+5mipNgw0EiQ+I4aMIXIY4IANGxraWVLknQKmZatR010+cBYZML0jk8gnnZ4GG5vdXXf2t
m93dhPvWVTSoE6M+JLGssLY/CzEK0GsyU30JJNeD6TJw4vpeUfwYi1QGxQ4DRSRKlKqJAnH9Cqws
jaAgbnAs2OoCCX9QiefFPyQjM3SnjAoZTIw8q1aSX5c4yUNY1k9kogI4myDIofcP4oawazfbEg/d
OiRDF9w9+sdHG1Zx0SuGdoGb9mT3zhN6XTd3EGuSWN9bLoaHNXTuHmMmAIKeAs/9PUOnzLdHrPX9
JevvYlp1a+Zp9eIdQ517McbweluyJjLaLIoohKl/2+eSIh5xox9ABYBPc8kzgWPJ9q640/HRcngb
MJSv6oYH/ah1od7403mgs9MrGiaqkc1L9BRRge5nj9pQ8wAmyFm/G2nFHUNV86V2yYWv2+sefHGI
PIrVnV9M4SHRBLReRCKBSyYqyZrRde2hv3QTqBidWsWMLnOEAj9/DgAE3+ahWAf/qkmt8JJgZJuQ
EBAwRwNU/rNZsSBsevJNcY2++yn73fFn7llWSu3GTJ1e8o4wXdDuGRXum6Jh+IydNkoTg3yudJua
v9kOxAgHBSsCfb3dTqGfkQbE15ONvPHXUf89OeMVlwnIzyKjigqHwEwlNgm/wNs8DPBtzUb6knk2
vjkcp96fZC11AOgIdJltwHrvcBEWtzDSl+xOhG2AoP0vEudSIJCBZRps5udjAXKffGIdKcG1mN9S
yoI8iNgf5Vn0zCypAbQVdxMTrCahVXlWry2Bfqh+ey8e+FLWaT/6Op1ntTsZUQRold/2M/laEkdk
5MwUm+9xbQ7g07gbsBVC/+e9AMawng5casTCwciZlZ8/Um/umuNS9OMOVmcbSw5Ohbm+tOXnVEC5
x7TPX1N8TIiDW8xJ8/vcxEbp6j3xmYJgB2rim2GeznYigDSp0rNCwTBq1peB1yztDyn6J/gkFsyl
oMWTR3PRyxozwn+j60IZIRPXWSyfQ2nyHcAy9G889cSXa2QdQzccnyVx1CltPH9mNyZ/RdJDpnN2
ZmcUZldHV8snb8GrN4X4dV/B3101AtgFEJWWJF+lc60lL1CtRpEdBTCsxdHPA6G0A5kNiC4UxWBE
Mc2tI+U2xbykgFaWILBOSkf0IizAqFnsaIWIu1qjNzx7Enb6WuEpFNKLYW+N28xZdHeqNEg/blqd
dQqRby0BA0rrGjTacPJg09wjeML8SVHOs42eUDQnCxqwEt9eb57O+KpTPMA1Asr6oM9tPUH1N0p5
lO4/WM7NiRxaLNjAxKuOA6y9mzkacpDs/gVq4spIDex+jnCytC4IhwPpUYyzYtNUIzTYzshjobI5
lEHOcxE4ddl67PQkW6dNCjcVFy9kNJadKCb299EHUA4Ay9PWMLFshbExwNpwYSTayrGelnDk4SrA
Tg5kiMIz2sMyH8/lHV2Jn+bTNRwTOF6oS/+0A6xxZoeAA5nmulTlGigpkKV0KRjmzQ1sMwYPXPz8
4aaclS+DvPKfoT3nhE8+gTFelFBq/eanAtDLOHg74whe6QL4otj8T5WoPW1hxbh0S74jDJ10JQnW
wjQhsRg3hN0JsVSMzj+HZiyga+Yedc9s64YH6dVLCuVvWByV+LConEbPuX7KNdhkhn++S2uvcpiv
EAwGt5tWkPO4njvidnWNQJ2PHFA5uig2Qc3Nx6t1sUTiRbJEoPePm3AievOh7jN+Nuno9sMI5Uh7
pQfkaf63xWgoycUJFWoTI0Hbd2Vq/WB5Ww6Fbk6vrZl73f/fWZfXvVy9e79jdIV+FLsmx7dSGtjd
6Vo4tCAhoH9ZgL7JZgu0qC64sZE0D2F0KvlQgRIPyWpGz4OjOJ9RdmoTDmznXngii2gXh5sVK2re
rYTTPB05gOURn2qYd5G8NRIT1zeNZwmIBiKycsswqYAhyMOP2GFvppOKVfq19Lgg3GltmKh7E/so
CXF9HqM3hWLTvhys+I9wvZD5AG3/oDrswK9dTjelDt7aS1SjcaVDGihhogvUWY7jOW5We5+9FPoT
IJuzt+6mBYdOG65Q+T+8Xz9h7hBzb+ak+NYyuWpPr6yoCo6ECypqIP01CgKnmHJkSp1acGlkOVw6
ZsNqHqCC6wOCdCVBaRGB8oUcvBYHDT+5pyBkPKH2bWVcxjzflp467XtnPMkxnRS6Lo6VOoeAcm2V
1BpytuKwcOVvDKjdHoXB9TIpXW7mwWt+xZq1BbzNnaXrBy6ekhwzMs3vApGjskdfdbmCLYm3fDE6
6YBIV9igC44/hIlBaA9YjehaPmb3zfiQ1HQB9e2ypKiU0+sq5dVsyApfpAcvgoTl8f3lMlMSwZqO
Bc1nBj7GP7qEdTdwSEwtgAIoL0FUzz9nimhCwoEHwNWdj2WyH8BBTigihxwzifss7yVinik5Jt9i
fgRvHgzsE1j37/sSF0+JL+4zQOJz+5RHhXtvHtbOST6Teab2dgqmWr2EQYsKXLAivVqNC0yJ43iG
fg0tYJqVEeOzv6lB2t/jq5jz/TZQLBujKWy5duCHtgGN9dAoCXwvixnKX947+uTWt7c5iE43oWVw
dBhbKhzbN+G5CuRQusoB1o7y/ROFgRpOcSAmzC4bK/5QM3I8FtoM+d6+8PVXZ3ZeVwQpC7jCTjeG
QpO30oJlXq6uCi43DO0B/A6Bx/4Djxd2KAgWM1LqnGg5YSqpqea4yRA0DvBWQe2P6MhNXtAj+eXp
nbmR3MO6Q8lrV3NK3CJcdOqepnL6lFsiShPNZd0FeZR8Mcs+CB2x/ss51uFLSVKQEVXb2FWPUCl7
C8Rbdlivnha3du7MdMC9dTHWhjuIJcjZ2WLgL1iJ9+UIDstqOKOLGy8ljIbzmgtSKj8KedAjF478
q1ltuwduJ/uA3ba4Gxx53hvgQnrj2GxP09SKSM3IYNhjQe51npmPgPxua/mrFKaM+Bzk9L+BlWfP
sRAuYbq5HVgRAXJatT1v+7R45DMUcL96glvdvnni8piv4ipRwIu1nf3Ora5oUyDfMQbEtqSrT+ga
Ey1JvvpcZkax9ItIc+sIzDuZSx8BYEVzMpLmYJtl5lAEIG6z6b+v5GzbahZlU57xBRkFqWodNL0z
Qf0FmI9CtiiDR2/wApcmrnohcjt9uzGFBAe6dw20MmvecEwlt98ZkAvM53gqeYR0I2WQBYYNBzoC
9m3rpfZNd/sLOGBft7LoWmPkFVRk4y+MaTP+OQcEYAIQVct90BMJ7K0zesY5QnFz9S65xqCnV/xY
cXSN88qEYFm4ndtJoaYz7ly+cAWRez4z0JNkWWZHb4EKp4RpV0s+ULL//rA9Rwb3AXcTr24Saq03
hiuWajrIVLmJ9otfsYCWETnnV9Mezv1be/+6x9LpUKBUyYvt/V9WSlhXBu9L2Ejn+GazVDuqZr3R
3TaEe5lF5og8zrC9QEvuVYkMa21eVgzqa75xpGZHNyIsc5RQjxQry3dU9XGnUx5f1FXqLpNnD53I
J6acelDtrq6Efku7NS1bA1HG+bc0duaLu7pfJDiSyKPB6aGo1olIkfiLWBHruUx0yyQqtGfpOEz0
8FM+47qSLTMGh72zOv6U0fc8aF7zcQALn0hKzXbPgMCF4XHUev/w4bjwUyZuWG37Y9gVTvw1n4eJ
0Ygz0a1vvhDtonLZwnH98kHHmqkdkkOAxvt4uJab8kEc1h9vQOF78Ed92iPVT1xP9GT2cToRZzjf
cCWCa+fr1uO0A5weNIyPYv0wtfVz3uPj8LwOstA/8g0pT12arczETHrz+AHhjLzp+idXY9E2Yrw+
M7vDFaCE9Mxm8ERSNlzdvX68QfGPL9GKYdEcJzottgIbGdqXMZR8gGZhK4aQHJlvv5rY5bVdocf7
6IN+5y2ty3BORnLgunqpkAbaz4Nw64bY6AlbJNpYM9/VXhPrZ+yC6BPWlB/JFMY0arffVUzLzNXa
9TWpM7K0McR8oIcOZInVxwktcUbGiyzYYoBw3BoRYreSBzP05B28wSaXx5OjnIWijQcwxUYSnSSu
imwxYDpBNnfLuLWGVdD9JDe+ssOv9Zm58s8vN8NqBo5BrAOfRdaJO1sDqXbxWskv+TGipf6ubPvU
RkPd14ndLJBaS3ZJ92iErPDvpwOPvP38QleVQGUyAaYwVK02wMgvq70DbQAIg4MtkT2kEqjPuO7w
Woy/xoZZjzVuH4WHZgUl4WSvdRg/d7VdZOmDys88egiWU4y+zpBFaiBcfMwheSbKMVJw7fLloB1m
54i3K+pFxlyDdfPicEkcEnimZzl1WSmTvjN5np9DTPHDW91uRKVvsMIrTZ4L5rWmzT27XHW1XtMp
A2V7kE6AqFZsmCRu1wIFmEFLf3Gljm9ne13IZhVSbQB7V7D4cX7aHg54jDEafu4mialiifl9UnUn
M8aJhuLW4UvlUV8o274aeMScpGXqAAVFhpVcSANTlUPCh7qT4/coJmt5RgMIeQQP20Jt5KVPWveO
zgHXT7ToBeJRHczKQ3kEOsHi466Mr6Hp/iOTRDUJEB1zW8dslLKzRAhtAVJM4EOx4Qm5RRt90F71
f4G0/p/PUIbfkKgZs/DrK5BaMs2Dy+f+DJalsspztbZ2vVQWkAvU/csQdLedqayCVmRnS4Oar/9W
utUbrZFZt3qHjOLlWl3H+pZDVScR/VEn/yzryCU1qNw5TFM6IXIOuYKiqLs4IPmMkAr6drlmYP/7
cmuqEYXOuMOuvdiGL5BXnyFte8wMEgB1HR+jRUBCN8lSJHm+m+l9pp2rbOSRSFiJt0abMATLHkPs
uCHbVjiPI/2DXsEaXDW42gwDDSrm2i8gTWMTHrOrMcuTzOAEbiXPa8P+P1drwI0Ncd4N50YIDw7T
XbASHXcFHg/1p2NlKkzFCpynmBWPaede9LEcgnktlGS52l6e7gcdL8mm4y5dhR+6lU4r8h0LuhEA
ugJo2F6Om02QRLxT2xNhwqNRlg6HEvVYlhV3z64o4nZVwEwU1Gfwil3X3gqO4KquohdqNd7oCWXh
Flv0bEjPScmCe7GHVrGLH0Jb+In5MzNSfslmKBOqwBTVp4gSmjUJT/WBlC+gtblsgmV94EAaN5wo
j1kT4tGJjZhVpXo0zdztqWSWXJbdhx+QAF0wq5ncrwLqJiR/emq+83AKPNB/MCPQV+jVKejML31w
sFU13JRrsbN+C6utlmrTmRBpqJPYuP0AW656m6Cnb0aO8SOEb4/ToK0I2PGbie5xZly/TcJyHKdt
wv1iFn1WhJSnQX8DRt91cPfn78FP4J/52bLMQVq1MTn+E9Q0rC1VrJ3EtQGfna2t/kQqOtVHHbb5
tZz3auyosVNs1oVcL//1OYSRPHPR9YD6CA1vC50MJ2gqtKOSMmxOJl4dXiJXTpZVY96QJUSxpwL4
52bLUNMguQM+GWa6TL7NHvAkBVnTNWJK7xRdhZ4n6Vn8KMyTHWIcKNUt+h1GHGvKfsqsrGSd82sB
Mq51GDqj5o6IHwLRrPYv5s8EgfmTJOGuBecf+NbZ8thwAKvBNy2czaq382IFhy6x7W5M7q4q6+71
Kkv4r5fVbgEOaCLzK9XPdHMFe2Tt6x3ds4XbpUXlAZ4KupOmeXj1VfSMP5Cg6Tuh47YqHk4w29KH
sdbl1FAlDv0fGgxbrdzsWNTKds64aMQK6FKWgk8ES2rPp0VLgMXdn6/CPfQfByKdiqPcuACWXxqy
vfIrfC71bM8BULyktvSTSoQnEW37Ejx8lLYwQHYKT+tDOTTtWS+QISI7jAMoEhOZF5a/Kaj5Y9CP
omZVgSG+FK3asTgqPfHuW3vO/6iQ2DAHIxeEpoKJN7z+iiqhsaxiYZRq3gY8aB7oxH27HvkBfAt6
jCg4tn/q9wnIOLqojYlNwbEkJCsBWq0nbJQ4/GJM4OPwdEpndl61Ki/U2urb/NyWcQijflk0SzT0
BzerlLNFsCljjKwUHPFeKJKDtRcCcC0Tiy8BRkJcZ3zw61hH3NgDRAfQ2M3oAZJ4itIhoADHpECH
afTLICCyFQJWByODbpGueVJsp7x8EsDV2qhY/Nyaha6avQ0VlzX1G+QakdEC9CXOweUprungEyaQ
AtR5HUoa0UGqM6wnf8I+8sumhj77eynXsr7wNymEYcJF/kMm+7hZ906pL+imH+RfHAMnu7sQXyr8
P8nCMKDLeG6Mv3txDkyw8aWx+Htzh+iqlOZm11Rps+DGMDqQynPjh7C3rpz+M0y2oS4KqKA6e8jH
GZaEhVuPPkuvtXMiv3C8hktOWaMHxzgu0KtnVIRvl1R34F3lt+DDUIvNtsC85r1X2OVkQ9BVpq2H
Tokht/H0eeUVavdh0OrHrFBPhBfea6nCxGGfS7I8XbzrNQb1f+4x5fu5DRP+ldY1/kVbWBqyRL60
gJh+OW6x7nSOYGJLb4rE3ut5PJ5LA0qFVxS8YTBL038NtQKGErUmSdMasjVbfliK3JipN3OM2tYw
UXCB6LqSDFEsKioEpYzdnaQ5T6ZsXV31CZ/7y5M7JmId4+kdvVlZNumFAcMlAn3mfZt6NXeVCBgA
ECqhfnPgBPwWf9sTCQqT2/aiK9FY/eZdy0R3JF8jVG+bVhOsNrzRbwgKABmJ5fhCIW/3CVgzyNtv
ujF++y018i8pZGvrxHg8I6/WVl6ZBthJojpLqMGZZJAsrktY9vf/8AzlQXU8qDNocpAbsUO1JYUO
uPK0yyhTaSMaSZJoU/coANhYUEZQ9B4lMUuVHCMtgopDhosmFFWlfvpdOnbZnvFch2s2Nkw/HB1w
2wqxMs1GYm7G79QaQtydcxt4s57c0//bdgZTZKeYE0iiwqjezwVxdFgVHqrxUfS/BjjD0gJUvWIS
FRyiobdaE2S4aT5XHgVZk1hs6A6dVIAUdHufIQJUfMC2syTqdxqQbb8xIZ1me/r82UKziyWj31JT
wBSUU3TY8xfUeuol1UsZjat4RFz/kr4mBYcgFYaCYgNXuORlCshH6+DdzNcxQ4tUszGxScaGu7MM
r2zJZj/UEsGQrCJ9NFtOH1Vw2EL6jKdReKLH+oQYOJFOy96x9ToilxFqxl0/CVZyZ93RZ+Cr2nQd
i7S5WxzaLGS9THSXDDoNw6EuHBb1jfN9geNh5l2JindY0CvPamhWC0Ws7+9B7CNsfFDEcLoXlsQK
j3nX5KAQUyGYowHqrUp1CVvY3OMISk3yVDHiQ1iIdYw+1XdBa9P9GNfrmHXJTrqIqGKIstd4PmJN
FL65LwlFRCctyDN1Dcbge7dwEUZZOjG7XXlq4rJtRlKwz2HYFyaND8OkHgTdOPzwxmqqkJIizTPw
yxi+Odx9Gzh/j0MBD3CnQlb1ID3+t+d8Oj/bapAgPgvH4/tfbmw/d3bNI7S6LZ+2tOOle00pi41s
mzfOHXmKU5ee7KQT4R6GBSHcb3wa4/J47O/7RQQgcJsuSpsYaGbXWMJlUQNEsjxyr827GKT9QQ0f
RcQfda/m3OdGJ05dq9Jh2WIZAy1rmwYJYScVhLFOXopjhZF6XT35Xd3SLpkR+cZ6MQfLwb/RaJkN
WzMwj2ty+abnU6I29vJcbXLW8ri+gczMYJL4nNsqDkdj4O5zzrdYroJMV5LjM7rkUGJk4EKUPScz
0CrfmL6ex8WHY0hyd93Yv36eeEWQLBKbdpV9VXv+tU02i4nF98myl+Sb0FJ4wRY6mGVmH6mvLLGh
rc7SXQGB2mL5EIa9r8x7AImh6lPbV1k0vlO5CQmqb5aKDa9SMW/6kKnM1yIp4nIfgMD8xzXQxsS/
2VJgz5phnn20dTG4DfMBOvTqd6bCZKLawDUzGrDMkXWFUe14oMuV1i5nVCcgnGxREemMUD4CopRf
0x/+cs7TgIjMxTNnucc7oih1++u6MJD071rVv957UwmoQ2mBSQsQNDRfvwuePGPWHYOj1Vk8jhrV
YvL2FszK6FwtPGkVveM0YpFhaigs+vjBjiFKlZE+79cEZL7dJC2HeTfOS7Q4AC5oeFpDoG/RdbE2
mHxR6aFobXuDMDOZhpkbDQsk8lC7uBAQy05BgGEhrnfiotIKjRFDZArr/AQ7oQS4q9YWwzDNd5Nm
4DBK93VAIsBlkN+UW1Qp1tqaSFn3EaY6BfvOEZvaSHYwZ6XBRZDgR6zlxh8AEvxZX9nnXko/130R
yswGvVQrNW1zNP3Iy70lYSftIRLe2rQNTTr1ec2Ho2Em3DnvbF3QJmDehyVxsUwxGJ3C4lIDgRZv
0ks/DRTuBUarm0Xxsn5FpkkkPkZnE5sH9rRaEitJySXE6Eh9Cblk57IJ8ZWtJu6ac/16B62pdGlN
XNDSXEDJrdl53GAEAARt7+VluXhyB4lIvZfWXB5x51HULXlJUV+zXMzg080aycw6H+i1fSbyKBHQ
6ZtEjZhkACwa9U9uS12znW/C7paLB98c7FZHgTx5CpkucNeOxu0Ir70gbYVpnWYUTPqa3ajkIMKD
YOh/mVIEs/IxPQ5ENenM6qJQ+sFBc/CsTWqERAHT7TV3RqeIbmAO+JClaIm6Ga7rcozQlRCFDU2I
/eR+hX218uoV9d8ML7hIG2snnFel+YPov4ALsGNUZtFnqWxrydNBz5XlfVH0gzh2m1/VQ+agPqU+
vV/wsB6L4cA6MwosaZf9uCPnb6Y+rlEWbkX8Ih7Ko1wNqOKdRsCM0iHdMfuoVd44WkIloi+K6BK8
HvGZehAUcOhKbtucwjb3M7Pb6vOXc2NKoSJnrv//B91AzSBJTlHdz3BqYKOWi8A+xO5tndSgRLS9
MYHQx/u3+Dqa8YtlfKJryD3gLWQDciGx7LNSlGnKKVG2ONsFZA4xguQI0jnqKajIC39kiVw2fTJZ
73AZYohB/Li+JOm+IjWGn9B7aYjfRUHZCy+UzptxGovlQo0KZq4ZfAY4dYlstJQGCgx+qUKwi+WC
a4xb92cRWDsL8biC0YkRmatk+BroPPYogxrTB9Hg/sTEuqlqaRz8Z3k3XYkM5nAr1wOMFALXOurR
ST8Iowmy9/5EPGXkGGWBR1jB9rgzqbxQ/BfqYWBmRRd/z1xsvaSRt3ZiNfo+ki2uIHQ/Bym78pLv
9Z4WY/W2fdh4DfnJ2Nzoi8XYHz7FiIdLSAQKInqxe6NZJG0G17g3mPG/1qoVtFSgVxy/csa/d7Tj
1MBDDHm505BQyXA9UZC3qImW2cHyTH5BdsuoDuNGezxiSpGvwjJXMwwjf10vyz6w2DXWMd019pjH
xKfEC5P/lUQWmkGhiToJiUUP1klkvEDfmgUCw27maeCctYHHQbqwWjM6bvlNmbD8ekWQT72yf6/T
nkElNAftC0A5R1wDQOc2Pj3DwPXha8p6WR925F9455KQojJhU+LowAq4XHb/Q4pLaNltDvOw0Ufi
XIzQmk0FtHL+sZP+KbA4UPKmp8Gut6r3hobY3+yRYPBJNw/4fEoWClEbUYjFeL7TrNCwE+cWoZWv
QlXEWtFzOtbRLQ7dsdjfx8H0aPycrliiQA9iVWt9/tONgYRC0jHj3pX+mfJCJLPtl3gEmE3lXpxP
2kH0D14rAL2+FoGdfQJgbLGsy8Raxn7/BHo1sQm9TmZvnT1k0oX58fSIaJlC0KPkBmWTi5RHetq7
Bqf9+GAEPJ5HaJCxBY2+hMcm8twvDPJ9Tn+rkOdm8akSbZujKVcZBwFoavGwChbdrvVZdEKLN7CN
9Fw27rvSoB+OoztmVxFMCAgrhYALeWOOYoaHJpawdqF7c1V4HqoBHM8rjzXjBDR2IqpOMKycnhh7
5OD/c9xbDfBzPvi+lVwFnCHEV3hIlgE9VQfWZu/QmFpVxNOW4OhAaepdRguOn3MwruN+bmn0TJOU
ewJC9YWFjnIfX8oh4DYBmx1jC2N5aDIexHu+MzackXVBXaiSqmU8K2141Ou9KtD0/HASgLI3KNvQ
ig2AeY3B90EBNnrpRN6ZNX2uoOZjiijEJRN2Xb5AFucqtFSCZHgKD8DkUizCUrxUQMBLy3kZcqXj
DUCIaY0pUCAlbiXBZZax0cT6N7r8hKnv1vUorqe41IgmmVOQw9J4GPXwEFRhV7T998k7JKVKs4Sw
mffPQReaXlmmkYVy2MY6Vxb/0Hc3lSHMTQxYp2NUgIVAbn3Ut1Z+9bOQoeczk+4e+we4lzpYT8+T
8OakL35bBVqS7JKrqdFy7uiQbZGlZsZnLW8vJJrBmQXkXl6U0HfEPtRANwjSw+Zbs7jT9jwV1Jdt
8hQAP/RHN0NaYLZ6wM2cgPWskHjJNEszpz7HiMiZG16yO/BZlW61eiVBHxDc3AsWxR9yDyDVMgz0
OLk5rrawoqvjHxpuof+w+S4nUqwuQswKTL+cMllaxNA/XYebGvfVkw9H1TI5fZjYE6uUti2iDIBd
nZXYSyBb2ttf+/hsRYWU+yOlnAcETI0HBQc8d5OJGDJDrSQxJAbuZ27pmNl/3aBNizs9XdjiEj3t
ROk3ABGinN98SmJQ9pv9UxErH9pJkxgsCI5MZSH9jEWRUOenxTB8oumd3+Y3zIgkH3qYImTSgeYV
o++nVq7ZE9Ky5QLoV3dIoS3PzN2dkC2OSATTk3rGzXDEe2XUA10WRzAZj1q2C8ZpxErCpm2vn8Xx
Mn1mEvxrJGjv4mPhgPgPWb1nP2DcR8bbeMvqFZO9pWCLo2o9HyBlcNvGULnMB+ZWYnIfZy2dfP/5
jv452eTjT8BybIX7EStz9Z+uVIlc6WFO5S8MEfHW8KIh4Um4GEc6crJ/zXBRJYTw1LXrQ9/uq5Nc
9PmWCNMO2qdHJ8IMeNW3TO7nHDzfOAD66I8d/OLuVAKWCmecBWPD8CtYP1YH4hxioqwJzzFCNM1t
XfcSmC5F6NuJ01n8K/YRPf/rKGYszs59P3oIc22PqTJUVGQginY04xiwAuaq4IVAMqsyZ7hzhco8
Y91x9klRQaAPoqS4SWCQIP87G3TkI39mcBxI3t9Wiim52sr0fUw266Fxcr+vqwBszsMyP+J3GbkR
uyGh23V6bzQBg6vTSYRlmbPvBq7Iythm4BX4c4Z3/j8QRU2tHkSh181Wki+Vag88TXuQOk2zNvBb
eic724GX2G/gW9HrTAT86wdEhwI8vn3wfQXZGGdu8BpJw1duUskJKSgSIc2q8jKxF9KNuXcMICDn
mjS8XEhl+64RUXMni2JjVyd91dE5lzggIW0boJW22ZaBgEYvNchV/r1U0neZiBgh+qInk7dHCgiK
cAr+awm5giPF9Vpzfq3Fzc2746IxA5ch7tkymGwubkrxiK/uZYwC2XDo4NJexEASH4QubeHbM1DF
qr2afcs5EZ+SuC8eCBxD7w2Wq33ifDQW0S7e/4xufIZ7VcLvY7zHPh6J9UMdc9N98yRIbLhgAL0Z
+n5aMqgViAi+JiNPRjn/fvh+zD9mIRdZE3ltOIKshN1HmE0xTNCX7F1eeIie4E+aHqVKAfpcDRiQ
sMagMf4E4FFERCklimWYSEp27Lo9xmZWJDoVClSUwDSjPIvySemvtL3I9b6aj+USEr7NBiKxBn4R
izMJHHBJcn5L0x3r2SXAztuHItZvdkAJg4zwJSCC8WjDWjHqIftSwgieWvnE1mx2M9PIGx99mcgR
DpXzVzGVgXIpH64Prs1ejLBf7r6Ua4LFAdNDHaG5fLJ8QbrYqbJu6f6f1dJck2hIV2RVuM4UBD8n
aFYwqQ2wvxIabkG5zbkQXXP6Le+Y1VcOl2ZdNVYnhaOv8qBk4khxCfvL8B83u2FM+GhFZj5sWmQa
REF0WIez9TIHCN0xuwJTG9KFp+igC1AmxhmrIbvh/+fBTTVxLL+snnLmyftIJ+xxchuCZcxmzEP0
zBg1k9Ny5fdRZLYt3Ly1Ysbauh1K2EEPAqaUgzZKCZZKu5ApYgxkSrupUes3R64DRQ0CzJXs1xOn
03IUHPbnsQpuovTFDDV1FGab2eHOhncFMyDpwrMsXU+dQ81UReloI7/LFURdeusRCQ/WIytQxFzU
cJ6I6Np+SCOoBdFOouePNoWF8Bu6D33ygA1lBk7mBQeLVGKvuJRIMBJoGiwtWDvXD+QBCf26Z2mV
flQYdxHAFqImrlpgHPm7vr9Cv2qaLdCGOvmjZl/Lu4foFemRfk90eu1drQgkJMeBJA8TxUv3fEg/
vxf93eLUSPE8LAmA+9WIGRgV2QqrfhuZpGTmsHbkK4v9LiGjrFcrF8gvKG0xIEqOb0/Hf1aMEjn7
Bzh3a+xFVeBpsNkKpB4Yim8O4e57IHQa2HTDP4v5CgwoXOO32nM8Pry3ndmn4SvXgRx2s+Te/kLn
cppDPUoKf0JqP2jbSMH/YocXjAqEu4iMpXm8a6ioK7k+BCdHBv8Wm02kEcHEhGFTapfHdB65BBq8
HVin39NqpjLcA3yAz8zQ6S2XdxXv6sF+9PSXfGVJV3IxLIryFOsopo48kLFgn2tjOP1F82CysY5a
E+UD1YBhkuz+m4ETMLG8nrfg136NRxtaHBPNAWTqerXkoPXSGrjL27MSbmYZ61FRFR9b/7gxKBY4
j1Dz3/WHUo0OqNhnQk3CtnVxBcd+TUmm4iGFU5H1f02DGqUgEecNs9bhr6UWoRHG1umpjFA7gY0X
IiW5sFT+dchSGi75Bp6x1THumrvsvaoG2rw0s+KjEn98E8H1y5hmF0A9sh7aBKp/oWvs1w1b9hQF
Im0zz4w/lXYxw8HDzKzp18kdysD4doooDpyw8Z6mtUogeYzOpIjMI2PhV9737dfEWfutiYgUcYGn
S7ZmkQYQaPpAVQsDF3v7+1C2IVEj9QjwO/TlbTGQ73fqodb/BNNix/QOUkWlvDgO0Y+l1zC4fFUN
J2unjRyhOyi7d1rRi/jJV+F7vtRB+FPmNglwKuz9SvnI6eCPKcWqVZje0UK8Zdq4TvjUtqlXvvsq
ycgVectgubXzJSMXJ9e1Q4l6o86Gb1nwMCUBr9gJGCGufQj332k62wsRuF9aWRTg2GWf+U3FcqdQ
6yYRV4w1iP1vRLU/1vCDuWMAHvOfDIqYX/2gC5laGFitj5u/Xqq+BU4xDTNqikDM4WY7ndlC3tk5
nCfbctNAjYno4SFEdRZkatt0qhvvMYsOuybS6qvNESFiZYYaBsPBd0tTZ0lJcYX8eseRl5ZgF6dx
cdvHabX73j1R8KN0fvCFX7hNSJGVCXXke9jOim9MGwrFa/fgW9kIpwevPznNw8xAkTZHA2PEkrq7
TMMrpIWOUAhUVbiVWhimYCR8o9MzubEg7jJrQMZRV/mtUsB0XfC4QmdX5+UQJE/tTOy+HIPHK19R
edIXhhWi3wHVNHCReh357GKiLvUSkDPIsTm8/NVZQfSjioSR6lTIEA8oFvqXiO2S1JRK72iBoNMO
VqITqrmwYBwKiJLSRMv7aqnxwaUg1xsLAuUZ0EFB3RXTg51lxURIP6cPWc2oqVSfP9GtpBtUgLaY
pMh+59wd1uxkQoTwwwdu5+brsu9sAcFyzerwus4dxoxHkyimRM0THxn4cNdv8DsH42S1MktSr5Nk
24ODN6fy1zBUG//3WtV8VnPBYGPD9fO0vU5S/29ROsj2vm+2NPs5whxbA9h/6+RM75UmM3fnyAx8
7yWP3bMo5wa1AtnQEWU3m/JZMPddYzz7Z2IB/4QwH6PdaWArDXy3nY13NiXnKzfZIbApqTJmOw1A
5zhKf6lfLNUHFRD56uXASKEc1R2a8OsAhNi7wInkvrjZzk1XVbq5k5V4jj38k3I4XYf0ahURwbmM
iWF/bvnYqKpdTJMsv51aaLgpNC1XS5gIL/+6hcY4oMLyKjQOgzsau7cF6IlEeNrE2eRH+6f2Sk6j
yTxBjGoGKiftDjiY1kqcgBmBbx4zW8Z39frOQr2e31Hr6tXm0F3mVcsoYpSwpAdutZ1YiycDnTus
NFu2PBceMK8UeG1mI60Xr53+GIdfxt3SGb3HuBdSjpCzXlWlnskzMz+pm/V3vZGCunwlWSvvtl+Y
E8cN0Am5suvRipIDn/ISiYFyGePQO7ui+D1eg58pRxGfZHlz2GMsrJZifpt2a9WfEF6mCxWVUNI3
Q4CMDjZUdNtklcFvpQU9HfKwzJCvGKrUUjrF0DNuGwJRTcCTKZUuFy9ZGOgAWgoZuvfewIPTgQmj
AeV8Uply06mDocouXY2wZm6vx3A+nvTt6L/vRVpnMIRFStVNaji2NNtwaxyqQq0zCPhuLFSs0WIF
hJDShNGGd8kxQXHNrN6/d5Ddbt2kxxh6vNh64QJrDLG30NObzT8z7WQT1xjY3ROeO/B8SMZvJC1n
S3rU94b1YLmgjlAvqa/IycG9blD6mpqRmUl/MIJf4KqSNx42hHNkoz5PJ8hZqC7FR3HFK1sdWQAh
tOofZ4Yhxcxvde9I3KgqGS6HRx00/1PWNqhi2qed95EFVOK3Z2udELX5hVfMh7ph1ICQ5LqLJRl2
jj6FRI9O2JYzxfbNwMGs78DomiuX9Dw+3+2gKZw0eo1Ut02M680RrgtKg4bST9USBmVZOiJtvhER
r6Sa4XqEyY0uJ0HE5y3z3pQNHpTI6qCcJigpgVUvy5mz9PVBFJvF2kYBehH4RAdrcOiILRCx0sLD
V9RKh0hvONEX6VTKJdARFwO4KNS6J7x5/Mtvd4z9DOKSYVabv84oM3b2bbsliMhYuCoHJ17iuJhx
vtwW/2hIdM/VkCq571mSeo8Xey/8urGiVLDSEVfyOBc2Ve4vyRzuorDTURIN//xl89sWs4Vt8BBG
YjZTm5xc9ijIjh2fs5RaXvueMMk4EIK0jX+BjqAqgIwesSVI/1vTbe0EbIEEHiYualP2uGwVtlx5
ZPODtlSl+hxh967PIPxIThULnIt0H7YkOnVzWTYI4nYTzbKyybD933ATpXCnd44fAdjHKXMsRYdy
EMMTWodqwwXUgDHYhz4oOmEI6EaUop03l2tT+9sHxuV7WGkTlNlIQ+bgSJmgNKbElNUN7Diiowqm
mKHuyBeisKKx5PVYqicWaqnwYLJMHukaBW5T4NP/LKDCV5PD1W62jhGKGt4SaFIv0pyah5aNi/15
OcMjmXWNC3nBvyJx+8k/0kMXkJyV5P4XLGdsxplzNPO1GKkWPRz6/5BpWGdsk1lpf8ngofRQnRi9
viWCDEjB6c4cyw+vVdF3ckE5UGj95Fpq9QAUUVcrhbuNOv707BJ7b0945xzgp5GOpERjbdLOGJAN
RLAv8IWlcl6LMvRPAXpTl0yxCVam8jYzKZmvxW0u01VfsOSMOsBqYJX5OwXHOy0+sdsnHRDUKlfg
jny0Nv6gwQq9dEzk7fCXlC5egHedHT8REcK9f3xfyw5OtQWjCTwYi7Bp+SMNGgoLy2Culev/KxPr
9B/RX4mrA9sql5q/YUyQaY655DauOAoefTcvScQ1YHth2IC0YilfjA7QJvoI67IKe4BWSo5wM4y3
DD60JD/gais06bWoXqM/3/As/xB4QHzBL14ol/C6EbM8UTEUz6g9rk8loQhFXvXZUG4Qh1Pet0em
MG4Hf8VrH5VQZ4y0RzhbrcP7yHlgmQqe9PNGxwOyW5bUPRXwaTJlEv+keoaosjpol1ZW+HCt0Sqb
yS5z/coSwIWqDtVQLjgB1wYINUkdgRQtF71mXaLiafg2ftHGvKpMLk6swtdnm+Q/9fTTQPoAkd2m
WBYZpsSIFERt5kbMfTvXR9gYtPxh0jzHl1H80kurXRsBCSxt5atEe2Hi2Ja0S6vM1NPy+d0v4E+O
CMVGOpguX9l8gePVVMCIkQiV7AO6GleknHIauftkfjpm3Srfj/uxn5R3Cu7NwSehhtiVivZD4sQm
bx0quiMN6UV3OjP3v+Vbk020gbLo5esrgU4NKG9pQ/lub74DlNt2Ba7JjKXtFIIQCrtZQ4Z+wcFM
3kNd24vr6WOIJq4GIk3Oj4HWY7cJGIDnUDBuKqDyNSmxZcYEUkOVCw2hT3QoAbvmBMZfl7ZOeC9W
r8UZZ7vwZApedJpg4ekhode+6PShzkLh0NX7d/aKz9MnQ5hiSUmgKoLBgBQR1rkkm4FgjC/+NcOw
e4AA0A2Z6it2MmDjlpPOy2lcnWXLsU/nRkxZ/NDwbel225iLsZN9HHyIyTwnVFBcLhotTYG7ReuY
6xZGgmPknsAuaBZtNxqTGS4HGNszTrXhrnFMhB8n9dXzbNJL/7tGHlU7djhI+f4JBVnLhiTWYHR6
UA/r+tuYNKlJSxD3TE9aOGE/UkybqCs3IzaW6rF88YK8Vuam8gmxsYbHiCy44byc6agL+EAGktvr
ZlTNqR7ozf7ywSSpV2Rvkl1AXvZo5kuFPYaVOTvZoilaIQQZY0i5VVxfz2W22+oe2DTu7UlOCfZD
E4Fr9WLbLFcqzkvFVKQ8/aX63RWmyM/mH5CNsi86up58RuYXXlLHgSNgeai97mlpWekadysFN/8A
FvxF5s5Rdv3GgDsVCekOtM+s19ncDZe78VASRkPMXB3eDyvZH0tJszMXmVFKAvOvknOeol1DpTJ4
Dwk0jihsc1/4uHwGwV/9ljqj9zxo4o1GOarbLr7nS9+VfN4/UEv/jfeRCOVFQHnI4Oiyv9S7EWTV
WK9svTpe+vGDWB6vH6EuDfWI3Z3ndytWljrphc6+UJunzb6a9CFYoWQtgp+gTTqUbgl6dRH39IoC
g7PeAXD0Nh9lf287vKk6oq+dkUokCxWMpyVmTYUV2vQrTdh5NAFObKeR5kdwHBpI8DDEJR6OeUof
9BLLiw+cnX8cqywRtc/Lxh51WLMPo394y7sEOpjYICx2C44TUSIDnUCL5LItoHXFrELmwzT4qi2X
HGH12ZS6gIV1C8/b0TuUPyldMG2B3ctq6fDbYQTm5DgmH0THupQ3Ix9DbTPtOuS/wm4pwjI+M/WR
ya6hrn64Q12aVnDP3xHcRh1Uhp+eNjOy+D2Yht7XwE7p3Zxzfsv9age66fJiyHeclKJ3rIUhmeyO
14DTZrWCPTmJvXidIzMTK7Tq5J0wnbNfIvNHEsU4gKfmHhEalitXNxl4zLDDXXqEVWnm3ZeypDlF
U61jujiE06q2us3X7xyOx+JiuV08adtjxs5FYyLgtWbBmknKooFG4vTUxtRBlwnZLh8X9jShA+id
puPVD2xqyX2Mhy0bVcM+UrtNUvpG691ZJZkOFPpPa8YRw3p0JkvgS6N3xWN1KmcbpjprkC+d/LNi
lo7sHx5X+ds7GpX5qR0zeCmCT9774sBhBSswX1fd/IVkQX4MolfDY6BBlNhMAFj10Q4WrVn4mP9S
QDDNpVnS9/sf1nPI2EMhknCJdR74Bb306PLhRum3ZkYfC3XS4WRSFRPJsg+FbkIV+JLxjefCDQ78
/zMga2ryrtuSuUuWrsMd8eOH7q2wqeIGZOd8k2iwqCWjf0ksSHKDFOKeUefmw/nc4qj5xVAMHews
AiEjsz/ZPWJ+qkRo8qm4NXgJBdibTvx7RioHori9hQd3NsBk4Bt9R98L6J2n7yNHZ9n1WFoGQ/5r
WRBq570gLd5SCtDFx4045l/LCkRZX1q4VMiMXFYG0Qzxshzp+2fP7qQ3N2I+lW+AREIftkd6QGC0
wjJeCzQSMZr3/1c656iHipufosCpiW0uv9h/I+Hr6ctUTaaq1XxkUbbixOQ0eXJmy0+0MchcbVsm
KuTZIFqfs+t0cQjSqUlsuTHsPxe28ydjzuHaplvKuPxtSrgt5MO/VZWycxBsFLlGVLQ5RERvilMC
Ae/GJeG28nBYLIoaLhrj3PYoHRBRIX8LVB5/3HFWRVHcV3eQPwkMvjA3IS/ftfgJ8PX3GMkaGUfQ
uzW8aQTMRFXtOXxa1zcd8T/RHqUVF3XiAUmwoZoJoAKt7Obl/3qzUzNX9rrwkpP06NgtwJJUayJf
bUDoW8aMvoAwqFNuFEjZ1j4+2di/pM8sqaMoiOmXu35N48nYZsgtOfle5xG0LCXq2h4FC/1t3hiA
no1Brk/ZhACyho1pAvKQrCVJvcWOyiV8XewHNBF0UlD2fhHhTh5aohiJp4pbw1G0dR3KioFq7h61
kEuQmc1d9qpWLkDJCkCOTu3S9ZKNFNsrnpPCmifGpuXkMumdOj1gR8o58gV2Lbbs8FKI9a9uqvjW
7SqKOkbSOCrVsba9mrWkYaqHZVQS/m8TU431cWjgCZ5PtI2Ae2ncWbUmmyOWb9qS/UpYpL7QLP7r
y3vNm0lZxh2u9FhtWsc1YyDFX/0alk/n/+XoFtn5bBvFPVVx6tTv2l1ZbSlPGUHotWjfxyyk93te
iVys/xCUFWqnEWc/aFpKh9EQUnYKEk0T1RlDjI7e6rL2haucTWZvLzVjCV8gpFwHSUry5/HY2jzY
Q+qv+K2Dj7a/lbXe00uOLGIZNPjzi97bJvyv2eGU9OTP1q3iw6Pr7ZnGf8h0UAjYx5aajfk7Xxj4
VnJxujk9Bg3lTMI60hqczABC6pf3ID0QRB7Avz9zaJ1R/eVQDYidX8ws9MJaRMrauKDt/AXFvbzB
jGLoFmfOrMa+NmolCAlTYWO/dVPPvnFSb7RMwj+6EYaiQFAd0fPzBZxlxBHDoq14JaUw7U9oyd7r
jlbvXOtKsWdWaAv0k/fYzLQHjoF+D4eMo5NLT9PHv1EWldvgNPTpATpwUQ3r8SBHkkjwaQ6KD2Bo
5GzParv7HwNFJTdRN4TOjtL0s6Ae98b6ZMOtoh3yeLX2lu/LW+5SFI9P/ClZ+loHm/19gJsIFVx2
7atIQwAjxiqOFhuBLuX/0legsu4zyF9OuHZXg4kwPacV2cSl5oX2FyUa4uDjrlCKbtXZzqtb3zzX
sAseZGvjHw/7VW+l6SZMdpdLdCAAtYHd1CGU3Hev5zeu8InhrRLthUgS112g6v59t9oUQsMjIvs1
5X0HvI1lpyHSG2oIgYmtBJtAoEdWCHCyk2C60cPyhiJwzUTgZD5fiU/OndLX0DzuvKEDGiqlA3Tj
gZH4fz+8mVvCtXWpkiWJSTE4RCrdq56LpA1Q+pUaOxQ8V7j03ntAY+BpnkZv4nCBt9Ht3mZMhgjq
loZyqH1k8RY1TplaJvfD/SIc+zi1kJz8FD8pmDnabW2iEW2x0zO/DHfnWLIMxP52gmCob/MDX+W0
Zi2khCGQPj81hWraJ8NNouIHYSLtkRq2UGl14d1HTFdd/5qvQEdB1Hnc5133j5exFJLdZ6PuK9q+
jv3++fJbmm2EssYSkAQeDsur0SDngsZQ3x7UAFcfBMAMA3TLeCMJkXmhWkGCK1PKtrAFAzof/cFK
Fl/V0uNIfXRQ0VPKYLRXt38Ysg0V6Eq1QJFxrpEyB15tG+/Ks7uF7kPOqAL4+v8J6s63rAKYhx/O
kyMptbTxvxe+fphzN9QhwoNjUWaZLXs3e1lNrEo9tIN9jY3W1vB7/wmnxBkC45loxVdUFxBczg1/
8cQNobUEcc7hR+hqanFagbbSBQywM6V0HY9tHH4a0BQHkq0VUnBM9WAmcpz5CJTU8QgM2GuNFf2s
B/UMyV8ELaQbZZY+duKXZ/HwD8SRmeCmWcOwGl6yggdBmlwoebF9cz4WlchUG3MVI9oHcvr3Acie
i6L35nfNrj8BGxRrlQhL2VmbkLHu9+tdZQd+6HZd8fXy9PukH06/DRM3EE3Jh0WPZF52vZhEXPYh
x1VBLMpG3mEOAdizfQd27CIUlyqa3HVAAVxUsIxmmegu2X7P2aO/i/ZAej/m5U+XTK0yasIIQK+o
kZlz93c67U5RgSjrfomM7TBDqY3bko9xZBGLADbtYrT7Yr/8i4d8c6azoQ3oMUiCuO8VnlGqriqC
93LOtXmNijjureXiP5eqY4tgSUeTiHvJ7EF94dhfH7eQ0lVruyAYHjJ95JgIHrNEhmaFmTmN+N9f
dJrJWoqGL0ShnynQhxQQN9hfrGxWBKuq05jk7lTM791JrRbC6l5mP6Hm2SETzM72RGrAP4gC7lLC
H0PAPRngDCE4yDAYLjpoyEawNUYSYebA8vH8wY/HRx6igWUlldGPEJCh5jkwBIVo2QVQgXWEI3ve
QzOnEvQ7qxa3pfb4vdYTPglUQzVyv8vi1SthMJj0eglQbMNr43Aw/P+aGWwu0XbfBsGdZwmvT2ty
kW7VD7aIPA3pdDZC0aCs0t4GCNkHfa4FCLswNOfZkKjiHvzgFi9vj02gEB4QOj1q72S0QD9N2Lbx
3ntoiB279hKzXZ499Yu3dGNAbBxo3tsDorY2fAZXg4hjS6A/sjCx3SFtRhroLkTDBVPLaEftRgUa
L+cE7hvHvLxa50Ucee+WDyahOQmWWLJXM35ROA9fwIFiz0bAB2TM4GJA1uRlNNIp49eW7Ek6vgg+
2GBF0ZPOSEor8iNEXG4Q2lpqjEngozk49AXrAxVIbPegFAk3OdSNwPq7+3qrAaaHmqd1F5nk2r4q
dGeoIKrw2pjL2fXnlY8BbrPFet+SOn1sLuAcyvKs5X6bzkemxFLJncwK6eM5TqxUqZgUARewWtvc
Ra0ZOOJD9toe9HzM8R+ub3/jjlxb7OCfJg2SMPw6ACkHjUPwdukt7nBywCYGeSY94bA7WtNVKhtg
RGaHeyrTOj3KgDQqDn8HiNTpMt/z+ubjqVmeVC7MjtaxCFmC3PurwbTITipTxWu4RPAiY5iKPpVO
RdjaR3JDC8lxAwifhxTiU+3laJUuCrVMbfuDJmcq5ULO6UldT/lvQa7EgaCwfzHs0tQ5qzKtp/o8
nBHRFj4ihAdi7zcGSd7U8oGV1l0D1xvDZgjnv43C4YyCRo3T3nIfWua4n7d/8sqWl780LBBOfwVP
6qfSK1hMYgwGjqYR+8DF6x1fhiqke+S6cXct56rPhK/X5nOid8iDWadT2mVuTaSFdJGahIpaXcXq
ExuC6t+D/4ENQ12ns2Bxy+YdhF3J6wFtIGQr0vSI/GE3UBwz5WLnf33I7c34yUh2hhr3Kv5UavyQ
QByMhTj2UcbsVq9PktlUOL0qY3xlEWM/l7Xma7WgyDlf3LuRosajw42COuZAo2d/WL4G2n4jnWYH
IO9TDaVxNDU0SNX5Pws64s3Z8qqdqfFWH9Id5LatEgyVWI/6XjbDpVjHAKkLpnfrWYJWZUAWsP9n
jdInKehVzqm1B6lMTUrOgIfVsxTqpQ1Yi2yBDGGORINHZLzRFLWJxc7+pUr42RUxR8uQNSlxRWNk
eWoMtlNU3MSPpeBvsEHHW/UNx93MxLb8M+0G6/4+P0GOW/ZJAkLIHOPhqKkyiSl4WK3kNgLduKpl
K6jew+ZiyP3B8gk9MTD/qL//ZXpk6Hj0J9m+ZODkcUmeYCotddZUZLKnXNXsG1UIuksl+vCe4D4W
c8bA4GJi5rFbwoMIkcaFkbTPXRhK3lPanOEDbJtHEhWJkSbBMIKiZ2D2p2FO8isYICjlBEOkeCT/
a76lJ4l4gVJkaeT6qs42OPHT5HQevEKq+GM/cxbRiMfLhvKWGYSbRbmEE1d90j8m+pdlTCJUstTL
1foh5SKEIuhbjBVpByN7lMa6MibUlhJjp1Xoe2gVpEGUEpGFhJIKKbAwtcZ9fMsvjuQHRSxhFFhC
9O4kmH7xH66rcbraK9wj/iWCBm1sqSvTYcA7xAKjwb91uKFK5iYowR+iKBXcRRXeNXgWg3B2Vgmx
Fyp2mjf3RJBUYlJL7VikrPkUF2jfQNB41REonPMv/k5HWfc1kdFAZncv5mM90bid7ffvY9SM2++R
nHQJUEntFSXX8X2Qfiwqy6x2JUo7NRJLSD6eL9LpYY84G8IE/nw6Rkne+p56UVs+s5GXbd+PGibM
7+tZlizv3wvE0KK6bSZz7GQ/5IZuX3qQBFMs9hwNEhnE9N9aYXzT1JFcocuz5IHzrH7TL6UpSc9z
URpHrDCS14WL+2MGYWB1wwmrIzWekz0LGfqUmSJkHFz3tWFPIlpfT3hhCLTHzv8w/Hb6mZDpLMIe
02ajY9c3QB2UQFAEOYgMOhBV34qnuHohRs2s4YIDm2uB/EDw9BS7MDi+R1cG/mvz6FwrLgW+kz1E
9WZ1Po0Z/OBmOiUW4ZV59eR23PERQDfjC3b2Ow6HI73xt6tbiC1uIJD0KHhu5XMyYmVL8RnJ+pQa
bDxGoYvpP8oLk2IPY7jmQx0IDllQ/C4bd1l6a7I5OFjfJMKERG/MIkb3T6bK5dbRFITSEJbkEu7e
oNKBGnFfO7GhggRHUDoFTqut4omJYA6UA7A0uSfdOoR27kzQ8+KryfFl3Vp/p4rjD4tYsLUiByLG
J7diXleFIH8MN1rlq8ILdfy+I2PY0nCZk4w+WVa1JNPO611Y9S/9KZms383fO84ZJ0qU2kAnd55m
KF8EVreha/SGUadUlTZqezPeBW7hb9zJgXJ82JCJkBlJFh1oKR5UMla1Sn6xUliAM3PzthjtSFei
3abVSdFLhL8jch1zHVwbCwOWKDYz7ZRqF/hg81wsE/TLT7SdE2H/WWuGucPmMp5zZaosiVO8/1RC
AdxVrHDcsBKw/4dPBMtTyfga8B/05VWTo13yOHYeQRVK3gHQoIrrCnauUWbEYDzdq/T5/tkY4DAW
nThMxD23Oa2pAYkjSl3z5GqpAeufrgi+Hka3/jJPGAi/896APMvTefSNLSvPYuc95i+r9T9dtK6b
0MgSloNQIZdQkml7BCh7wfkLuWtw5JwGWT+3sfiX+5gQxHCcyPl+Gn4dVVnxQl50wXTRYeMC3Od2
ijhUlLE/f/5wh2kxK7r0jPQuTyi/x5NANGeg57iYr6gJQgAHef6EPqXhFqijtFGfTifr46N80eXA
0mRUeE8gzqIZBnbdmUTW+/KaezwF5b1y9bBHSQWXqhPg/xB4yYy+khpCcZjyMZ2Mn10ZAS5bZ6N+
eM+oJ1x5eSLTkHuBzXF9YZSag+ujpdhZLxrSg+qONuYic3Bd7Dn6hOPcnylRFTfjGbCBfm2XGNdU
EqcQaGqsKkGF35Au7NFSVdGrgTQsEJtkZntLNLPLz4oguc6Gg0oglsL2BB/vtEYaD6vsJJ5o7G75
qSMZoZUPgcVf+6aIul0m2OTavBdL3drjN4KeQQ5saaEv9PZtIqjY53EdAnu7cbsl9T415u4Mxq7/
7ZT+1IGkE6kNkpajt+iABg5aLvhTz/XJMzGSQJHSG0VtSF5zt8gnsMhe1474DdPbczN6yN1OQpj4
IJ4iUf1D9x5obXIuy9jCJDNSGuK2demttrfSmikwhukr7SMtDMjQYUWNZdSDyBihfwJ9wds1BpVP
xAAhXwYaI0TPNHxQIXTcWQHiepvc3U5Fc9ndUmKH/T2l15EmLVyiFyYjeZe9nwhunt33KO28Dmtk
Cbn7Q9tPMD0wJ8ivJGBESMu8mrUUWrzU2AAGKXj3NzrUV8M/l5avLOT+qxZDmoRRLM3mhQ/zB4PL
4AjyXZsbnUD7zqgNzqIVO3RkSAewFrckU+0H60lQQM6ZTIfrbITOkyo47fvurbshTK48J1fiHu7c
IDP8XvqksHOL2ENBHo+exqg+v2poSzQp0r4vTEv3xOYx7RqxiTZsRkC06eAbCbK/0WqkkZ+GcvVh
4pajWTH/6aVBjkBvUINPTPDyaCBttlpDm+2/2hXnabpXxJA6yWGfArdtxkzEgVLiSu1d2b6veQOl
j5Rj5IEnHLvM3vMWeuSOV7SXRuaS6wHfLqsNOzbo/fVElZAsHV2c9kuKUkJqAhJX1bJWFwImEANa
/bfUs/oiSp1yxb0J5zyP3qMfvzu+JQT4pR9wE0NZ6Ap8lPMZN9gJHP4nxhBayQDWxYVIcHc5EidJ
LAUyOnd6YilgalTqU4dC30C5A1QKsgF7vQf7IynDwrIOOiw6mSUKYKN/943HALvAANzNvItKonZU
WqrA4aUYSZ0uGxwYoQBIyLgdyV9UsWnAhHZ6DWTZy/fZU7tzj9bWHxxiOquQAmwx4pflJUoF+01V
YiXh+TADw6sEX+u1YoLgiOy3s7hlUDxw8Q+1vbs7w1Ivpo0yPrmkeUtEZsUUitQmoB1NFFtWhf9V
ZjQ3z/M8cwGxSr8PNrxFOiLhqsXuCVgc/XzeX4iOUQe/NiqLdCdJWckQZqNsZUOX8uFgWdta9HMz
VGlGkc11wlCUx7J20p173kNXTA9IJyzi+RkA1i1zQbkOhTZchE0LpDwPJeGhbOTjcyC0KhW/cD4l
t7hLx7v0rrr7yilxm8oPoDc/PPNMB7iacUVp63m9ZEvtQQMomljOCJtaFWzo0J4G0eIBMZpmxKFJ
BM3SQRjr0aX6mtnFF7Aok6undJ2LKx/ypVLHvk7uJRj8u1JbybhYD6RMuBNc1ScdxIpv8EQeqb7l
wVMHAk8xObdBN6tAngqEz9xG6QhEpiMaTI3/tjDI3Ij3KXVGsgcJ2NtwBivJPkVDkOaIf4WjfMgR
wP0JdIC4RKI+EsnNQo8YKnqHUrTOyvCoVAacWXuLinDlHLi5au/27o9tOXKITDQBq8lzYV3jqNi2
SAhJLXyw+4hmpPLkFjhkKKKuIz1XvGdWXV81mlOvB/MikCaXMJXj3epIqQX7OSX3N3pmBxscueqC
C5u2C0qugZfZVWcKsTBdgSZCQRQyZ7BTlVcIL7RdPkJULrb2zAbST/ELAqAdgiFcuPfzQCb4a/kr
af1rg/meGANsGsftlyYmqGWZZvyXEt4dSkgbRQIwyOKIXt0nDVpWDCYjROs3IinRYA296KLzdj1m
MgiZL5Eg+dWs4kdPGKRNpQKflSmG5Q9xxsNZCd+Q4gGg1paNeR/XCOZ/BWZq9QKDGNmScum2tzc9
OeNcEYUCP1Zq0C4vnuIetgoKwBsFXCLv32fs3QGA6JkdW4OYfTHBw07b6myWehbvO+n8GTS2nT7G
/0dqsQzWlB24Q5WLGU7/jP4xih0+EVTpbpkUiAS+eWorVCmVFZ0tSP0/sDKpp5EShpXR+NjUl+dA
N+fytBiMqfoAXCuNy+ZDK4CL4wlEZnyp1g70NBeF5QzFr1QW0jxDny9XT+3v508/cjwJbbXKXR2A
R2DSYI25AfwLZD30cPNLRwLo8M2T/pMRK3y6XhtupQBs/XDbY/xB+ksRkz3cMrdU+qRn4k2WgZbF
gslFc7q5vTfcUHGwhJxyfv89KMj3t45Ki230+tsRBfGaFp4Pk1YQ65SCuEau2V2A3lIqWUF9aifY
YWNGMkeJGQQxQZhA2Pa1KGJf3oLa3vE0wDYwPVl8lW/p0vqu8QFOYKOMH+42EcssLyfkJ/XLTFhs
U3HdBhXtTdONRkSCxzFnntupowkwXccJDX1xuBSX4x0Hlb2IWPKjUtpnWyO2Xza2NLYyPjSJIGV7
U9M1/I9DBvoSDNQzImRWfChfs80UOVq2PptjfISkJnvd20rHuwp8HXiJab+rk3wRjl08Sv17HSeg
1wQF/Et+6J9wqBFip91LZ6noigVaFAoqy9AEfmmhDjSTrIFtr21YMSpU3LIJtu17ElXaa1Nnc2yt
Xxf8CT0ftu4BTa5obhFcNiaS3ZxdCaDE3XTssz7E5hX1vHhtnImt26uaV75jESrnfm4r3RvmzNcv
eJUyTH7vYR2VAe+aN7wRCBSUrrvUjdSo4jfsGIUOU5/LIuomnwTucsDPXmV3FoiAfGNSr4dUL6oP
VN7UmG3KPECEGnd4l2tX+cgXA0S9ZKFEF/rvBi2s8FexnVdCo84u6akVLeWtbopzz1I9Mg4A/3Pk
kHhTbMocZXEkUM66LQ8up3x9E3W5qW6y8ahaLgcM8vwUFT2zkCqQGCZmhhhR0WqegioRJ+UhfpT2
wWh2RQxfgBjO8e31tJIX+Oz659ti7RV5tkJd5vVeM3Yhbtd1V0aS1qPt58gu3JFxGzjr1vaqKw3D
wDzm9dq9bAA13SxEnO8iDVmKiUKlsapGWQh0IhVLk1Oa3PFKa1xayqAhv4/gYV/Fj4Esgi7DJJqw
1qO4x1hONAzVg6mMNcvdilKg5igZmLu0VM+7aKGH1eGKi2XLHxggpD6CiA3gbgocSkqoxn8CTycm
SIBJhmAQlGnikAO1A2uyljxXc/Du4dui3eNbXYNjHplyhigRdiApXegkuNOTqZWrjPZEA3wOzGHx
S9U1lfYuINnMiad6IjxjO8LDTjSjyaJcoPViztWhCcZuJgq5vBMCN8pHWfacgaYkuQUYHCecLIih
qZmUmODs/TkGWMd7jJXDTYVkzSXi/MFNTn5IVxstqG8uBTeboX1WJSgzSvL4HvJUDcETGMiy0aE5
fWPMETVLmJqlfekYlK9iDDc86kxCPfs15POR8HGkiuJMLG5ryjI+tyy+j5M/MiTmdBXe8zjflhDY
Juaxx10u3aZMRt1QVi0Pe8bZi9VDhecTb7BOiFU/qtPaswA3/4VwdDG/luInbdScM/WsoioYgg9Z
GRyo8a8l06oqKptN17upcfe0iXU92K8rLJL4i8kO1aaz372sM4mLOWrUJP8Sr2IYPSxjXXI5mw4X
fVO+CdgV8Q/P5iq7JNPdHh4c2C/RhNAC1xIOSLH9UDYtSc7O8nkhbdfF4c9+QviagsWJSQDnWAyH
DC3zvO9JgaEb2rzQGThs5SovNCoAKsnTForoxj0fDeF5fB+cTK298t0HXKnlS9WCmbfRyxcwtSyc
2XiIBVD0QeDWXqWA75hNImhpmhv5aZrq4Xou8fbrylIKiePmLLTucdBnF6LoRoBlDDkSOrxiU+h0
gX8lRGbcz9iAmPd7Zs3o6at1yRb1BwAu8PPUeLnMTjJgajjbZzuKk+Qf9ruH6534/GGRePv4tQaT
QZhm5RqthDDh/I9p6luCyUJ0pHd+djkeYyOKJnMuQic+OBAENsHTKostTyOWfJsfJBKTbdeIvZer
LJlJRpb+az/NRK9GSE/3M34M9MwlSEAiCfb/mUdObbQOqIRp4ZKlb5uPbliKxDOCTG9ETJi7qbEX
grKf58iDY9LInlQD8/nVhYhh7iuKnkUOknIPl878+ONuW66443kx4fmcz4wKt+8qYRftZxS5d/3p
ERRM8u9421MWP77QpmQx6mh3r4PLxA3wXK/HpaWNVm25oSnUeZRMaLqmgvLSSUSeQl5tlE6kcTc0
hsYeWLekS8JSsH2t3XldVWtKf7HO6wErRMAp4lgh6rUa9ugGfKlgWYp2nfGJlsLj+I0EyDcavNXh
ZJHx0MomcjPPb8LTvTq6HXiHASP8zoDvbAP9vgqVs4W9mD/SXqKs299ZyUPV4f/mAWce+MByxF56
bhzxSL04dE1yu5MbN9dQKLNJyxqu+uYZSPRKzoDH4cMY/Cz/nzrBUZ/Up8kt55LaTMcaHPAM9A2O
KYydJcM/oaRn4Qr2HRe3THK1nQl2ex4yEDAuIxxTU1OiuOZAD1vF4ATEFH2cQUiqI3uKLqOmchXM
M63BBRBeJGv++SxSsij/4BeVebkl+NI0MF7r91sMCfyv6QEp1RDDeFdH4Hb2zOvunpRnizXQJ6E0
INXVqGwzmSnf2FV4IlNEROwy1ECwg/DXaGh7ce5ysVjViKTkCzrZ1xJ6oVaKJaQ4cVFeA+/SF3tc
wRElMwmgGt4fcQ9Da1AflbJcUPmRxZ2sOtw+E1nMS5QTAaGp95qbNM+SsCN23suVd+VHCcMMuBQa
quXlM15k/UHZiP8xcn4UCFgChc6hxliJCN3tHJHRgOjK0ZDiYrgHzt8+Y4gfGPIqb5SB/warlDhZ
l291VurvgmdCfeFcplMOEgGS1xr97u/W2lp283c/uoGjJyAc3pBVab8uqe9MPiy5ntAVf31n0mGf
DIYyVCigvTkVu6BHZx9l1/ehXgA+jhAjkCR7RIA86zO/9kFguH7t7nd7v8C1kB7Udci6xg95OXzN
OnZr6saqCB/+VIx+nVfns+BhVV1RiCP7s51WZVjJkCiYyZ464ACuhbDeeqhIkTw8liEhypZYH/ny
Mb2r3Y4CwNC49Cxz4L4rWZd72hgj/58CgQdUdeRhNpasWCfrF6tP+/poeNklCc3+gFP7CNT05mGl
SNQsPnQAUX1jmhA9U3HJGJnX+7q3uKahxpYvYgPfOLxGCwqA6SRrYG1GtmIApAhxhU9J00GRfEL7
6a/fGiSXD+ppjygR7RgOQ+GonqD0pqVJIJW+0RAE0wYGhENw8uqCHuCQ97uYV1SVwHf9gXh2251O
k48h2/FPq9IHgZ8RWKE5yYAyoYl57X2li+KCk0aWgHfGUp0wwXbgD7OY9+QrEum/tWiwCh8L841c
57XgM+sHSnN3WKzVGXeer4tGntj0qtLaWWFIggW00jTrAkT1eDQOw5XtgbXgQBS/axn7b2BUxLRg
KAQuGFsULdBXD/lDkroRqIPwPFJI+ItD8m4nlZ7qFh39W9aGrNYSwua5qRQ8gFBUq8MRuOdvbIim
OI5sRwlLOrJjtdr9gvkq5BtYVwXHOAIC8fJPye+RueMD54IwCIYzhmzoSi/GbyvwjKAu3i3pqwnS
rja6z3Kks1msvuYivPxQZF0Lc9xHL0hDenpwrEkCKtoqvkP/dIlmRTkpS4yjdwct0DEr+a2uoGDZ
+tgbuaXvOo1k9/7r87U6DnkSO+KffRc7LR2RVQ9SGk1YOsMsGhGVSUh2zxkk2pfwTRwqHVpEoHyq
pYFFXl1STcAtswOlQOQ6mrGDVpI+OL/a18V8zjF16nqK8ZbvFP8+ozu/oHPHjOdTtVROT1HPIVzz
M2W3BirKFPtKC1/2SjRwefAZg/tOjZ4PGRuvQgpJkNvc89v8LtGgixvSRqPOlT+UM7snweCN+Loc
UMQMDFBjmqOj9IKCYMnAZBAKoe+PWRviJO7jKAF6wSg5lQ+CLPLv7uwX0/kiYukphYZHz0ZgvmE8
q8z5uqTQeuGRZzjEZPdSd9sX/JFyMtHX8AQaWfckT7ohXgiE8NgpmfXVqUM+NWqaMJhMjdxWNU2k
QotzMCIFiqWPkifkNMtMfU9KbzDnUsjpVEuWA3ePX2LyujNd6nW57LECFUQY2EaJVIXwUyl1Hle2
NpcHHhJVO66ON8byn1z3b8vnlW0n2WYbwnhd2i1gT+gxeppe6An2lQkaoROBbBMZKa3CBJfK3PPS
0cv+95ykBfh6rD2YYQ9L8cyj47BI570f5PtiK0KwJspDy9KQ6cZ7s25Ib1GF0Mt/WSI1+BiPzA/4
HCRr2S8XP89gYBDeAU94YXeTb6buHb5tDVYoXtEcmemR7hZ7ksVLbgXMOzLz44nrH/pYYTUG1fxV
hE0eXWhw+gHoaPQ3PD6yIYZ9/DqWWGO9TcYnAjiAZjC33P3c+vWSVpiyPikWCc2+sTWNLGGKi8nd
j0qlGTs2jjJQ/GqHTTh/vRAPFyP9PrR/QQG8YaREqmdchzZc54vfYKsO99jnziF7PSiKJJo4A/Uv
5hKmzCB07p8WOoIcrZxl/t+CvwwUYd0KsbC2PMsk1RRyZMUzN1qb3R/JxhLBruYtvg5BgsNnxdYP
Kz4HtwKXaklfjxGR29xheUcenxadsEdDxj2tRN/wllFpZyAg4/1B7+LhAE0Og2rmCjaWnHWS4mCm
9Ka/m/l+25pxyAaqQGov83jGQpLuXyit4CsuQB1CgTwEzGtJvlZG4DyozcthFoiPiPtm94ob0i0n
h7GqCPc8EfpKlJbudM92Vyqo2mteW1D1PQaDdnZYw3NSzEiApkwuopiDpGLgjIKb07h7Uud1ClWt
Tq1t6R6SYSlgoSMGw0kIkgNcWz/enGEgD4FHSu6FDybMgtmRpHCZYAP7WvfhUomliyUwDzXOpF4V
Q9Us5Sje/H5GG+xGYiPbjO8zHI0RcaYJcp2OsmuTP2zo5G36/b02wsgDlVyXRcY3dN89rk7lWFMA
ITSG8sKxku/sYQk6DmKjPPPaBfFdUyJDKqeuxTky5dsarOua/eB1U5eec1WjghX9so5TAKjFxlWd
C/0zXcSbuejglHLGSAR13ilVpJGdV8iYMSfGpSG2hSkqLOiZ0FVCpbM2hAfmNUiUvDJLZshE36VK
UFbtWABTbyXUHyHVpErCl14TB/tdGqvSDgpUdmgaEIlfyixKSVRAx4wvTcYucq3cVBABaGEEgXk3
vlrNz4zhhk41m2Sw2KdyV5LHOhkzztAe0E1QOQ4lXqlwZhlqq9fm3BhwU0ZHQDtAsRCArUK8td3j
Y2lORBQf7HGj3Qi2p/Zyo9mt3Uz5p4SwFcTh0ITUD9bqdGyePGSzLZNgGEqUT6KBeZn22XG4R9To
TE/cpplKvonMm+XoMWgyAxIWXBNaN4ZM7ju3NcoiBsgrDoPaAbWV1QODwuP3wDn1UNG8tZha6e1J
gcUW/30YkX1uCG9FXtTRzetKdKYsgPBrl6xmkCgU+GqUmZquBqyqYC98vcBaDyJVCeagf0Uhlj5B
RWnsml8v0vFM1KEJsmJaS5isrMJd1/ryGDKm2TaUEj6gp3cMAn15yO4FQr0BNE4AvoEIfMzsSFqJ
gdwYSunnQyWEPHOx/VA4aLY+6oy1wtdvzJ1gX8g+GrbYhiSOROnfLkYZTnd7pcUDBdKNxtaPTBFB
BWjtAN50UJS4ZyMQH6fcnYlxAmzcGD+zvEKXCjmpo00KWrpemwUquppqxOfgHlEDdMCIYAwXRWuB
5lnKHa/3W61ZZ+ZD1NeJ8uw2BA6lRDzw9tgcgLmueJoZ0gzE3LZUKiN1DjU8TcHGL/PedCd4LSgC
17nCB4qAGBJxOQ7GNUhQVAHL8DXNkrrlOy3KJwsNaEt0zdtd1vd6T9ig6jXtOiUAqKK0pOyLh8hD
9ZvslNj/8GvKe8G5lBXjvoo+doxikNgUTy+MPK4AEVtdHfNMuL06Zm0Gz43o24id4abvMquKDwOL
VLIyuEVbowsSSsch5nTVhmAD5OE02SCt+QeGXfMcx7HvwUliI5MbHLQ3ysuNNb8TByoFhb9gIkr2
0Ej6WQLSEZdchwg1TPLyoodik20fsvJlNl/kD/54hktZWMUXls3Vv4tvTEqlZQb51lYvk5c/U3Eo
k8+OLJFCwjoTXHWdADPzBlPD59fr6aFRQ6rvCiQoFXksZOqSh43239AAKuo6nysPFcjYgHTWAe18
85rx04ctqG//NF5TJyrB0eXcopYbOs8fgaa6DI0DzHUWZB6EEmhUzR7/6ZbgEL0u2PjR2hakc/y7
kgE8/8jl8uKKEBCRU8tlmzZ/OIik6myU6SklwQfZckdns3rGd7VeogtWl67NMfcHezH3earSrnT9
uPzCHfOkKs2Kt+ByQYPpwY+s+RcQs4+9cZNYdZzinF31McIb0XHXBqj5D2IOO+ebAwet5nQEIqQY
bbU5YJyD/Diu9jHXC0y0gSJSAw0KvVyEE3gdxDT/CKiI50bIMw4QKVqoY8aaOqJA28Our8sPHaXA
kdtCtvey0IG15QjjN/EdQtdFTUNBbFiG+AdNlekCOzjepbX973DEDvRtarf2PR1MhsBu+H7Ywzaj
myoaMDjo/xnUrtBcr0J6im+plob8D0oyGxhKCg5tZy9iOOsb9x0CXgwFScALjRztHcEZVp8jnIjM
z6nzFazrDYbxVkB8Gb1Onrv2Ig3Y3gcCy6+73K54POZbbpS06jNMzXMlz3Fez9QTe2AoP7sgf/Ui
tVICSkMHpg7CpUqri9d/cKfFBkMEhFaP2ZMh1ZcqBaCcxOGNuaYwOzLVYct4/FqrwiVXJQqH3vRH
n9TxZBrmHwQYBTTd48ShU6yLRE3wCEih5z3jAj5Bn2oug4o1rI73yBD/8ycYcrXNhK33whx1A0kQ
WmOPzDG2fL76aaIUaWtsJJI8ZwMMHP0LbMcYmn7ekAONZ+PcE3qYoaI5OK/dyKFbw3kSCkZi38BA
18oMqtK4ZgdNuO9wA0Y7O8JPOKm7eDmnk6TbFjzkVpbIH6WwKXEhuUVsy48TpekE0hLBPJNjhy9A
vVKmomGs6orOwtaafSbe8BDANrOIWzlpGZhT+ZkkzRFht/BohwzI7gxAwhFyGs6z147C3Xgmpxkq
yvQc9bIpARmhdtj6HoNeZROa+S2tW8Ew6NBExgNoHLqSfXw1c6okcdcK+fJAZfUYkrEMvgE4YzuO
eEK+Krp5AxBJ6pEvsn5qa22DNBriGQcweTF/TCeZSrjtj2x639WzgLLHDkkX7QMULtHj22Q/EtxE
ItWTjYueYLo8e0A5FZaaHRoUP3z5wyhvkaT5JyBI7pv2nfNNoIWeoqpxaCsWS665KUDPpoYDDoTk
6dFwIMuH5UTD9UzbR1Ll57JIIaAqKVFYvvPMnYnZfTqsm86pNwWzObBcAy9Pj3Qc8jwxU0DikaUr
ncr0bp8wLIPqtzRBhxh6KZj9+uUrrpgkkHks8CFquT6xwDmsV3vnjbHZ1kqrpGoymGbWVdMvzlZ0
/S6vA2Pfzj/dwugrVWw+0FZQfXu7M9GckUJXIpruZqM30lLmDFfASRT2Dr5+sqbOuegCksQ8pzIP
puQXjv2UtmlF1Lp/gTlNm9y1x6Cr2dsJ7wwhHP7GwrA+V22vQtN1mBPsF0R43ykr28RwooBpaSH+
uNm2IyDh50pEOjmNXRvG9UZ/oh3diActf2+EASXfCL2cTh6xe5Mw4/t9YEx2Ng4nZIV9gucMrxhG
wqQfOYBSNWO2IELWYh91rBQvHHWRGJNbIvWvEfCrSTnXxSlmyfY/94wdv/Yior7YbT2Jz3pOZS3P
iUtD0qONCeZKrplIzzVX4OaPYfGTMPMSP5eoJiSqIlobjdW/o7TBDH1x8Loc5/RwrOqE/Sb06D6i
/phSsje390yuobiVUb8RXPssrQyT+TyhLz98vQC/y8as63ckVk2y6KxYiCY4Qk/LYNWSH9khqru5
d38bnG2/1VoVfcA4yeU1clUKoNVUlZTt7w9yUXD2nvDf1WcfTSxfrebzeKlj2rwk4HxAi58M8LC6
eO7jz6z3KVVtuBnJmtr09L8IGlZjDSJE/Av7vqVhWmRXHEFhIHdh1CTSSCSfOOB+Wjy2+ZioSdzY
DEwjHqlZY+qNBZXrGHtD3jqpUq1EOhnFjQN546DOeSDN818oY50LDbPOF/LnsqZJZMYNiFKtceoz
sRstNp1dqa4UgJQSImLMNdNuEfDpf97gtOh19d3oRzQyUQzxkQUdXF1BtWZ6483QW5kOzhXYlM5m
2BlsCD7NAkkzyBt5hvadkbgNLjUiAW6EU/CkiLAWjTw1Lpqt+tzRrTb4kiFvgkC+Nc4nPV330ANi
F9+J2NwY/JeJ9hV9Td8KQB0yaUTOrQvJBkyUj18+t51dr1Rss1ST3TpU4h6IjBewH02+6EY+hzQ/
EE9pmKnDyeRHHRmi7cdnmMMgNPEyzKUzf4grquCYifmeV9C9uAlBuN+2FYxNu4wjbwPO5ccyodtp
/53RAm5a+K7ZI78TjG3cAG8C8QXpHi0FhwWnYV4kpXNZ0XXK3NULPwkPENfh1beVz/Xz6oUw84KT
Z1BlVkWiPViMp4Sb8HkbGqj8/91m7lGdjVUJBNPq3vvgFVj9mjJaCXsNG2Q9LCH+6kW2Z1DCyTpJ
xEg2hugLX6/i6zIfdRquD0CCu29HVoe5UYjic0oXWi4inEdEoFC5XxwVnaZ3RxrMZkOnWXRN5T+6
3tK3HTC7PVZ1Jjh0eNzc6BhyqDH7/ecH+POvCHcvjwc1uTs5wXb9OYVbwO8vJmnHS9ZOVIfOLtK0
dR66O1LaOi50wz60c5CYZOBZV7qrbNvP7xn1KlLqJI1ridc/ui+2LZ5+la2cRI/gt6F6KgYxV7SZ
wN9IOQI4OsdxNk+cDY07bRBFqgUBB2vB4QnCzGAeTxKoDgtcv4QNT7GOnH6UDNuTB+EJeRRQxvLp
M5xYhR6DFFGNJ6gGLAJA5yUQjoNDS1U9tJzU2/CXOh4yv3dguAuERpjftvd72Y21W3qMxZl6g18M
jpAoxFqNMTRHXUn8dRebWe9fo+BzR8++ur8JQzbV9RLX5nzAFVtiwQxbt2YF3oaOJaoXtHuflFla
XMYHAiI8iYm3OtGpLmr29cDLzkAQOmnhBZq8iANHIxGGhu1TtHfPwvF6o6friNQOgHrcVQPOBDpa
Qg7cPaPFLXd7M8yy0A3iPAWDCrB1bi/6PeMnmEHv6rscnvzqIHdERjX5oSOWnSIngV58WHtYTvWC
rbQDXAhdzkJu/sfgg+oU/K6LYak3iJs7YW4zITPc3QY5Wvqp0NVYmy+zkeBuK/ndfdZbEX5N6ezl
szMqSkKkQpPG/vwd4VRL2RWan2mOqZHwNhhqvdsHLIfED3X3kEGy3SnJs4gUhV9XiMbYPldJl9re
UTTJR14/CEUoczhDi4jCxVtPTnWNMD4Ihebr3bSnNNtFZ9BQkMHLneUgPpopaxDMPfskkjrW6apZ
m3fAX7ZCRF6n0MD1BIZ95jHNfrNqF0HT5ss/7a5fOUhPCjo52E07PId2NIZyDFc93+XTXvwFLzLL
AJO/xB2bUKRYpTJlWMWoLpks8ChPGBK4PiyOFi3fhHnJMyKQIcyrH0B9qzkmE/dDC2/MAC0c6gRq
N992PpEtnR1S8G7XU1W/W4e7Upae5I/z2ajiw+2DtkotbWH5Kfr3kapWXSrvDuENNJTq1WsdffsM
A0EQu+Dk/zloXvvNtX0olgkg7QUBmo/N/ppK/TNgXEV96gqHDixUv/EcuOfXTVXTDoBqksKM6sqk
iSqUZQ97HCQ8UmTyp5VPE+pasFRTY+oVrU3d+Dhl8Olx3FthdSeP61IMb/XoP/yD/v16xA7kekxS
ubuLIy4Ato3znY8AE3dc6FQw7xYElpiBDwwDRTrVYzAMawwqOLdNqwrAD6Uc7DFwUkU4sz3Cd4nj
7fwXMs8Eh1DknzdEVRDJRiI5kDADjlA31kbdASAmhGdlZ3BmpIXQ/vqYf9YVk1LmvXXkoiLPwVQC
AeCcdviKs1D56fppZHGnrN+gGPUzgwc9RwwzKISZIknbEZ8ebkZwiPYO6mzDXrFJRnlhFjloHyEF
lqhGt+Wm27zeBNbbds8BUiMd+YYB0MR0pO5gf6L4JpoGuPgnMXaR2pMNix9s4OKBuwrFoBuwCknc
1yWwddiZv9G3ZS3v6P6xjXllAlBx/BVZxEo34UDPpMSJ/ype+RtzX8t4JfeGifFFZzA8Fbn5v0dc
kqNHwMTtSYi6svOdydohFkMgoPzCEHbT04X863zUrj7gSptSmPlTWXjqmCOQc4UZnedvyp2ypD35
sJFDLn8uGdBs46XXPXz5Ol9iY5Hxuy0LzBxIHUO8PlJMMaHXvdrFT7uuEPdj6ugFwQyvN6ad+p/5
v1Sim9E5dQ6rpcg0LMzQRpsforyf/+4ySoKQL43tuPO6gxhoYyfmfea7Ag2PhHLCC0s9mtGx3LVi
wS3HP8CIwSKNjpT9j9+URtcw5Uz+pqxSz8nvmqTB7O4vbED+0frN7IXZqUw1Cdr5LKfimfXS8R8P
OYHVqN6nFiN9ONC+hNSZHz2Eg8wLUmGUSVuGHxmR/AL1HabfFivd2Xh8Y07IK81lGOr57WRIrUm7
S3U5HXdldq0NB0YiO4aqDeHtgNcbZlWASX3TOuQUA8EtjFRW0P8VqX1Reu7h49larwlAPssMBad1
N0GTD4br7AUaChs1HBHXbcuiP0t4hCA/In7GJGSxopW60/q27eHd9OEYDMeJdJO7YTR2C7m8cDmj
ZhZ41/E0YpEiK57uZuXdu65U3G1Q27GKNuoCmSj5mfzwI58ctcoH27DRD3vDLPMpHQD0XCrTvgB/
AHBwoh1TGZMI9qlhz0bhuxmiATrKWTPTOTn0NDpI9Iuw7t+UBVDrualeWqkYlLdwQAljs2Sc/nmO
EjqkEFBzKu0HhGv5qVIL+z/RD597tGHg9/zegewhHex9Md/llYM+/Ae6NbTCUnp4/vJ1hU2zhT42
U2IqOl+FvNpMHQfpqCNgJ5ykg0E3l+Ld/93aUZD4Lisu1GZHBoDNxEPGDjXrVsw7Y+LbbMatK66G
O476ZClpLtyMCKXeBrn4T9E5bfTQ5OWaEmwsPIZdFyf4uLZ8EblLk5n32/5VvI+zCSFKSAHs6Qsr
4ljcdUclV4d8BxoCvSBChhLijMw9XJVe1SpB3aQir6xRDe78un72yCVSKAwHkBsJUC4zNJSlnWtQ
FA45JLoQf8HWm+B2pOrjE4vBOSnCvg5w39+8moJIPCykeqvqaYLvb77Xw2rPs9+Jhurg31ogi7U7
gzHoaKZSoRoXYh2/TSnsGh2QaUQIreST9pi6Lz6dw4R6vX5SEqe2ZG7upa8Btbc/1wutpglijM6A
0i0Z8OnBAKytBjowozyxN1DWvd7cDVCrKEw8zLOqwgl5NY+phwfvlYRsktWFNdYABzRzB/zIUMnQ
ky16upoc7FWPV06FyqU8xXBcrXt8Bl5WmwWtx5oXmm3OeBJMH5ygXJPJiLYvOf+BBtquap3YTuTd
ShefCOHGDi18jDIbM32bv2+tjbaVvtG4rbN5wqGmRNSZRaj9oZ6ZkjJX2SsCBve41eqBDPotdete
ocC5Ojq3Fua5MfqiWYAriYU0QepO43dsmoiZMNqg4LjfJ3DSvhUE4xGH3kTQHRJ1EURimNhoMNul
CIHKqJPYVAteVQ+Oj39IzKs3yyFRO5C0CzNBNd9Gthc3cxwx+xz01ALggVTxmIY1WRDZ/aV4cXvY
KrFe7qn8eX6ebN9prxpf+fu/vFhhjN1DT0rLVFNqQQjopDrcAFSJRVEIcDkFFG4IHQFh0AqB9+ie
w5bBBMiE8d/QgNhQ6WSheOe3/yIhS5le/hdvWfUlZkfUKLSxA+mv7KRDdty7ca+VKqYspAQQaK9N
7/b2AwMyHuVJDxz952GiO8cgubpduQPHrRg6kwjoopNKyUCtA3k1jX1ROiCrryGhiO8ro3j9nAlD
+ZcA+Keu8ruL7jdxMPPNaR9EYLTzdUj99Dfqnw2URftW3j5tZskwXTEo40pLHAi3bcRyrJCS8Nin
Lio/s8lqR3ABa0QBbzRoP3e6CxbOPlFU9yTVw2YIFlkrOry9pIk8gN4kQmAHx1/qvai5qcMtjjOC
WwHdkd7LfNN4lUtzCdmlPLWRGM+VGAdM8akj3Vj7RxKYzC4Aw3y4ZocS/9qOhgIQYN4kYrCBu7g0
33pgo53rF6Cze/V+zRsgZhFZENEAo3zSLULLOAlEOh8GGeCFMLF4Ed6et8cfFJPQk44q8oXk7Ets
0xlQ7GrSCEUtM9nZhQ6NmW0FfQ6GgMtrNiTwNYh8tFH2TCu/NR4WMfykJUxYEi0VtB/91Iy39osT
UI1mRc6VhrAWHfbDviRpiawnX9qmpnazswYY9V+ubntEO8Q4uK4q4BWy/FWA2YKRP7g5JA5G7fJP
+Q6JGFIYFm0D+UYGf265RvDF7zW8ADMptlpiqO2juiGZd3HAgAXhNFlXrRnNnDwP7eUap52cw4Nf
FoP/w2mu7JiUOJVXnHPVvb+8Ou73gurD6sne1h7K7ubSOtfRc8+6HSYqhezz3yjeTzXbjwbtmjU8
71BPzaMHU7NPdTCgUxqvhw+pOWdQh2HrbZpRAllX2UQ/27t3fV5L1FZgj4XjJY/HJSsat905AN7b
lB6+Cl2rXr7jv4ghoQvRZpppJMDXQqULPWbdcQ+Wjzq9s9LXHpztV7FwNjwdfWRvMdfXC+VRqWpf
B93JjlsWSt2qGnAHxItUIgoJFOkOjYz5F6tbHn9QBKdHLI8HxnkBmEZoBVU7hX0akhiX+1JzWBdU
ejqIjlKBjrmPdFBkVs3sh63CtLHbhzY3P3S4HOcDqi4gZRsigrwZ/bl8E3GjasNcyBa0z5UwVbEJ
ztjGRQWH+Njf7kUszqt8z9TEbvlUcu+LaecZCZg5viC+giJhHvdXUXbVEN+AE8MXT6SPO3iaKbgc
l25ZBA8k+5zzyoIgp0FO6F6nJJSYo8F6MWiEKCTJ0E6GvC0tYssaXm1I63gh88q103bFzVKtLWNr
eHFkdsvukJLKJBujwkpItNLkDDoAYSmiB8Rdhbec8IFzem4Q2it9N5MkGRaJfZFtmyiI6lnU9r+i
PlXeWcd10rb5H7q+w+YWkq5TdiU2/FpbzSM/1VVK4BwwDP7ykjozAmU3nUOlg7ilAJPvAym4HKnL
Sh7o3VG/1M0aZZ0u1sX+5bONgmH04ouxrsz08G83QQ0/3Z7+FqBMXm0EjuoLnZqtZJE8Y2KrNXAZ
Q+FbeRHmJUX+aGGaEtfdo/ECOcVDWmo0RfeUAnz1VrlPLbDR97UMP0j3k0wzeSi0PAiGSxnzp7mm
EiVJNnYTjkMtAHv89AC0gHsAcdooRQ1SscrVyBJgiMnC6VigxbN4ADme8qks9R9eKMNK7clnijyO
+WvFreJhUPBecLUgoCBHaxE60ygmryOgPjdRCbMphPvgGULc9Bb5EzNt8LuwMHWfIhd+1Uxkttl1
uhbN7XqS4yMuEt+Qt11Wyqba62sZkoP7j0hPuNerLgoIJGK8Q25203Lo3QLVdPuRY81polyNCMsp
1cacGXsvJElOwMES8S6Z9JWuCwU8esbb0g2e9rIPbUeXEfa+KiKWtfFodbfTGOz7HJzKNlM6aHAn
FZO/hG5oPwDSgWGpG/68l8zsl+w/U6WIFaElxLkcaeEneLx50aq3xW5YxNVcRfyJMgF21MQnSAED
JcXX3+AofrcocgYoepDjG9TwZrD0+ncVMXl0xEmelLnHo2NrViunXiVGUgRwCMdMMwPRZ/ZAb275
M6XiMVTFV5l5Ur0WI/OeaaBavWQjWPB0PKvHe08sCtZqbaqxauPp/FQpRy81ld7ZGZbM3EhExFsR
G5u05Jb4aGiVXGUVxsKGgdJmMVda/xwqPleoMJWFjUn9J3P3UDanTZtygfA6DhgSyf7trog+5PZA
/UTr7OCCtV5a7RptQbO2X9WbfWfKyKuhLHCbm8HyPd29XblVspqeSLEM063Vh5qF+qUx7IFK6//I
shZRrgfG+ikQrs9Goj7+PzHgUw/xAuuAiApCaU3tTe+dyFQUbfxqhgS4J7/sgclezAPPDT0uuhHR
fOMYX+0S9gb0qPlX29CTgnOTwVxReK5a5HiP46AIY+pCFLp1NLmbwZOgrgZzfmHsN6BB6DCtuPu7
Kl6SjDkCTVISjUYpE0QX5M8WDR1LsWsfCyPwifOFDsrUYbefkBtN72+jnNFkkJjXXCgGnpibvmcs
eblUyKFfl/ghlB95Onz2MPxpnFgXgutVxNbRYGzbtBN91DEtLdg00fttk1gciyyL0mj334doAUv9
DivWIGikMStziSE6BYC169DKWlV03vbQ3X+Egt6N87RKLIpwPKjn+2Onx49ws37lFEpDCRn98MaO
gJdOT2SVI4eS2jGFsD3XJMwQS0WzTvAj7y4ZoYH/uo40OqozOOm2gzM20Czv9OMw4IDVAVyATlaz
uFPv/VGCAMZJJqnMxkMJKE/1N6/Jd4ue955iIdv0rOf+nHMvNuB2wvgzS+wubDCTixcXG5ZzPG24
2UrZkJtqGr2QcC9rw2pH5ELLsDFkx09sE7mOvuO9AF1fpR4fvJcZQVftbqTK3wzcZXVfj75MBUBt
R2quyLCOy17+E050jAB39om0L7DrcMZE5SsSt7o/Adxkax8RSU60tCKFDB8jv9VFeR+//gfkuheq
BfkD+tqZ5ZCz+GQlRWTQh7KsP96zDD1B1yn4ZIdlO/6ej5dAlr66WOtz/micE+52Ydv08QV+QzhH
TKvKlYSAgIvoc2IRFEFCITbZo4QmLN0M8JAssu8H8nGnN3iY4PX60UZIm6HwQ8cDSG/Rl2XDyJ6o
D00MpdNAfRE02ybUeGN0OXCaOmKGNfmtXZ5hizaPf/660BqlQwWe4fbviJObQldVQplvHcucpYf2
nIYvc506D3dpiqnFrXaaIcCoe51CMrvIpQhYm5j0Ow12HsvfuEAjFOZnKKlZ2BQ/5nVpnRn6D8U8
QQ33NzcRsNOmtY8RPu6HqhvnulIbVUZ6eaEnXJHcRMznfsgFESZjjzhsiRPewxXIw++/VnNg+ELi
hZ0TTg/NC4THs4h5LfX06cooTdmhcavkfCN356Rymc/fPnnU5QKcGE+lK+VdX+NUuuiWjsQQmurH
ay47s3LnOu2SFbIErLzpCpxNKpCtD/iP6AFOEDh1vxepPn7Ud3PX9fo5oifsvUz3D682PWJ/9PkM
00xzdq26Eo+vv3CX4ePlJZBKG/YK3qPvifZSeTwiBBnAgXTmLJf539TxgzLBQeEiJT555oEzSVx/
p+Y+hDZIkJAZVRr7uiPeIdD3DiQuph+AKSOrpzeybu2P6HPMWbL3F1KD7mTXwqGf5LlZaX9ifoKy
TbR/cVjsvO3C3mr8JXI86v35BqifxIryP0c1VzQQ7h/XbCGnCfdny/AfNlEhJrdQrfxqNdPlm8d1
cdNYZxcyD06xTvRdD6or7jmmjtGCnrT7rE2u1AQtd6ZQZb67Yi87idL81t+9n+tAfT+qgE8rgxtb
OAnK3tbcHukvWa0yCfrZ4cFutw2/l3XQzBAnYl03rGyb3pDgixVt4tmbV/E45qRjXhG5bzTYbyHf
bWgURFUlXZrIwuyCgGtBPVRAMBNGTKRMUZjX4QeYrNdDEVVpTAvdEWjN1tWxidIOrJw2imAq7fh5
FlOy0qvxgrSkOrhKyNoEkLYbAdUCD/rveMCsVI51gfDC9/nXIZQVlq5ZRm4oGK8vvejFLg00D6Dy
QeGudbZiMbgoA4Bh7FAYOTOJqChATn7C1aBRqsyRljwIGnNF68PfaiqfgpbZ1axVgAY1wGTSmnEX
lnLlrWdpN3xGZ1xRa4Z12a9d4GulxHeogGXLU2aQ3srSFIxSbEfe0iiu9D6H76NxfiOmiyH9cOMK
+GAWht7HJDKyRC+1zuDiodFZTBdsxT9wY4N+NbR6miltWxEFowF57vwLeKgWG9BT0L6GH+4ruyvk
Gu7L8+lrz06FyfkHa9WpTd3LwSgYCudAbjjl5JYDp5fHnwxzGT+p2LRAxYE2TOD0a4dRmvi6/Uw0
c2fXh3KaEnlQuxdrhgZLkltrNoZKTckfDTUvwZyP9+MDpoCJrO2/OS1SIZh3CwiKaDK4Ik1W6A3u
G7szLjyxpWOVCFlbDkKpaEoYtqaKnQHvWKvaaSLaL6RRljqhTDATV2BV2wYSm2Dgvc8dLcx0+xrz
yaaRpyXwTkghrQoBdRwcZYcrvGbSvfU4YcpqRnJnt5PYjLHkkIc82Dc/VYgfrxIev+cd9HWjeFUE
DR6XvQASS+2Vyuy9o/5ytSNUBSVMcm+WfYSCvpSriOwpb2U564pzZPJB7HBjgsIVWnbvEDUbTU9K
HRxi/YNzYyGPzUtFMaaNMx9CvRfZj+tigg5vUALMvcRMLZi6Yi0a0jClB7lTVM3gq2R5QjD9TuSQ
xAx2AR3ILCdOgqauytgecWZr/qtpC76xlH4JnPABVpdBs72w4fE5SpvxerdJW5SWl94tSjZzWUCz
IInZVtp+87qDg1FSm0JeefY7uW+BEoWPhkYswE8Kji6VuR9i8Ou3occ/GOsD6tYCW0IQFXKWL+To
1xfiX/AVTGtvaa0vs4nnd59Z4S1GGdwn9FKBJnvv9Y51U+uVe+yeK9HzCyFwOA66NcqHOGi7QUpY
887GdolhYxiQo3HSKv9ayZkrS59cjBfmD/zBOTJ+7vx1Wsyewd7+9on0Bja+o+mTncXGyXlGrVcw
A8CvVMPc3IveQH2AnkLvrxE/7N2t2uv+zPc0YjZWM8HdtuPNSyN0J7rQX/KzkiiB4qvgzbyEcGU7
pkcIuiof1uAOBO8KEhbC5WV78kb4Pl23+1Q9buBdvfms74g/gcW450J6mpjorELDy2AkTxzRNCcN
2jIUuoDOtO5QJU6ari73J/eGj5M2UKA5etReNikvb+tlkeRj+U/785+JHBxyE9TSdPFB9922jo6G
/IVHCBO+Nx47+TtaWW4LfgTXIszJMsLm1v+RtZ+bdLA89VgZulMVKNCl9g0Ebd9+JKm4fH2+uWip
I0lM2va+TGsPeY35U+7BR2iLobMSWEu80/IqOuV6j2lBMlsuBHBqSCAwxHZ5wnA5fD3z0CieC2QL
1BSZV2eLujdWpfr7VOgENClGB5XiM+/3AoBNChZ3UBxZDINF2r7iwLZwS+h+AB6hcW3SD5BD8IKE
k6NiJnd/TBNUnL7oO8J/EukTBUFRkSzWr/V5XL8bV0jeQYxaMTokySQAWWZf4Rofkx4/biJPRpRh
RM1JobcYM5gz+/OfW+nrlL5TZXodnQma6seW9kiVLJU3Ryi7kozgun+9eBmLELHhsomVngAO0xu5
2x7HoMg8QxxFAtDetNya/uybRWNevX0/l3GU24p07NRbG6OK9PX6I6G0iEx+u38wPmWiUk6bzVbo
igrMlqwzjToSo/uatO4wBntGbWkcEb2LLRqvGCOI2u7N45Xvu/dlEh04rdxseRGz+AUqY+4hw/zw
ZIBQgMyF//S/JIjgDVjvvOWkgmHJrRMT8fb6kdvFm7t6RkKB9E4r0kNUIn0bER+ATraqdMUgy8eL
znU7fqLxduLMMoawyLnVHS9M7P/oEVYlxYsT3dWfETqHOMC1t91qgMCTcqpvcsGpbeS86nO2CZLA
u9FWMJyOT4lAA1uqLzZo2AzWvy3RtNHmgkTD7kurz/sHd2/bLq3H0nAscJx7+2ImswmYvL43TQB3
adozZLXyzvFPVoHw1nvpLaozMO1+v4fe3ZFVMgpjSYWAuj/H0nM0Sy5uDjJdmY63X9eP1WCSot0J
Jr1uRc9SN0lSRJB2adsi5Tifg5avGaQsqJl8aWB5vjWJCgdQ+e9Zw+IzU7NUlP0fTczBAXd4h2MB
vgPIZ5yoU8Teb7DlvGDfV94Unw8xjSnqe4FbU841hDLeXoFVwabyOYsWebPvpn1mMnV/8axPhnHV
uGRLwtRzbcIEAHI27vuMn4TJb+HZVhDruxIg7XsHI7pvu1GwPLMP7kVHHCKy7O1unZVT9eqJmXph
F+C4WC9PQyiVplO9N1Z0UT8f+v7cuAfs6pc3pjXjjNhWIKL/Ov9CZmlPGV/MpuUHD4GbXNvvoXV1
EkUps0c6HJrPPv0pOHveb9kxRWx7VgucUyq2HNTr8jyfHB4CpykJL2TiPShfWDg1SsQGNW3R4ZBD
uVjQZ3BhHVfRbdgdRpuQ4X1tRI+NCK/qBUvksEjF2vNyRH0jcZB0fDohesu7JKWvwXsWNE/JuGwe
FVgA4QTdew9BZOZqLy0lgUbnWBw+GKECmZlGCG/sGah5a+dSJ+U33GNPFQ1xLet6HbrMJp+WCAGk
WILTlTl8biYw4H/tS75/wEMJ9OHqJTfEvZbd3UAoCiV/iu9QMRIAqFRbAKD5MpnDzR+C+/l5UJKB
TZEl/o5TeUgZNM8UCvep48zqn8mK5bPb4xURQcTt1PBtYHIsUag7Uk7Ls6/hTo0q3rQ2T76MPmf1
oUfAwPlp3FOk/jRH2xEoiqIKaNBeSmAq1s3A/HD1cUrRfKpyr/Lhtek9noHC9vO0M0DS3Ki5J7Hj
fdQXVsadNM+yh4A29heDrAXixfovBRokAHkwzOw+yvtdh2vripT2CHd6uFKGKnvrb9NQikW4wWKo
/SceQvGbQpET0Tg9gXfIoXzDxShE2pmdYsSOf7DeRmjndt+96o+vHO+zS5qiovdvh82q+SA3521j
sDzzFR/e7insTOhYceSCLe/q/h96OrP8PTG/OaZglSFZTiMoVcSwYKMC5dH1odfYmz8APs4v1PEp
bgc5dLqPh1ELfepM8myrvyYrKiPBalIm2u8WTzCxZ72t+Um1kD5weZ4x0D6KzBKiNW29ZKS8nNoL
4kNYwQ5nNss3GgNk/Gw6z6yq22wgqB/tawxFg2Ml7D142TuGqDgwAOTItK8LN4MVsSx5IRFDtFSB
3lM/EoxpFNBqBoKrfETiDPtWYiYEFuOn/u50JbJQjxgINet1IdYTrIPVeY2aeWanfy1OpKoW442J
tCGoYpmV5+faeGayY0cAWr+tWKivKVAnVFR25YrIJ8xmfuKeQBj3lOpeO8ceUWkU9356+umxnSQh
ggaFoiLtrCzvvwouqPgDLg+H42FKraZPEp4M6u04vKIE7+h8LWVEBSsq59cqz/i2xGdWUGDB3Tnk
j1MtrNmu/JHq4CTTlIXvQn6PoB+9b8WqU5Sw8iwfMsAKO8/BovmhxIdrA5ooI7PzZebumBk3QkGy
lgGHnNHa+gSIKvsclvlMYTEQL9LLb4y6xkOUlWDs4+2carWK1AesnHCp0Y9njJPpBN5yd6UVGbBo
lsWl1QEf8yOXrbrjg7pS66DzHVj1atCVDpLk6XrojCvxKl2lt9rDepB/342kGyr1u8WK/bSRB6l9
zVX7iI170DfPEqpLHPEAtpubEhnISnZ4M8LRxVTu8KifnnrJgQypv1EgBcvB+3mepWSHWZXO/g/A
tNFf0+OEs0UQ+HOPsdwvm9XTgCBmUbq7wwRoGZmtRDG98xWhPkmcNnwHEfLH+k9TEWbh1rfzN9Lu
0hLlijCd1SmyNJuJ1HL/af+2K+1DyDixOKoM5eiz5LI5P1AGeT+31j7OExY2dHPaCMEoLHBTJoal
dOtvKDz0r0S2CATlpyxcLXFeRdliW5dbHGVGs0+mvdtdnA2WXtKHDgrUXjpTvT51lmSc3jHOxrJh
qBTFgsJ/5GY6+4Zb0WDMzoBm62MWIUEJufCe8Qa1m8m26zXwuxENTWhHKzAbSm+FSOw8pZBLJNwk
Xl9YzDXgaX0JZzwd3AGelpJfWnKbhQoNTXSUh/mb/YFRRBDjoI0iOmaJaU7QVSJeuis6Op4/sNR/
folkToCqqYWjR1V2U7/eeI9+3NlIodPAF0/gBMYAWAb/nyhmz2x/6pmzJr5Ltv1fOuu3CyaVu9qv
hT3kaNw0VIbH2skyijfTzRAJ3DQCLaJ0v61C5k+8+/WgGreGfbfDbTZO8ffhbt5soSg3UXRwaSZN
OjZMw4O0NWPfllqb5nHuJlKM23qygPN1Qtkj6BK1YmUx4HYs+kRaqt+iYJ/A6QB6/bZcA8MouOD8
auGdhR4CsHyEhUBnAalJChA/D4LWH+zPkVuuNwqpB+0kLmgBZ7QbxS9VxxpDgrmAmf7IFUZAhj/D
gcVrsI/WniUEhU2YYmbp4ffaNhflsspuyzR1WVy/BbJqKb44X7AhcRLrz8HgekvAD9Ilh2niBlTv
7YFHYwyZ+X83lqA5Hwy1VvyqK6M3/f1yGwi9rRvGcdA1GlGNNWYItgde8FNFiGNbX1jWGIVdaXWs
bD3guTs7JYemOX9kNl2oGTZy9U2P5KLzKbNV1lCvjUsuvQGkTvO7I9MzbxmhYd9cjPZ0nmogN+PE
RRV3n2zGnM3NrJM/xogQJctWY0kjD7G+u7cB0CaPK6qKZKz6jmrInIP+b1oSNqEWFG6mr9YTOxsz
7fZ4u7zgFV4OqyQQXTKq3XVWl2x/DJaQs5Y69Ma2003qrWFOkvZpw/8XGnCMvuPi/KxLNoHebo0W
lvifjDfrp5DcVVVJY8g8IwUxahVUfWiWVVB8YRrLtD3K/nG0No34q55o96XmQWMCfB0vLpA8Xyjy
gYQxWQSjZavSyW9ZqDXUZWNZiQDT1FFXpYRTKFpdK7KG0cU86yN3P2D0tCxPV8cPYUTTMqmdRm+/
jomzC8rTE8/RLeUNZ3o/OCy2K2RBIrnoDzxvLs8Fit0w+9NL0e/AUKh9MRQ2Q/hAB9IAbuRsmmol
lZvephfzmz6Nak/HXUJFe13UHKFus+NFPoNMmFv3sjOlcCl+5rKbd8Kx8qmGveBW80BWnILkyZDm
Q+GxBHNnEjXLJfMz8lblAmtz/d5Kuodf9H10n3JzLDPAop5EaqGS5O3tm5/FRILs0GpjxB9+mDLu
f7Ua6JaYW2bhci8ysXrpGvZPtTEcUQAagBR9ZvYtxDMySKZhZlvJjfbecer7+P02zSow8tnfiB6H
FirF6MyMOUZumd8DG9qgbPnhHMOYF/BybeD3HlZ0/sLGNPwrTESP5x+GH2kgy7Ket4mPpAfMk2wL
xxb8YGC/38Q320fgauNVhNmSqWnK5+k7uZ+NYwpyEHyeWOLnQGuTt1jHhuXK0gTYJOaZxQ6NdMZK
jQ1P0NoJsYgsco3Q4CcGcgTlHQ58tRi0bdyLaQxeu2kEMxmpXeNFOfJQWA3onQBSDcBabMvflIzl
cnJlsi7qOp6gsBXqZJZlQtw/R3eufT5bd9K8ZAm6RgrKbPw3aop2W/JQMhCR9vGKsUQz5zVcGF7W
KQ2WwcFpLrNuomfv5eqlhFunJGkA6hJjUpY8Er5/EmRyYp+DLTq8jWaDDc3k2w0GDMoxQf7mmvsB
s7FALIhqyLdXNKAGWMdfxt0dExgFZyLB8DWyKXMN6eHExT8VyPssh3A+BKRFWfT9D1Nv27kWakEH
2E1oDcHUB4S/5XSb/E5B7T9traIiiyoHst5m7KtL1N41X7i1al5BRd5RA2I3s5EAI6t1orUR/ccq
LTWk0SsoWzStQn90sORRHLceCRa6DAy0twxFbpuvtpg9DanfFYF0eT1UYLkj2yFJAPVQIxLBoYc8
/zun7gSq3wkEj3rugYGSfo4tHyz32CeDGZj/45VwY5AOqD2WD4qgPutPa5BuA2Mtiz27c0doHzo3
tRkNbirNpixzCdrd5V7IUWupNyatqcbopSN3EuG/P5aHCATDfjx1zb0sXK+0uCTIFQoeEyWQEcWG
u81dmn+H2qMLSWhDyijQo4EUhRyAgC5XCpzH/Dee1yWoa6nuM7iW5ttMn5nldDUHyhQNtWvgnJ3V
uXze8CXSL22TqBwZxKltEgWNvGBmW/dnz7cAiQC5wznOiVO9TAYJfii4LbWhADQdjoQR6sdAJdMv
eKOCN0tkAi2QaQ+Y+TXUf6I1f4rJQLAfY2vIg3+4NES/+GW3gqqtImF43T5SgsCtPvZYyI+YYSP5
X8NUWXOtMXAz27xTC63MxI+mWx7UtqB0VSZrPb4grS2XUx/0LlrbpP8/RofA6rnxX7EgcAUHjXkj
13G6xZcWmxPEVX/O6/ZXdI2KaF4gt0uBAXrJTfpdILh8dRjH5L0UpeeL2BvmOQpfvMXg8hP9tExS
XsK05Zgfou+sXEF3fgJAn2kzen8pyZgbBxfF4utHXD+Ux3ngvzd7ZYzFBVdC7md3u1orcq8YhTSw
GAwl2Y3M/aSjsPvGTHuZUdf2F/88kcgnkpym1HtLZhrTqw1oY9rFNq9TNqef2xeikPFHENzFq/FK
r7oitALI+P2OksxJMYQ9AKrc7cYvYU82NasrNgmL1rpY4sgl1+/cGDFfZmqr54b3v+EM0xvFN5FD
DeG64DqeUDh56QqvSBHldbtkXSRJjF8H7AjQHuNR70H/l0DwV/q61fI27F+y+lNPQCJJIG+hhEdY
IwJ1mTvhLyiJGvqRIjXFQwYdxgMAYv4oH5yOIhYODWmqyr8Y2DJatGExdL9KLMk5VTdgeJ3AD29H
Gkqdcp0b+yMQS33OFyEEor56oXWikl7g8QW3xGrOTkSg/hIn4l5oxI+vf1O1u6ysD0fapnqJWfW3
PWPQ+JMo5S+bLPwEUHBMF6P7kP2cBzudg48CyhsRfTitxwegRxRy1Yc1sM4USdgHjteIgDJ10uha
PhS9n5YTNuSwvxxO9NHQsXlIRQMjFo5nLWrvqTr48R2vzqcH2FB7ht+NHOqiIBQTaiNqCtAVpCom
sVWoWqTPZV4yQRiPoUYDpoq4afcT+AAgku+h9p+tlSYwZldsONGuOrfp3Ez3e3bwAG1bZgUmF0+d
lK5wh+A0VV6NkOjT93PUVhDPA+jK2OkITTcx4EMFV2JaIMRD5mjtSTJUIbkA9QQ/PPXCe1DiLr+h
6MTCNtbKFVh+rOOodfGlwn9KN584P89K3esOvMFErlr9txvDwmrsvyQxEDdBjWKoVApE33P+3sgt
8476O1NEtSe7MIlkWH1CYxW3+QlvdW3M1CgMORNvK+DkuZxT+6zGjRTL/eNsUB2mSUHjLTWUHMhl
lEKWzK5345xVcSOJIk0b2cerngyQMYCpFtRs+H4sCKPh4FRlM9MsvlI3YgGdUCE7ZYYVY7aveJ3A
dko38yAqI1JqG/bbtnqKavV4N3Io+gPd49xb5TEpFWr2A0NwCCBFyIfwWC9LSGUWzr9AL7KLAPuT
/edqalle++D7kLshbccDC0XzVLmlCISyOBMa43zj+EDq4DR1WztNJE5k3n8WmFfQsgojZmt3s+Kt
WbmE4Q0vDenBLDR5cNnLM3wr6B5fKQKSYMBfhWUASmWSmdTJVcXZ31y/bN2wfZapiNX66NhWGPGD
smR1ZB5UnnQmAxhXJpW5/QkjZJXx2NMdzRf5hVbR/qrPZsgsOTgf+tE87lNqdeqFzHH+essr3Hx9
sx5gDELzzp1c6WnNSzS2Tc3OkwnfTDH5QGh7CWpB72b2ssW9F2+80E0bN9ZvZNjsFbmmLYBW5Jij
VFflOiAqBLmTk7D3qQ/rR7UXn9WZYcnJncYgpapCEcjA2bzrWQjxXlfJMJAhj15H0X66wge5D0qy
OyRBtCE1nPko82unTZaPCnDnSQhmrR7XbEgkwHyoTetS/Kq+bc5097heEvVD0dWVfOp0yLXe+pgD
LuiAfIwdViWdwFbS+2+IKaF5m03Jdjv/qih10W1+kqv8k02VIq0sZmqvQx9kyFoBw1GDopA1rzbz
pB1BM7ZNitRZ6JALvyRWvYmlvnq69/tebITKej/JrCQt9oSdNjmRe18kTNk4MlULQtYbcP8PEqm1
iChhubJY3sB1rb6+LlStp5yqlRbX9sYn6wMZBw96GVNkYM90ivcZ7jKukhmtAE7rHE8zpj9eieHj
JQGFyVaM7cKFXFz7BtAFjb3cT0HB8IZ4SFiVmqCCLTAEUcmonsorhnWRK3eqYHJ4BQiFvXleIK7t
a8W6tLS4fShUXhpriMCWhPr8Rdv3MaXSfHc+7hVvU/NPFX/l5qG8wwUNgw+CGba+s/A4ArlJjOs/
+nUH3H/z8h5yAWNdObaLXcdOiCtgXpbexB4v13ScdCcV8hOujHaEeN0hikydXkK+IMvWGNFSZ1S/
Tdfpro09cNjBCTWB11x4oUmJZ9p92vhDXEeQloo7YKf8jpo5/LzEIbMPZ36vJqK+wzh2f0ICUlvc
r5L2vG53sb+t6/EE6GzYfBtNLwTRCvmHUlGYGRKwwoQvungSUj6H2FrK7RAwpKRnc/eSP1t8gB6Z
vtLWh3Vl0t8rEcpNEMrh4KacIv2Wz+8QNHj9Cor5mrYjKXwxHSr11VAV0j6m4IXa5pM4Am+gORdP
wbKiZn7MvM9WvTNeLToqyETDZtniYv+z3srCYw9Y6KjVqbnhUnIfl16YtgVF26MNjZw7813RwmVe
fMV+HjWIDhT2KA692sePQHZYstRphmY/j7f2kgDAXUaFhi1vLziQgb1i1+kkBK3VuvFsL7S/j/jx
1pHyMNIOZLaADpAzJrrjROcDyUYevfDyYvw3ABOMI95XkczCdA3C7D/509Livyt2X2klEzNSve+N
KPNYDG2su+inX/lYKq53umwRr8ylT5V00R0dbYGBEGTQ2VtCU5xy3FIdHGXAV5O0W8J+IrnkvaoJ
gZ5tsL+IQ2mpUxX3djgUWImxESQzzY9ujx/pSN9rEmEgPOc2vTjs6nEdOno19W6spBCjujNG92K0
1ULOq9ZmqB+q9mPTuhK/wqODtCRp+BqPRh4HatFtbzVR87pzNUQ7YNjqwUqHO7+OvyiGZPTZSTRN
1Qmy2SYIStMuIMz7gzwpNG4m4dOxkXqhlUmHlPWTSy36c4vlXdjQQBPGAzJHDVKn5IPkJWIxXkW3
UoLY0clximStPwVE/zS+fZ3ny+7a/E+7B6hHZjadnYem1e9FuPSdROkO9MqomeUA1i/krJvhvPbt
UnP/rGXIvsEpK//+hiCxciw1dCJIat7jdjn+zmiBpE1tUXVbBYbpxSAfhrkMuVtj09OwcVkKBzGO
oNO0Vv7zQgTTolKoupqmpaU4miaJLAEBsP4O/qcNp4JVG9B/s4KByVfh0vZ8aj47hm/tjYRSdzTZ
k7ZC0OMygyIflW4uBLQmCl66NuaCceMvePX9RFKZOCYGBaXiJihkKRk+zORgwzSkpxCH9/fussuZ
/vJwH7s1GtA2Cx0LIBRSzIsvF0lZdvbErG1itxjkh1G22HydJdYE8jquagUn9bsJUu5M/qF39KJ4
92qZNwqbDqHwLwhYB7kncyh98a2bJ27u8ecYP0egX+e3DUJ+yTqe5OArVRN4SrZFe5M+GhXPenY9
rRN+RfSzkW0zkkFXt79FLbmvpWOMcdLq+agI6Daw3VStSdq9ChLkdL7z+IEL/aT+InL4N0Bx2/jO
QH4JbYASNRrS8aG993Dt+Rp62JZOMhO6HIO+yA+UHro0YO9HAUG5QQrm8QlfJhqwKCGwqNPqjVRv
n/ucBm8XeFMn0s8dhi0E8P7UqZrDT4oxbTQJ+L/e2nNdko6+IauSzqmYs1FA4y03CQuRELKXtoIu
iROk7Lj4pTQ8lkoj2xi1S2329I/8jC676mPO39B0ZxiWNsv/fiQvAAcmC0Pr0NvgwtivqbFyo3y0
nZ2Xpzn7ELHR8nvoNPVjxWAdzYF/MFdtA+Ly6NVmYElWYKXm63puwYys7hjAl0zjMrvtauEhHFHI
gJqbWEGbgYRbc25CWAPcLM40gxznMtFKg9oZpvAARSIsg69yCQsrz0QXVVliewx2HZYxJu4fVn0N
1N8BRbWe9h6o6INAUeeXZ0rIr2X/iWBAHrMP2x5CqfAkG1nRnO/AZsl8ogLLP5V5tieYuJk/Zahf
6Hy02cq/ls/fSWP3MoRyuHYpXzuIzuBqWMVtYbTb2E8bINBdRfY0NwxqImv4sBrtENV57KjCttK2
SxEahmvG7OpJhPWhIHNQvVczBH9n3L0uWGwWrMb/P4QuCX40Qw2hVIixWyTbEDwmJnZqiXCICnI0
1C+XcJ7wIE5K+Py3CVrmloKRp5O7TDIczH44nm1bYZaPUMAHt/PpIIUkw1fNJh4X2ShGJ+f9uMbR
D6Uo4v/ObZ+xwL1uPT7ldey+hIRv0zjwb4oyKTKrQBhh08FBqJyhLFrgadxlGMpkxPjYVjRI+ZKN
Aw7F+yBR/VBLGEMluEdSAt6fGOT0JHtItTQ1jZm+Q6DzMfj3k9jbZ88X9oIOx+rmt7YZuInuKzb0
mXU8FAskVGjlSMh77MfHEWvvFBZB88dCWnfOLmNPWo3oyG+GAVsSsl7WG9LCKX3LQLQK+TtoFZMw
WNR57kTSnSt4akbcfs6sPOCmnGvsfzp5/CFGONbiIaeBDh2mXqZI7vNlsfzkJ+spTT2kJt7hu2gj
KYaiFWfarSCxCxADbKVhVjvzQBxLAlOqxnNJkVbewHXQ6QCfaHpGrqbC1zRZosAiZDIlnARDDgHY
wvoGKqJokkVmZ/ZD5hGPU+VyKRLUWQDhCmi5NXbfPxVCWr6thri6zv+GyCkerAFiEZjNYtKNuJq/
BABFQ2V5Lk99pMOGtpR8w4ey+q6wxs2EkH/1eJ9njKMErURMROJflOaM8cDu+Ua6F5N8WL30BVHh
wfz6qM6vl6MoRn60JMwgfqxKq+xqfjgOZlSOkhR+ejqm9i6QqVpTl1kmEsRt3W2aOHSpP3K1Ugwv
aEnNanMT/RWXR+lANnqKNzJNme6h3SBASHT5E0ZIzIf/sWq/2G+Ddk5Gr+2zAPifluPn0JmaJbPQ
56sPMlPpGYsSRDP4VuOmRsBxTtC+JlwPzFIfd6Wy3SSmdVUQjQOk486BL7tMg5uD0a08RE3M41nG
WH2R6dCXHcEICO+zx3oWjrTrYW3I7uYpUrs0NAcEJlV/hOVQsY1yt2k4yV9MQLadzmnytYeRKBBs
E27BNZAGTGIdxyG9ZYOoRW9h9dhY3l/jV9MX7m2SoQKBw9vwTvUxrI57xceJGotlt7+fcE6giAqQ
FhTBYyml8dZHLoMu/7ioOfgpql+7ELdotissQVYAIPZLObLL3mrFcv+i4OJ+PwtmGWJDz6h6NEOo
AEeKJ91U7F5LT3XR3Lub9wH8oYujmLrcjfw1LlYRnRC6pWe/CF3crY1eKWeaZg8IV6cJpdJB1aDl
Ps1U3Gfpg+yo17Q/VuRpdeP9BefQbQAvxIwmyq0i40UKAmEslC/WHo1b071zjh6h5JmnxkY+rLXg
RUYGaQHiJ3TKlRmpvcz4qfCamrYN0YuBXmDLQS6Xqcer7JK3RvBd09RRHx4le0cXC1NrSQiNjsJK
tB1HiEbQ6vf0ZoZJSEBuOokv2l0b00KTvYGVs/2fY9iCEjoinEWBfkjx3PVbGGfMU/44ZAvDSKet
f70HIVIiLTkD3SCvif4bEegjc9JuySR6TOMThvVnN7LReBwUmWmuDB4kT7znvg64oDlGQWqWU+Nq
1B/SlFtFWkUegW8sPuqoY3FLIJAMvEqXmm6bqOVnIIAnxx8D0DiYeSE0ZGaU2TJkwncT6Ell2Dh3
z1ujPK7YDO/q5ybGIsdBBze7juSkGPR/u0u8DyVZoakgMrQ3S4bhqaCXkkyHM4+np4yM6FK7baf7
GZDYqZwqrTrCn6jAcVi+464+5G1hQ7Lss0CJEu0w7cYrA247jHFW1j6UpWQg00a0Wy6rO9eE/q1S
o7snHzrQd4qp9SuM3l4/PKSSPn4NpGz0MpjzvH/At5X6pzUzeYcxgSLUMyvzCp24wC+l2el4h/94
7gKIM0lbWP9nI2QlKpUf18jfhLmJaP4kc245h5QfQjiYF5WVSSgMltRyGEyCjOPV9OdVBDm5EBZe
tV9ZwJ9ZykiQMAI7dgU+/sNqVwqt9PG+G/sqkRyTQjtum5fymFwIeq0OTVkI8q5/jNy6iVgiqVu3
cXXO3Qo1Tm0pvduFSeFzI9+To2NLgq418EPAlSzPjDaM+uH8L31iflZZCzN1tvx/VxXrLNt726bJ
kt8kfjnknPvbQ5f8QqBQ2P0da3C2/yEFqFO01J96SLqdZScbxB1NaAEiWaH9WwPRS1RkX7ttMFE5
sgrbN/27gzRj8JtvV/iWvvR4g3ysxPB7w7AKnjPPXN5rcZw+FlA1VPFQxxy2mMDabNh6Jh8QVkeO
BREtsrYgrA8B5t04gxbD4AY6rr+agiNxef3QB4ZLqLLxFDe8R27OZ5kJMCHE3lqdvgSWLQewwriI
nyYQ9Q6oNtrIlcbuwiFEgCwqPNRiIRVgLm6MyGFmNCRgk93weMcc+U1Ugj6QAt8zwUgkG9DykM0A
ATdrTJytpuEJWldaOkkqIZslnSnW+3p9sQTPym5puTErV9O99lLzbJ/Sro7fLsdG5hVtgVd44B8z
ihTatWl3bwYsn/Q4+ga9QJpcpyOkmNPi1toSR2Q6ttK3PfueFFCPKF5u8zOB4uESIcObm3Wo2ZnJ
B5DG/IW7AFlJ2AFX+e1/Q4vv10NHCqDT9mwt+Dtx9qUgcz+71fA7AtYVdNN/aiaGCXlCOp62CwEV
yQ3VMRz+yi5z3JMinE6AgSfh2zrQbjtO+MwO+MW/tMV2xqfZeD/zcShRJl2jRZpGF+ZLJjl0vE9b
zNaxXwslzxhNecMtWawBZrkipeVHa0lySgR3p3esSSzwievJLLjFRq2pVn02qrJbEVDxYhPB9R+n
ZJzU5yMdzmtKd8vjM15MxYkymZd/BuHg79fVYf3zVduHv8HM8toMCXPu6W1qFqAbMFMJsXQkpkdW
28QOYfEztnQ+VyNoWJZCDPU3xVwjxfR0qkJKiEQY+0DUvBxr2OnW+3HEgVWX3bTZcyjkqlwrGQr3
Gvkq0Ro8m79Sy8X1QvABx32A2muQR4MX+euxl9wxzj/3VkIDAxYf6jZVbMq0qI2ye3mDVF0R3LLt
as83D86qbSRFvaM/j0nL/eoosPLLDuLt5pcCtdKoZ0fVhZocBh9bSoIGe1PSbNNRVqI0nSl34h9y
0MpPxgKaIS2uPuhAQ/GdSBL5gWOttv2V5ZzsjlV8Jyvf1YGTgk5M5vPEn1qEKic4W9LQPyyWOwq/
YYJblQ0gcK/GAdnMnaDVENzhzPNa8cckiX5Rg+lAiXKBiMbsOpDjBQy9rlciG/ZlB3nDfaKMKOME
s3055/lquWtrRfVFnrvZe7nP6mQfDxjYo1eDfUkrdnKE8xjjj6C+vGHonI8vtfAC/yzGaeu5ZHUs
KPISosCghvVpa5Pxijml9LJLRctp+P1D87G9MYgbjDwTayDC+u7SFkFcVEh5Vjhgp+dpF6wM8MOh
Z/wxe121XQPwO+wOOGXgU1CW8z9/g6JHXyML+3ZD5D4vOnyCtE5EsyT1ZMVTwA+A0MVNYlvsGuk0
7h3d34YZJM1zSA87yla1vmsgnDRWNMBxZ1LcT2+h7XgtGm/wx5/AClg80NltGlqJQFUalQwNFmDD
FlKI92uHK+hZRVx3JDyWn5oz3P8HiJwfTArhim142ciC3910QQSajDpGs1gJkaIJ7vLCh/g3n+Wi
gEbpcWCR8atTvXyZ9Io1h68j0StKGNgpTbdLMVh2k2xfcVGQdEzZN/PEVEUIR2m/sEIb3Yd5M61b
V+8PqkzFONE9sJiEEJF5i9lJ/eOa0Yt4oE8KFgxrEKAQB2SUIkVQ0pC3W2tB3rc5Zcw5+KNRXQNs
5gjoHyAEqFiOyWQt1Vl5wu4CGS8hrGSZBrjVTDCdR+mqj6tcnkO7Mil7NBMpGKS8OZPVZvTU6nX5
3iQz3YBcY+UYj3lClY10Z63rwo3ot7PXel1nkcbPa+mc/K+teXhmUpLAx5zzliq8dOc9VHSNBROi
ToL+CKghuYWWxHaodeY/yUClRy589cmO9BqzmbsNOJ3ksF93/8Ta6SHnLalcjP2EMH0Wsv9+yuyR
TGa8lBlaf2WlMDamAkba0JJaBLM9rc9FhAg9IwLbgb5Cow944tJkAPyJ2FL/FAnOrdvO+2+E31uP
xVZSXueYDAVPmw1n8319xDVIm5w9edGfJJxgu5G+DhvvMp7d/Na4KbmfT/IGO11nx4svsJS59n+V
f2SjJCAco9wzwGvyWfBbjwWw5Kt6CtAcGmNON67Dwa5k368/EhzkM28dY++iJt+1cK9i/Q0ISkEh
BO/yNbF6F7cIIgzHOITqVT8ff8VGsRjXc42Lti0oiyzdbH2KPwSqYDxUzsJxLhjwAP2PZcOL7KHn
MPBcLKr++YaHbX4fF/DF9p8zX8/XJzczqtkOUJbaQIySz6+lWSQYGSzrU+3FPH4yJyoZNJvBz/yO
nHCKR+dDbAHHYqLs1RB7qwpMRL7+IiP9oTThUB1X+ArOg5eZI8znbCSF1ZR/GkdlPWRJF84kmI/6
LqSOcKdq3Q/Knn1WGPoRnl3KI1eoNQvGV63WAeAzvMymBWf3n7S0BKA/lq2MlaWpouNqAja5PKWp
lqym6PL87uWsIUWQihokxFlUJAjYm4+89+AoXBbcb5sE3EgR827vfPs9s47mPexzwwXCJgiblKH/
6IVaLaYP1MXSoAqo8v3b27K+NOUzI5dCOzjUC0MBDYVX3TqllRwU7Ma+eypvbPet7GGLpQTfYsV3
4J3dcubDB9zWxVtCzRrjl85vLMKxzy5JTXkwcgn/0C194WkAXAeTxg6ZEcTyXLpn/W3FklmWrWei
obSfh+65IuTSxrOOQ4y7U2NhkR6A1fUJ0ih3EU5rtLE5BBoiDPJY457CIiCL8eiZSfpu5mA3rL2p
tDXycVg6huof/YIDpmdy55FAD9pr8xxWvTjZnWGAD26q5c02jdElWwYb7yDxaToIjpUv3xBKufl6
CPIfaLr0x2ufo7juJVmP6DLWpclN18A1ysg1nbdMRRdS+n5pXSyELy0Khesotc+iBiRp+NGq8Izo
5MgREiPYZsdkpBCICBYMWba5V8Dc5n81ixXM3kKMiws4OnllKrz3yHjGDSaIVmS3O5C2gTEN1rGM
Q4Txm7gKiWYO0Z5zRKKl3UAVatFL/4BKicuUBYU9lDvfCrG+ORXXSG1wEe3ca+ZxAA16evg1lDEa
a0RnMOIve0z33ByLTzzv85d/WT2/NI8GUSVQrNOF3itmb9PmBkxl+ribWO4bdXQkOjYs0lCYyE/F
i6FC9KGqsZ+Kh1wKgVYZlCjVNj0L0icg3FjMgajMAfVyMoPfIbif2QCXpicQ/FnEeNVxmJottlwj
VUOzSrUlenuk3gl3sIBPv88MREI8lQ8O56l9b8iP32A+IJWBduq36Hr4njgiScNWMlVQAGYwsSk9
i+tVqeYyQ0/mJUEyLc/D3M4ZIRNsCmpQQzuKEkxS2RZN81x1TMSx779cmgK+077Otu7gueVZ1X0F
cj3gaNgumikntzn2eF8OiPH2zY1zlO4ie2ZDCLq9efPFzXrJfAt81TCOd0Ka02vo8ELM3MyEWn+l
fVzGxCSiqt9ZrSS0cTJFWBNBiHCUsSPZkOHQr+Mri2uxGOe5QiFUJMvzqfqO6pmssDgkWaPE3dt1
+3fnb6YHEM/hCYHthlRG5WLt8q1RKa+NgOF1q4C7I32PQ4CKMs+ES0rl2D+4ady4UjMI/i18FQtR
qglSLqL+ii8BBIyS3esinRPJ9q29uorrZVGQBjWKA1KWSrpJkGRhCVEfWPSSJsvJbNT1oxkAsX62
/bt8mHcf/LuYcu6BfsMxnOhrHpEXr0RL4dypwqfV1gBxNGDKZEDew5SnihorVO8lWfJY/8P2iIe6
FCurXNrgD7jqPvpK0ptS1/emEgdCC/3+5M2GjkTnqDyQ52K/L5uv+u2whqka3IiN9scIuFgJBlEs
k6iMERrKKq1K2Ne0zGi6LL8iHzktoE/k5fmIHB/I3yONCR8MuTkoW/yzXf7bmBd7HrFCxwjcRJEO
Y5rSX9lQwm7Ysz0j4LVpBE056hMyEGCTw9DJDctwNpyxDtT6jqQoTHuLW6xFjEqrBJCBM9SfesAS
IOYjhumu8fQsLBspABik0g60Pu1jKx9pdbwImkzswKC0gJhAvH2In0lelRABUex2QQo+xFmRYbyM
+W+keP/aXx0aL5Fi5y6f2u2CderSYQkrYS0QDVbP1F4+T3oidB5YKhF99/b8ei0odux4WZGJ6dqE
/AZVHMmx33+XvQ2OxBXnjDWSvSWB9k0fN+QUrBbCDWBnmK0AXbQ5t/S6A+AvKMdRgDC56yPwcFst
Acujkmr30u/ScBzeaGGP63ptydf984K+nG65qAkoLCdGITRHq++nT4e5UoRVTw7Y61FAPnP2snwz
XAOgGHotF2QTbxCPeFWO91qbYrOP2hyiXfZu9/4WZvSmX/PlCibQsrf/SPHhCSJ220XQgxgiy8UX
yxVsVCwW7IGOzAV69xgtwxeZCF68TnrSxfP2Eg/82Zq/GxthEvQzjBnCk1i7kyKddX7zYrYH2WTm
WwVfEgPQua9GO2BWNxU/3cZ/bijbe5wdv50tjYWK/lMbMdGlvPy3zAZ0CoBN7Td75MosE97Ytabo
NuILDQTbPbnPyzboZ+siW00nuWSxuE33I6xzWqmHzprkeQZzYMFgxHiR6MayD0HDbFVhLJ1e/ZqM
Xm7ACoWPm42unQYnUBvZ+xh3gMLeTM2S2X+/qjrgjnLaBuKRuXtrLFwBAWZfMZb53zOF9ugqw76K
yAZu3iBEgOWkCLqKQT2XOJQmrRe+NEl2GjtPoJUUpf++kU5DkFJ50pv3T/BxFY5coRZ5US08rPhc
MFnEZogXRPIBflXDKLZYpIvVrk7U2bZQ0f008K+BfnpQHKgkEYUPpLVKuX85KskHSY2H9rOItivq
SMT8mDOh7iinRB7dm3/ZwdCSRc1kjkfO80dJITsYpebsbFE+cQz3i6hU9qJhY9UymHRBZfYs08KH
/1W3C+NvU8LswZQKuSsIjgM0z4FCyCom3NDwjOMjsRkk3MK81MH7VVjA2nwTTMp2N8A4yKt6E0cs
lR6xSy+4FXgL8J3+QocpdUlqi2oNd9QZBqterownJnUtNc/4d8UFz7NpgvekHe62DiLwyOGChT0F
U5NVnY2sBJFLerI+aImN6ixHt9MGE0+3Z3BVUWEqbNmgl/vmZ5X+FZELlFdQ2LGQT5VoQ+csoDet
ZK6WkG214V1HNZ07CVaHi4KsmAAucIUOxsl5YN1sRN94Z47L9p4Sx0u2Re4fXGXNzMDKw61fhvpc
KC0JZAIUdHt/I6mb3UcNT5VtGmKT53uyDajLoI/OfKDIv8sgKEJOYC0FeDeNu7zlxnZmiJzSe+8+
b7WbAbnp20vSPWrfOCNfDwzIkzQylZhNUUuY8t/98LWuC5/vqAutmFITkUGPAJ+iUTHLED0Y3clI
UCSxNb5LV64vspP97JtMe36F+3ebh5SiKFFTY1H7j1ZhzXRX73+XZYyyYZT3Wb+RLwkH7iQGts+1
LuKZRh8P6w62pH9tDs5v86IgyXrtpKpbWtjnmb2usDuR3Z81y+2MuRTXZdnjOjvPU0f92Tv1jxb/
+3CKrW5hv2aMBZIZ9yQHe5rOFXus7uRgvcDI74NySjDqPDZPYz6tehQsYzCA1TWFOs011INJ5C4q
rxzoXcZX1X5cAh8G9PuwP7bdrpkaHV7cMckEpR4qhIMFtddrJwx0ROMzbvMJ92t0/it1aDZgNBWG
GbmxLpMhN38uHGkBtun/YonasWIB0RszGqwn7e+9Ex5ydzIdKVzW7E6vtN4j09yGiqsgCvPYfEdG
MGb0Te6Nrano+0ygnmz7dqgUFv3V3A42xd81cZbokIXSNFIqSW9XOXS+RfXNAZQxfJTFYCc4tJfQ
lfzdNcfF7WGKAMmUr1UTQtW5GbmcMqJjZ+s3Ez2hjvCfDFGybTlOOtTTsxBAh2OumKQ5f17hks/B
GYPMpkZGzdg+cjqZ9HaebetrHHdgfG2rhHRcSryisJ8TQUIhYBMbf5GWu7LNpfPB+A5kU/J8Me6C
8FuA2qjZsl+fwR/vXPiAmsRcnKq8S9QFh8FHERdjhKnLDeW/x5Gp/0VqMsU95XpSWytba3heJwNP
LXi/qVd5YBu9yDhB061rQi6W06csfT2yHyJTXpBvdY9iN13YQ13KBGsXIcmDH1nvyba4LRv/6PYY
MsvEg9FtNN8koilLU2bxQqF/J59Hz8bHnbUp7qkQjTrQfaJaaJQgz0Y0dlaQGO3dThXMoUMIyr+M
FaDcAnn5lcP8g7F+5G2/x6lBzRQ4L1tS1UALjBdRCyzcCFnOc6yXIAOw51SfUbf3YlGk7gpC2oju
5HyE89lndWH487ItABfSM4D/4zKanh2CGWtKuPMKoExnmWU123NGNf6hkFsmuqDLx0VA1FZtcc/t
/ZPe0kpBejl7t06UrY8YaQ6IBtPFhjk5FEceDgpmMBAd0AgFMCxquhOfE57VOXLGe9GwB4mUQJRs
RwYg4IjVT9P8CPBupILsGJuIzHS1vG6rgyUtg1YlTZq5mIcTTK1rmU4Pbt410bu8mzWCP98ojzn2
zOSFX9dLD4mgutXHEQxOL2IaWDaGvZA+UlxbkShXc+T1nLU7K4rGrSyyWbaP2nXxcqwGLzRtkwTL
dMXGRuiIEIvNcoQy6sXfshJeq0ZmiES+NyAjpcVbuCi3ojuHR55DcAieBsNwhL4y0rsnMntPkhfy
4xOOSP+kGHb9v0oq6EfKy8L6mnjVXW+cPcBgm0wZSgTovXGGn0eQb97C93lE2gLgkIF0kyvWMP/v
AYuskZf3KHH0hGo3ZES+HIOc913BLIRH2f9TvXDVIHDmdXTTeR9OWMn/EznfwgPYTg/jZ1xQkBJ4
4Uge8g3quWu60yET22xQKK+IggeafkK02pIlIitUfV8ci6/9C6XWKazX+nEjfe/ubtiHi+2R38p5
u3p81+oFyveJNvV/KH5oCFQKriqoDXLYrlCDgXoYskHFUGjNYjOoSyW3MtV62czA4MnfyFqvAu2z
Oc88NaKXBhqbkkA/PoVvFXMOVUyfQbgyDp0ChFwRdK238/kZDLvc7qapBLd6SExhc2yzy353DkDr
sCt09mZ+Ccw29i27xNA3TdPROzv9XmKsCDni/XH3IBJbXxqdM4aenc+Pp5ZQGwDTzBt5d5wtCe/E
kXxxOrbhOJrFW4AIthsgaP6J8CnCYA7NmlsjJtdRgLnwGc5y9T4dNMQTrRlMTKzxWJkzE3TPsAhL
rIL9G94Up1geJg67RpLp1qG55LRgkOZDnFHoDC9VQpZhWzxN0QHNLjbyQT5gXDvbqxiG3dqHEn49
DjSKnvRQil61lvH8eCKqF46lgaTizv5NosGsF41tguR57myCWiCs6mbGXNIje9LJB9GE1lhGxpxm
NVWWp07Qa/9iDrKEHNq90exqoTViBMKuB3U1Wy81743wbMQQCr2igpnFvndysnV8/BRnJ3REGRyf
bTe3FDbvqm/45djaPtrlCkzM4/hVuYYqE8IvLXXLoRut2pl97ZeWJr4Ru1dd+T0YZkzzn/D6kP3P
VgBEPl0h2pPyFtdBscPL9KN1C0wBjQS9JMDFg4rBei7oyBa6mTHiWyMLwIkHGCRSjoD9wCZNl8RB
0h9Mwz9uPFldv58EMGFWelXVsM20Uo4GoPru8Cy/3eaJoBwCW4exUSc23dmKA4bqPUGWnBfwmiKg
xQNS0WvFnOIqHPslF5mGg+2FMVKyrYelaZ3gnSR2KwRZniN8g0iO3NoKXxLwiR/b/lGX0DOE4geF
HBHiGCrlxlv84SsLW1IqONzfvcDoMfVU5KRa1pQRs330UsSIWDLA4s9OwDW2bgWkUFKH9DAs3vEQ
TDfUgyagclkYut5+3VgCLd4/SB6hbRm6yHDG7CdXGQ3ECKuFlpqiifcQkJq1fNBRKE7SJwgfxgtp
OeL7UT8Elpil4ReUKz3fZCXJaecguLlGZv5ff1hBBzxv+1cu0ALYE5CohZikfAPQxN5GWxFN2Adf
FU3x01pRW9KSxBJIQkPcFFngeBIiNPPZN4GM/y7Uxi5JgqNuCpAt/9jgTpZd/IXsAlgsjJz4ezKE
lPL0KB3ll7eal/Iw5dQ+/U3ThAqhwKrHmpowwpJ37/D1SCz4bwx5FFTXQhMXO3e5zw0nmmNihTGE
op3SrwHzdopNsw0+7EmmxxhhYoAkeTFOqnDozxo/0e1kaZ9tix+Z4I5GW344dTYPB3YPZ34EYnsk
VjfKOAUsJ1nELJO1fkjbU8QTQZkbJRfLrbSlG8tzm5esQE8PKyG++O/y6dzpgeHaVd2aBTg5SF0n
ezU+yjNGT2LZXiMrVf5iGMXbxvw7pDiUnln2Kp0QblpPCxRhza3cqYeQBXvYEgpeF4ODqImSca41
CpYsOVxJ8I1Rplo3uyQ+c0joqsColdVtfvwCaa9wv+tWQuY9nMITPw3sfR79Qi5vCLD5Jk2Ny1C2
AhltjjOYpg2D+N+14D3X+ND7gMeq31NhP9pEaPGjoFL/HIRCLllklpaGov1cfYmE3qF45+tfnYyo
ahDSvP3Fx0G/1EJoL8DUoebFhMQOLT3Nga9XMhD1jAQTPruJYPqLQ9Re9bwrN8sG+T0kEFpZizFL
5Z2l75Obgpq7MApu1X4Dq7ygSa4Dt/j+77yZQRjtJUBNsX6TdemAuOqc5KO6ENWX2t3iRcTvgfD7
iuAIHKEo9arta/hnqnaWBC0IIxk8aQkjRx/KE9iSKHVQNRX27XCP03szAl1X8MHsVBJ/kir8UUGN
qxfICGKR+3ptCQD4gv4OvhYj1EuxTfP4bQJVlZX/uL/RdxUyTsQPq3G/BLlG89tNxZLDUIBLu5Y2
GlsJ4LM0Nyi9POWLY7ZOATJTAOIPFh5glEmnOtPIB74jQFRr05qYo78QxDr1tfDz8xWzwVlsETM6
uKkQ6UIoIqRNX0Qg2iLF9uBT5N+LSZJKsaynnA23xZM20ysKiOw3xFveS80yZkzePesD9Umxyjfo
sK9zKspT1ml1PV0S8YKJpvflmkQE0xB0RIA8FNau1Z56xt9KLUgrreHCUPeKF4I3WhFU1wEqErcp
Y4p3I/5HTKGSzeDlPKL1VlJgdngUva4Oeo8PIVgyy481Q/97zvEmJTqFqhVczPngm68bh/MbitHC
uHfImYK9nGljqu0eD0A5ieE/foI65ug+g5aAz/gVyCP1gV8aMklSewurtVX/q+/DTJGOeteirKvD
KD4f//GMTDqsOPGVgqBNgBFMo4FPSvV1fp5SEZgJ02tShC8qxO5hqzC/OMZlu0QaAjv/53iYuRfA
D6A1p6aE8RWVZXS5p2BEVAGe4/BvJrRTpRvxK+YkUxwUEHzpPJNwMv8owOfXHpnSt0LTrpBQkrj5
rF19b8/0HxNix1I4y+wzB807J4GfL8PRL1047LCIA/bqXC6G2jdhi8LkE8v2y95hlbPdfCj7RzJo
XfQx7IM4K+jtY0G0LBudHCht4k3OW11jguMb51ZrvoRDaZJr4Uh5SqoN5XnjluArhEoFEQAT+nl5
3GVifNQH6qCxRcXS+VM40jmx47xAOU+4vUxDK2nQgs8BlBAoQ69J7EGESSgpaqH/uFvlnU+Vxj9L
V+9ILLNptwZavkZK6IfEsQubfP5bjiYIn3xIu4vliYV6k7jcVQB8ojua4qsiY92pXPAgwsYiha4S
unQwMQytPsGfmROiYuGeZNY9VOplOJFyt31B76cFVXhJP3XwcpyEMSqdHQ7bqJUrj5I5baszShCG
XZLVVMjdxj8dN+V+NUcjX0zn5WMOl9Fj2sPI8gtQdByypZHFU5stragrlmex62hvbOV90ivRWlmV
5Vl6tcPMK+d/YU0EdmT+M/pKV+gM+OCBcvr/WvjogbZrg6GoaqGJk5yaGLoFxHcc8UYnnnPJPRnn
CtcIJmhyzbGMNDiefD4obFuVxWSDX+rTVqcMiUFVgGAD8+uSG2F0k/EHWCCJ+9HrSqnO/0yDiHt1
2p+i135R1tartyqaBs8pEoMnHyJSGuS9hOFgPrzmMd/ijcJxViJNsU+bjTQ2kysbXSCfN7lzr1Vg
eo3FfmlJ589FQyG59wlX7yRh+XjEvMNvfvvitXNARkETvmic+avvJwHDqcbVSZ8bjZ9Sg3J80DC5
KwUHJPdekMMA4Mh3pq+l7tMHLWf0Ubo5Gy8NJZY9bRdePK5EuCLb7NA+rDziS32Rqqwmfz7yOUy7
6S+J0qTc0Drqq4CKyXNVIDQUYJvbmNuUL5Ir6hcTPnttteOj3MQT8j37Hb5Gi7zVXoGJOHrv9vWz
Bza6C3Jwzu3AiWYv3gOdPZd5iNrwDK0fBFKKUxnGDLyO4T5kkTZyKTJVNR8o5FXai57wv+Pv/7R2
QFagRaJgZy74J2/Vom9CU0NbqTXpAtK3W+msLY2LWmJeh1HkSnRHhcvaht+j51FdEDRKbBxMuCKJ
FGuuUQx5tC8yM4BpFSoVbwqyhMI13F2l4rtSKdPmJV/Mvja+uMqy0o4P1HfdW4Tf25+sdsr/1Dve
GQ6ya3w0AHos1vOXEaNpLr6rj8pvezaD6dBWr8SWqNYXaZ86X6qF5cpkQBqBJuifd5bh3NCZOsDY
20xDc/4N0tiPtylMIA2h0vxj+OkI3mYIHb5w0r5MGQefcKexAehlJerda570lwIbDp9ptEz0BBcG
1Ulst36zHcx0eNU6Ib67ueeyYJDvIhLFND6cZQuHz/5UBTpadX59sxbMq7NCCDIesrrWshk4T85Y
+mKfKfelQ0TpnYMxjng4/Xa5xPRUqXON+nkKOBMpX6RriTuT2eVwNL4tEJ1ASoxrGgIUQhtZBVbj
WZ16QEnb6wyco3yHc042M+bJoXEnz51LbCtHScx562wTMmGi+cjybv5oa9AsErdwImFbHTaByZ4g
FBcPi9PSqlABuITKuj5eCe5A0E6921CMdzGaSPzUdyNtMi7dw07yG7+oP1O+4tV49C3aXlBlMCCL
SSbUoJPLTCL+cAv25KcCoBn3sbgZOR43Uawe/CbyvRNJvw6C11cg7CB5/MOiK7CY95bTpX3X31pJ
Q/cawn0qAwIqvqS5rpQcTe5wKO4iEkwePr9mYQck/Ecz+bR3vvbrQ7DNasKw8KxSJWrEg23pnLRv
eadkwzuq5UkTJQCG+x2QCQNh/zG5jeZwHarL8qFo/Qpmdrqs3FXs9yAFFi1spu//K3kNIptVfo7A
0ZhWjDJzxbH5xuIaPzBvYK4y5xJLHdEba8BLWo4ZBzpwxfSEIzscQbNqO4awoZfpkaNPGk9ZA6BY
15D2PSZVZDPF4dUInUrVQH4w8vetCdZtvlyxAnKyxlRLsHn6Zauv/nQrydnNclZhV07fE6re6j4A
NotvlzPlFMawMojqKYxVfaXlODNFW42+Pc7kC3eoqvaS5eiCPM+FjLeDUcfhbpTYPw1iVNvYy56P
mqEN9RjQvFV1v9VuR0H45ck0QoqMt5JedodIUfpWszRUDlTbKXgrS/2ZL/4pX+phd+0eidoQZ4dw
pu006CqcyNxBEZ1NfJ3l39bKkVG7TTnE3I7l26N97w4vxNAbLXyRbv5Ijbzx6MOYfUEzmRfnJJtl
/6SoSd9bn60wnBZu6nEzVQ6sA4iYwRQZlC9NaI3RmVfYkqk/OUEDMPhSm8/Z8pKGwBcx/LICehea
UV32eogMExSFGU7KHPdJz4Dtf1B9YLR2j7omNy4CwS0a3XOrNpa8JVjRIZD8uulZ2iE+hpI/J7x4
1dZY6zc/hTttohr/bj36STemgIc0BYJZ83/H0ZNWvwYQoP4jOY/hAZnspaKpDEafGuBf/cIuwnIt
7Df/ZOhA8wg7ScZ30iWwGfJDSRPO9sSN7vr4QqWwEDwSyGeWdPgcBdu1bhk0RNAjZsyxNsHhwMvz
aQqhZ4Ms/UgycxQTY1Y87dxWrHHnRg7mM2Ttcp/2hZycUb7BIyo/1l/W4X/AdhQnZXCVFOVUhBu7
5T2y2B4Wu/eLIVc+A5bU5eAFC3OK330jgPYClQoh76H+aJN58vcgh9ue+OacudjsqGVAyaawSwWU
dFKSvOzERFn1SoJCDaJ8T8ZFaNt9uBS0QFM/knsLBsxI+EKxzEIGV6+CUfE2bcCke5Pzd/K+oMfk
p179F2Qn5Hz9zUiwgdj4dEyomA+FH+WD7+rddkTIV184MUkVBMTxS/2dt2mZkR68c3MGvkvPJ3Kd
A+R08OhGFd3wnqxZYuT/FyJY6Dl+vj4yXkqKC9cEpAMXVs8vaTPF2V25nfb/OC+AEfGe75D2W5DA
jYTQxPEFMpiGpajhmA1CYKMpCO4rjWxN1+tYgRA4R3hx9fvgSbbI/etEDlKAR+UOvE4SZPUi/dVD
wYI3HUejEyYk34i16IYzpSt9YOoYYSyNFUV1rBkeESNynnP+txQrtYtNRBhD7JimE+WLcSsnPxoV
1u9A4BmFC7AIMmg3bmk/bpcAx1RJIcnWW5rx3raGirvS/nWeeiBRUY1dLnNcQ/y49gKssiW/N7mZ
cUe4ctNWGfG5zTiorVG0lmF3L9mO80aVrYHYNWhei0BWSzOZYXXFBnBgGmE402REaZA16w3yf8eD
s1VOJaGpfXhA/Bl3BD0tPMZ6zTKjNdNaTm3N7OL14PMYF3/24Eik7TSSdM94rQkEGM3njnMNfHu8
jCcNBQ6VzoBqmsSyPOqfPOJQquP7nyPxLmEl4nyCh0nn1yvI7NnSUH7DE2pd9V5IogMnXRf5VwiJ
rx89VmJ4O3Swurm0nSAAds1wkE3NQYUCQ4LPvOPqO6oCZgX6UsQcHLo/vgiXt1Fl3BZob62xATS2
K/MJg18BS1CYCEQXTfvr0zzrhltr1H/Y4rR8Ek/nbhbm7fSPrpIgDJr8hyWlIuxmPkYmxtEq+MtN
rogUXyua/nLwm3xODAzeEOQ/PKrZv8Dcz9rCA6+G9NCR1Hcz/K6vdHhHKiwgX4oQOCaAmbWPk0d5
bE8lqc1F4YTPGwuMQ8TYnZCLw70QjbJNgwDCZ5wK9dTOaYM8rrcIVS5idlk7oIe3yv67mzC02l5J
U5HAC+CQku3IsdAszBRgqy7qKz8IguEOHuJFA4b2mc9fWIsCsDCn1lEUDYQaduT6mCdBWoyD+TrC
Hfdm9uLlDARIWaDQ0UqC91xGMs1Q1NDTsk4pjWNveEmfQdJP8nbm1n5g+wWv5KkjR6LaCjxzcHWl
OVBRIw0ig/t3N3cDcCp/YiC0egVDBHXn5WfTh7PtQDFPCm8zI7Il3T1rXn2A0U5aCPKEmk7Ft8uY
bKcUk18UJxhDufL/FjXARaQIP82gWfhYQg40mxPvZUYyOXi1nIF9Nc1BQtaR8qFSv9U4NMHU8s9A
OmSRAr3iECvK+lYjTUmIt6gt1GrIyKZCgPBD2ePbzLrNGrwhmp1KubtyHGpLahxFd8L+ITO9M99I
01yG7KHnSkJbbopYVqyADbiK6/P5y+SvHzQ5KBy8EdnOVH03dXX4J+n5ThcDQIN78Pn/LHzvpKqZ
jKqgWzfEsiInii4k7Sy9eenleR7qk+K6fqUgGKPA9fduxbn3gxH2vwqnWalLCgMuXolhBkYxm2rg
ErXK/JGhy4o/2nKxEa5jnNmmv8kLhd/duM9e4QOXq9VSlmgHqvlkuT0QVt2j4WKlXYod2arVz4XN
JUYggMdY10z6gePDXEVaSqLBQOx2BYPIQWMjnq19f564X+7+MbzFMNcIvqWvQdw4OxR7B0W1lnu0
1NWc/rn1b8PkrtlySYICaN4rWW/WDhdKj54ViE4z8ap5CRfeSiNiknPRNBaj1FbB1JsJGLx5xkmF
l/c1CGBd7L1BpLWlE1GE1aDRMuS9R7OIJ2mD3ABYaZ7YBKvUABT2oShSCgS3gJGTWgiGmcgVoppz
ujkBNbaj49zP3+CcKxfgenrhwgwA6H8QoGnYvCin1F4FOM7ToNLPXDIbFIqCVcHv6luC4ADpq8RQ
GGT+jCPSCY9lSTEwmKUm1HtKoMxCv/xrBXE2JUxLePZMrxu6xoTkC7fHjUz6NwuXAAhFvWSbyyVx
AArvWWNiBUnFrd0NbNl5MznglnDSfSIOhn8FUUYY1K4nNbXIoGuKGp7pSLAoi5R3K5eNrZYHq17S
v8+Q9nSqcR1I8TAtRi6CAnRV5a8QJel2r0yIlQ+DlzfzT803Sr2FPVMkEKzPbcAmREmN9TjF9XQA
qZqQWfJ5z8sHundL7rF9Z1/Hbtc0Mg28nO2Ml7iOkVxbN8lFjQtnLKUJTBDvt9uvE+4PDxvH+TqO
f4pqVTgDQCNywPGugohv6iJsA7HBGUCoh2MqyWSqyjrB09r1EltyVKKqFKRRVjnsQ/Oy8RKTabTH
HN/ARZ5v0eIuV9YRC1jZYGY1Pu876Hd+JjziaJlCYmsD/cOYImbhQDHu6yVpf4FVqq4SxxURd1Cu
64Wz9VtAhtEAV+Ut8EAJWhjUhTm2hAZoQpQVa41HwxcMqoOyAdTew602HbnbTz066aoRKr1P4STK
YFobux03BUmGYFZIDcUa0WD2bzq3KaclqdWs3qMqjyDdp9B3gapshrNAiVt7lxMnrJXILrjqmUM9
FFATVpDqq3r0z2rYmIZwTSFBIuCz1GR/Ig5t3RHF39U6yDLGq4mrSc5/QFilQ6Dsq98cVzD9aO/X
6EsPc1oKrDWwjTEucS1WAlehlucjodfFa5VPJR7KMLTHCbLwBuq0Anh/y0K7SWRmazZ49SQAo8NM
aN8XlYE+sCQBuQpEM+XvSkZ0AawDblOasVOWvZzUDnES8q9G1UYEf6/TggFFi/qGibMPgzF5bYCH
LYSMu0C7gUWswAM2YZqrADYudJN1WGXrxAqaH+NJzwz5O/aviXG3lI4xORdf3pResRzIkLiksDMV
VDp43BGGnDARgrT27Hx13FQaRIYXvbv3zu6a6AU3FcAA8LD0AEcWz/1YUNSJtay5t8eOfhrMc6N4
ewSPk2KZvPNI1xIWwyLWxH0vIaHdtnyhmAu9nEwjDEycy76jCy5EaiyVBAo8+enbry6QMWwdMwmr
/XlQJ6cJeZ+wTAUVv8+SPaAb5n9/efa3b5IN35ptb/FyWqIDXeRkSwNNSITzq/v+qZMSaAeBAXZp
4ag2Lr8ON9lvWmjR/eQJFoOntS54N8ky9rwmfgG5xHmRXfZihG0gZ/D2q87QsT6B2IyKy7lky+pD
vKQPrUvjNp7p9jAlKy3+k/Uqjfz47HsAqJEnranfJ7+qGXh1OiURCei8JhS+vLqBbTx7QAKm4l8Q
7fCWONGCjBmwgyn2Th+p7Y3P+m/Qi5XRWaIuC/c4Jh2zDA4xkUgw6DLrEIVzI1U/kJ2yeQTnlh1p
GoLq7qrE9wyCcYHMSCSZvOcc0P/1IM6rs3MlhIfrhcxH/Dz4IRrzHqy944TiboToU+7JO1m0MinM
zileVPLWAPapt6Es8b6iYIkDVY+6KSidqL/D7/jw8656jIeduKyoE7HX50cTAKTB0LPe6B5K1lVI
uf2QYUEZDvtEGVM0ncn009jB93PaWGHGL6sUI5vFLueQq0nGcxnta4VWt6ij2mp2fFVTpp16ZU3w
2wdvU6SpfGzvbAD9m8AfS3HGTf2rzTywJFQ4E+/r/Ec+GXJpDtdTuiWyBS2Zr2tL0sX1pEF7byE1
QvHEQsLumJ3qbH6WtXzAgBRwd4IlwVxA6VzsbgAn82S9VIYHDBJ5B09Bg/xFRl8fTVBCVQTLBDVz
BVwtJ2JrB9nE7qXkmrsHcCeAxNhbpMwZYCnxcVU03xU7Kj6Rm9qHe/6w7HVzYsU5BDNIz3qaX8UD
VoJI8rn3Sk4D2cCf0iSgTpeX8/3O5fYeEWTzaASFCEr63w3cxqQLEVlK7aRw6EGb+nI3qKBqtJb2
UZ6kqvtM9pyfYSe+ChtuHM+L6gaHS1+23i1ZEAI4M0ZJxKbL6NojN326RrQCfbg1/enbmEVpVr7c
bHAhZW6PGvQQqji8HdKgL/ZRcUyWLC6MNbOaNpArMl37d0SqLjHWbALQoteYdLBOeHlpkQvFeWGv
gFYMBBJhEoiRmJVf7F1vm/WIhk4e4WrtDae7Hk8yHASmywuKjaUwKAvHJKc/JfSmkihy0YsooVI8
STOr1SUGX3i62nNNnZsTtjrpu5msXjHUNNqvjZ/Q2WCN+CnJcO7YYx/c8vJLGJh3Dh3LmonfR/Zi
oLvcODmTp7YAu29S7I6oESBJHY/g8wd0+Aq3RhWWrWpmo9PsIYmRQMUiB66MbO0RxyMOkuLjeOSE
Th2bEI260uSElKjiMVTIfSagx2XIb/bVef44lXtUP5wl6DZctq11muau3T+dvkvasBR+GPG7pPyR
oDzA+cpfn2VjsaeVn+ba+8W07n2A6cII/jZ/hGtPEujZ1EY+wq5K7PUs61ktr9neJdR/PnU1tz9A
S5VoYqeITpg4qzstMYO1Q44NTpGgZ1fFFAut2v/AljqSPeY9EJMHUU/SGL16K63vmK1tU1vSp0vk
29NE55gI9AicUtbKL496xj79mx8eM3vphn7tulkw0O3ykwSJ9PuivpY5ADyDljVqcF0aynNZA5WX
ZbKQ7UVwVFZ93sTpDf89zigK3qnsncZ/2ODVK2nJ4UmloTDFLIz1yiO3mNQo/Hpz04vIvkdb/yu7
0bA9rQEVfVSOy9OHiArZAZr50PW6RSKZQYQFduwmfbLXCSKkYQelaoCRRWw4q726OE/23gS+NKKj
1W6skbIU7xgabi9qXil2No0rfmhgeFdEywSM6zq1VsIWDcd4muRRNodharoOhlJqQr2Qqzwkxnxa
YloyqsOkkfArlnWocNfH80LSU0M+GzUhHxpM00Hl4zaX6FRg0OvJZW8ghOoPhXZECtBkG+7qsLmb
gkSGe0JKbxoOq//P9gmKpV8gFNLdjtNiKO/bWjzd79qdN4LeJfRi7EE+Y4vhBSVcg5a8V0LxreB1
bu4twL51NuoQMK7qxMHuI9Ub7SYSsSnw0QhL6rstcDaKmztOobsA109AJpwi4bFthtYzOiVSUb7N
RjQD8g6NQJhWJKWeoBpYDrIEtqHAOOBay4aiPwlcD1sgnk67tIs9cmdam6hz6w2giC/jvtXi6rHZ
OkqdkB0vIMZqfmysF5TkFO5k9bx5I8JUXga3OPJC2OcrVwbSCl8wyK0BnosR2SBbYRasWofGcf9M
TjAyfxcLi7qVw2Kb+EFbZWM6M3vuiMm4fqO/ymDh7p8JQ9yoPGX5M+Sx/kMLKEM/xIMkJP+m7hIV
BsP36xHL4QaBI8v/Fd15e/+bw+CQAp6Pl6pIcGBbsI6b7t6dV8+16wZixqVolup+CLJeW9gstht0
Tn7AV5E7oX+EnXBoegrkY9AL+YEw3BTmYBkbyAcj9oWHzQ8pqAG4B0XL3nW5ArPpsMBL6q1/t2KN
UyMNTRaTQahpkIRuh6fTycZ/HOPbOIBCL6JYfM1ZqpjGQg6yfhuIXTpMc+xAWt72sIytJfZ3eu21
AdNqDvVeRA0az7ivxxbcw/lUKXck4/YjwF1oU7mE6vc0xot6gqG+sgnWTXfJKZszsaUcvPisgdPC
jrWN/n2KuCqQTZyqYKWsvkTrsLf+LyoUs5sLOdSusrp+QblA+0iW4spxxQOAH4OGHX5GXp85Rrdx
V46QjAYbde3vRWKpwL8H2dojyt9pEMNbtZ0bvDy5aiDB/ZUfvE+PDTGxnPisIV7kbjcf4ya78IVt
ctAqB47plqV2uHcdrz3WGrjvUtvCfVufcy6rqWO/K23do2skgxaLRppUHe/zMsDIDAhTAyGpJ/VA
xqrOpWBsRS/is0OHa+fJ72r4GZAyj4TRIO40emR2UrD3kmz5XsjtB8nvcHrO0R9f7UvCM0Vz3sG7
ZEiPQU79oOnGAkT9KqNocTYb3y4hiQ+PdE4S6+Fvqs6U+qUe+SOUUTWqGXRxJIqmApvriyyPcpPB
c0nbrMn1UBXqR3yc9vBZO5/vZcnNF0fEDlrq33fyt8NBM1XR8luF8OxQBzhPugoac4h81GBQ9e47
gZ2iCaXIHAnepqpjjU5Gg2krhG9OptyvSlau2zqzNTiZTMDzZZtFwKZDKjgRKLn3K2kTl/Otvtap
tYe6yD3vGWMLfRijtSRpQ6kBgv9WLDuqtnpxOIeXUpSxWO0ou3RpdVtSNxzSBUxg39ebV2YxoDOL
WbX6C52jv5AFAt1aEBBD7qM5XfB1+MD0ummgl3g0VI3cyPrszYtTCDiosfJ0Uto5fMFUWiO41jLk
ISTkfou0Wg3PxUE4a4THvsu3zkSV9JR/Ww6HjfJSA4avO1BhNsglFDQcU+2Pu6K8XFDTJzjBThOe
3n5FqpIqJwkT1LZmE+jFEfE1Cf14cju0lhRNflICM4r0HINmqbp4+kjIYbBPrtc1hWjUs1jw2Njl
VGlhGaS0n/Vib+i1P0plPYlTIoOV1tkIgH71/6m2sL5MPF6GeznitPz1rBLf2z93JziLOZK7I836
G0vpybGlIrD7W5elSa8xuLzc2/XElx9ASqTUlPV/6tY58r/TSs0DZixPhUv5107iZPFfieG/YOk/
oO+OYc+Fbo+5DZJgkn3Rce6eCVZedDBcWZoIChtS27bexv4j9NEBHPSbtgYLFyyta5u5hVsqeaFB
84GlRuCwVxOJUgGqV88RBHZlKt4gx44bJdxaEa5f65wpbNStZpaDW2i2gOrlX0lwAsFxln2ije2p
GQZGjEd3zUljoCqDpw0iVSXAtaE7VBSD1vwRFjfIJtvkp2Xy5meShLF93/QePJ2zp7vjrctyOSBj
mHcO1S0INAPla2DgLSRih67zkl9juB6V+Lc6BBycjurMBa3Bj8+5On2wDEqqzP2mBGjgLJr6YEbP
NurB1vExbbHw70sahlMwiU1tli7sZVXWE/5fL+SJoB9PEqgerRmJEuru2hLTVvTwSVXHUWZqVsjY
i1FxggzJVoyfrbZcNPv9rY3EAIb84NgQOZR8ToRGSehNtOGcAdtoabM3U2Edm1cbS9vt9vFedRyi
QgmcbuIJk3qvVQB9hpWlOWu2UMGDOxj60gyLpTHwKduzF254KDJvCIgVAMYcqmTRj/YLf+GOjKQJ
dEqJztFAV4ps6qbspD6L2q2d4cqZi64Uh+kS/mNKYCmBqAj3ur6g16mXdjM6Z9NQd9Z+IvQRTr3F
f/tx14CicxSFWS1yp/FqcxKr8E09ahpzPKUTo+m0PwcFyQXuk3yvUO187ZPHnr7HhnyGAkCsXzMb
vw+ruQLMGmd/ybxZmkuQohXgBUDr1HLKTcmSysjg8LByMArNDf+CGG2xipXDeW1pdLnYQOoT2NxC
IWXWCdP0v07gK6KTFbK/HRWMBT8KZzNQqP4aUqu4Z7HRInrhXQfbVxnUrbmUDYzpUF70G/0F2qGj
QaBziHZmaHKR444QPYZhcC4Q6Lhakz2WcYvHGtgkHfjIg5FoLBXjFhN34Irb5O9tKc+IDwgP8v2q
6Ttcs9BsaPEsF5hR2/BzEtwv9hrGduiX/T5Rb6UY54aXyQkYWlhr4akezux9Ox0Z1CG1CvnECoUh
HgTKQm8d7UH139+kYDrCrVUSQd7RjbypCNaNlSdfWoRJy36boNV/XLKz8+24xGrEWsV02ofSAyvL
tuSHksoxzb8IP+rl2F6Fi4r+rYwIQeECzgza7KykqqzfbJEtF1PkWIoctgO3J1wOqwhjMjuuJexA
KFvC/5vKUYYHQZ78WEAPmnWDxfKMDZHyERWNnPLaVA+NU8gZsT5woK/OIBJ1HNqavw6SU+N5VVMi
4KsVYil/Qpf9PBqlTgt/28M30TT7svTkeKaIsKPGNUjzRfQlPnpm4l0nbgUHm8/mMevXWmXspM+9
uISjLBezvBOz9D0pPqq6W25+Ne7B3pwVVUMl0G5KT95JSLie2ZIGdGSgyXr3xOTFpTiKRcHh7msR
C5gq/Ml5vV7NeKhLYem6P2V/Gkg0QWc1PAXjUHDFmlaiTrEZwde8r3ft3cMCXhj6si1nQQMilKdw
U+0olTBxr4voSuWBZ0mvqTLaUeXIjW5GohZ5gGHpVmsMyVs094I6L8I16wv1VSXyN+XLEo8tz0/O
q/6AzFh0ZifHyeQAPwmuovh3/6SZhb3hXEP6C+8W+EICZ+C+sdiVL24xuqEGpX7BLhdVSRvw4CUd
0p3mmLFB8nW/QIds2+0Hk+b86AiVBdIgQCrdFBkLm9Lb4dqGTsK0vu/iz1gkCWadf6ViePwR16D3
frWz4Jqu8A4Ee+WOdp+bARhIpF8/Te7gcrvS3bIZzEPLji9eI+EcWS71jmU50ffzGvsdFPER/der
Yfz/iopNDjsKce/XDEi2trEeuE5vgtEVEN+mVKgAB1TKoqwwiGgmQBRxpNPT0xn6Bb9L8mcH9b9j
E+2XFcEV4lMnxQVhZgvppNjKeYU7QgmZAWiXgEDPrXW8XBWDzcNUPCBmW7ZyOo1wR6b1htiIWRHy
Bi/CYaW9D4SbHfCHTbs4DwNClf3MHhobQqFqp8TAf2U11PF2YmMDzrub4cBPdm3v/GOjDZezy4XR
ionw6uqZ9cLpZvDxqEpAXie4phxmPekWbqAOo3Cp8oqKKDhaTkZcvUaQJd4jB9IV6KKBQymMYMX5
g35+9lKzLwjYGb07zGIYWhQLYjxqQYORbGM2C1nzasP1HFWaOjIwm9Tmowcoocm5s8dwaxaXLZzW
3r8S9C4cbGuRC5WkkWFABB2OK24CcyMyeHgiIZrC3BxHLAfqQOMlr6x831AVJUO7/wvlS8PQ0syo
V4ZqsY9n9dfArOJD3FBvzmdzAC3cBRZy6yD+i/lokdzxI14LFXOqrAUU/gf+HdNdPpxp6F5Vb358
1RsyOL0PzIgfsCA+36d5styneGDtUvwoDtrD1Hp8j0S1X7unJ0oCF8HtktUXTBt9VMoFKisaue75
Q91dTUSWjK9acPaMWcQrn8LbTVZFpU7BxWT7+lZWBDIo5zcZjpec7zTz7ljUSBKBEf8FQ+Fpx8wT
Xk/jzulDbjDoVlJiBuwcbHoqiUtPN/Ey2goMH+mbafVuERcJdYOR5pERjoaWhEqFs/+uCRJzqh/w
bj6p72PpeXMksh/ylNod+LF/hw6YUe96l6rnuKNX4hf3aNtHkmLY7wv+mxdaeEAJGoWtcuMpUxmG
7rbQkz26VydhV/0pRxWlTp9WNEphAiUoYfAnPzxrXMJdiNld/dadDBdvK+M35yGVjh6tz3fyuZTd
CfjHQaQpZDShK4edejmP0rtccKEyY2r3DNri1zfwlsBxK485wrTEGwj1VSbuhHEEgGCz1KPvBx/7
G9TxhRFzuQnq995svu+QAS59UqE5/9hyuXhh51Ij3HQl/onXr8HeTtVEPVRFmjECUNUudU6/F8FX
cFXDZWSxHVjU36/Rbe0oDV6HXmldErnAtjx385X/9Upvp7rzjx505sPpEkCuvApn0G+DcApTREhQ
2Jj1xgc5PSpjpRcXBLvt3fi6fpU6Bn4IKPdKbpyES1R76zwWJNxEILv8UCBxfuuezBHc+6YWVkGU
69I7faKT+LeX5SUfq+nsazubGx9uZY0kzp9BRcI9vbYCyedqUSXuxgFoKHRy1oQ5YEsHDWKRrhVG
CqC8xo61rlUd5cD6ilTbRWCduubAtYTTF1rR5H76Zy/1LRDdp9RZL9XGeJc872nfOhkJN7CGcEpM
agqIlpwsEWTNmsRM11Tdr4aqzMK9q9wAiXhsGENbyEqnLkA6P3hF8gD6XtCaglOQZzcrc4zTgic1
VP60FGKl1+/RReikYqp1D5cI1MlQVBrLwkMcu4+PT+J/p76aa6GM1Wk7vF+xnentcXS33QY8+yc9
tTk/ijrcqQym+HrWtKWNo9K55z69pPXJpKqV2AWyTZwA9216UkE1YlcVU7V/pTybISfRHM4TizYp
3ocJRzAHbWOOU08WJ8aFOQ2JKd92xY5D017Xgb7OiJSNagRD5osQPdiMY398ftZIKhJQxSF2t8v1
1pdHgkUXXX+KXZ7sPZjAEW7CIi+AHzIxir+GSRh7qfnP5TAcIdcYWfm5l4AZ+rr5zIIF4dXdCzuE
98R65dbGoIr6p10y1pFTu1VTzbN/T3kXc5MhH2Bmyjq3sFZXfdGt0JS5znXqF+l0IrQ3m8TejRTJ
bFmDxsfRyqx+8gXTLEtOJa3ymjSaaxKouqAuZL6kEiPdjMzk+vJ+wXcLgspT6nz/WB6W7ci4r0d1
m0dIULLouI2szSn8QI7UGI6vSvsw7V3W5ocvd+AW9Trw4wV41I5MLpfwQCjd7n7V20EzK33lmWN5
JVCEBjP1c4IrOXIvwjgzajQhqUBlxQ5ntnelgwIYPcyO8d0W54A7xShTyxYBUup3CrgDzxqrij9k
n1YNQK4JU9bg6Uuj6tFWeg8p0sDTgwq6xfNFychsR8VG1eicrq/IxqlcPc7PHt1oZDT9saRRNtMD
0cWUEzqSrTxPVp9BjKpmBdQfRbwlhaykWBWJIGWq6vrwmBJA+Aitg67dSJi+25UgK8GDGgtGxEOR
DQ1por4RBIeKYpsrcAZxwXpVbVLkEJjceW/gs8M9evY19Vl+yt1gc1R9cRthuLZrAWwGBsOXjzEk
C/NeOUTIzPWtDWz7YLl4mNrkZ9KH4+JdkedUjWWK9GhTD3c8KTH+SkEEECsRYVWbc8ioTW0QdPOJ
j3o32yQypN2+XwDfmGsQBog/nRWmXvcdRjXiiKNte8b6JnueCQp+ldOaRIwrZeHTndfSOaxBfcKz
MJBT9it/TfokRhKDW0Zjg02OcJAH0VQmqVxWgyK8aESPAzRHNx+UNyaeDgEanBa39MfQZhgfS0FM
o8H6as5Vfe6KOgOsloZF/KikyIdSqerdQcN85zTrtXSa/ZRPFxiCu+HwAlW20lnPSJ+PVB5OLcpI
ccaaIbNQKbuOhOLDjoXXJ/RB+ig8sENag41eMJOdUYfj6zk1bSsJf3WKRBm27sSR8E2fYRg7+92Z
s9mhnMVaaDMORy/UigmN193nvGI4yz2rn4mkmbub+kP2QmAJ45ealuKTI/Rm63hMnluJtF/x+jXf
PRiw9Z9FplwlKHJk+dQezSrCA0M4hsosppo0g4Vp9uYNLTJjt6BwLv0qyyoPd7qrXhtnPC3T58AY
PRlh3cG6DzxH1Q9V96Mkl0VYhnSMr2NS1nh5qxG47aPJHc+N703rYEedeDk1cyzcXqzubXcsdSwS
BYUDll7my5ClAAWaCxR8VpY408KzggSyWm/S49XMkBGL/OW5KWPDgO44+qsAYLWmsSesBtY156ft
NtDzJTMvbwCAUikpKpeQWXBElNuaFkJ/QeRkFUF0w2z5YUUwJ1DGVm8NKTzhp9ZdzKobN2z8yit7
h0l6h1oze6W2N/ChgnY5MEjYLkJ7bO3XrRIBl46O42Ww0olHVVykTSf5xF6PcZh8Q3UFvvN9QIW5
WTTbngDUGAEjhwDDoR+3UnziMdmU2EP3Yevw35xUCc3yMCue+FZn7Ckhg5jrqXd/dQ+ZAEuqyXgC
2f3uQS5SPcajnF1300/HCY2sDXw+qPdLDMcffu9az8K2cqLSrLQrxEg18rXlfHGTejRoCUCGiwED
msRrVlJ9VsBd68Eko5L+iWUJxuW8kUzxiJ1WrUwk0uGes0A8mrR2fN/PB6MgmxAM4Td5obz9+p0c
iBEGaGKPsSq5le9X5z3a8fUMCmZ1fLK2aA0SotoyC+vWk94rwhjf3CYSozasdos1sTN2/ok41ouI
8pPgEbMYnp+No+/6mj8U5pUVcwm+Arx8qtgSkMqiB3JIG0BTLVkAWCCposOtraFzOv13eMz9KJd0
Vl/+q6bfoGFtGw3ryC2UKRVED0GjdLI1FKGBpt0fvKUS4YTEuZ0AbEpeuxcMommrByPM2NzUw9kT
sM5Js5qyx7aSh0skBlBoefEtTMjQfBKwRJQm1fLSsGcocHH97YwihHdWodl/eGrOISO/la1YURIy
d5CIHx2sTqTG2ZWYC2hekvCGDUEOwvx7KWOX+dx0AMddQ+6wJaTupVdXhZmVaMwoslfKWreq9/5I
p3ad+nmfgNgObMjrYcaPaD9CqEm8GPH55ugMQVfR+fIpDsLGxkyTm3RD6ckkSEwoqkIJ6Ls9sy+Z
G9XKqCoQkvefnlBm38vgWAfYVubNDsaZ2dQ/9Z0ZQHQqlZJOkjIbH13rEahK+Y/qYQANeNcTyc9i
JfBkPpLPrDMJsCcdOTyk5xoMCbisqNp4BznKkZ1Xyi26k/Sq9ubY9PoNPLgt47ITVXMAeOWgRs8e
g2tp4cg8lyLCDaSMpt775B3XwMJQB8TdUrloegws8B1JiFuQBpHpVo+oARaDNMATelNgnIpCdmKg
Uif8Cu0n1nSII+qWN+9sZgvpRGbeGKHfFVNoBY8MwOHFMfyxh2pPsRHJSsCSCkTOGxQFqeyHMO6w
jZ8nser2c/7helcfpuEOD4/02P8yxrQczxxbzwfTD/ufao9k1q72khZv1gdLX1cl5nY5hu++a0j3
JO17fWNnLx3tJUxKnA+fl0Se4HrPTa18quT+09CPwyktbTcFtP7m/2r71S0CRLTC32IgsU5ICLQO
5mBM0/a8P1WR2uLeijsFj2IoGZ333rWw4JHpRIwktzT+9lUn4NrWzQIfOcBt06UoAJBEi245V/bR
q9bxhdMMat31jaBTxGVvWBZzwepGXij1vKzp1q15x9aAT+1vEIKf8pfdODKL9Z9o7Zb5QVwELCxe
E7P4zHY+CcoDcVtEBJqFT7Z7y3eagePR9R5KtzR3rFTAgR2N9ToRPs79NWocdnDITZoz/B6yivY/
3OO/edH8Lq7XWpYd/+zlCZR40PKsnrxVqn2o6bSwlpCsSjJJTe4aMIArDPbqVxrxTmyq0tVeHN82
F1whHLpP7RkbHvYoQrXC9bRtkF/YGPz9fm023M2eplfsUgEPmRhmFRah6hK4SLr3J4xo+cHeAOge
B0u2gr30qiSt6h29MSrmDSzjNwDHPtA6IUEq7naJOKUUOoiveUsVb4zJye/iPY9BuSbLs5lVk3mh
4XzUpR0N9LB2cTTTyx6j+aPYWkBWDcT3WrzqswwaYu/5QwgrBlfwlEY9D7TsTwKRD8jmJk5ODMdh
HCjw6dLHNVUiiLNrUHuA/ShiVGFC1txFMBuE+7MzV7WiVQZ8t/B2xqV1oiWDhWlWw2J6uE8J7sgn
70qwWJGZeelBlKh3kbWOToshLYcx0hvSPbFKYblXxkOSFzyBxAPjxN/oDM4lm2DLJBpHL4e2JgBr
K6nUkvPX7bw3BQZ36uLKI+KF1k+9JC6pHJ7D4yM22iH8xqtCstsm/Ri0Z3KJSsaysTwa2vuA3HKf
ibfjQRBIKTL1b5qCeE5PyW5gMx8iom4rWwMWchmrGc8fRQ33AvLdBDB/3NuXyjUqf+KafFGA9XgH
kmPkHypiijhQKQdfHLs5Gk7rwdPJ1t7nPuQuXOJTRiHx2IUyAlPO8o3eVY4W7El1zcy70dF3301q
ZbU8HmTH35GGxJ2VlXHQTUn1reQTxm5HDNq9mYLIfo6hv7C8GyoxdUf600ZAFWK+RrGJRnVHjKtc
VOhEWhyJOGlNAkBhoP5o6N0soUlIoQqAwuqkSS0oc38TLq2s583wv8rsaqcpMjhupSVbjTXk4Q1M
6EKG4wvNr6sEiqUTeY0f1+Pzc8nhmf8ANWDbaaolECByplSQkp1SAd317nDIVgF65CbjAVSRtsGP
oeBVWbJrLK5sOCbU/Q90HLXS59ZddKZNRhDb/Cwy/DdWDw/ZT2qqH6I62V1atNt4OA+zgQahyQ6Y
PE+rkfI54T8c9yHXbMk4cG8h/DE1ehn7FxHFWb6aRlGOFikX+FwsMxZF+o8nd62zGVPMBDx+qfj5
0P/aKYP2rRW1D9IUgzVM5YYsdpAqZjLtuOzsmbiqodvW3e53fpk7VnMpuD1YRGTnMm59fIXJfs2i
XpZSm7ecHxamZ0TPp8yXrOj2jrSodSu0Watk9ClbXz0OxW+NCAPv8ojZtqN+YJZGqc2edp8c/gk+
BZMVlJYXtk5iVsF5eQ12mnerd6vIeLA3ggoGxnSGPlNJ6vV9obrudg5WT+qVQt9t5el3gsAkn2qf
45vuQk1ky5j5cnSd2sl2FLwT3FyM6RAUF02Hr3MLcuOgrfuExw7LdjD6CsDv5KFW2sIkCL/S7LiK
OF5YVHFy/+XuIZuW+6JLWeqfgUwdbPYJ+lFYf6baMep4hh7UU75F70kc911Rqg55yZVc62yYoF0I
CyWUjL5APPiml2hlPWB0aRqTPDf2SQWcWTqPUx5zzvoHz6vm7USQNHkIGcFC42xnl8rPZwg9V6gb
L5aQaoaKt6fDnQOO5Y0EvvZzlZ1bXwUcB8W/MiNNHIBZUQIQtWKo38ypnW15Q6Oif4gLy6X9qr6t
crJaJjbD3r+1renuCV1cyzsokc0HmD+EQ5ZX8xFECGNdQmSl3pUjp1j/bxniJpbK6sBxHAuaCiXY
iGYUo1Xfte8r9/yveX02jKz4pUYV6AHf3fT6a3xIkOcVajAW8Vkxmb5+dUoQFQ1CnWEGz8Ahzk5h
3P9f9IROtsbC72rN9J+h6HSxAc4JJM2IejpF4EXQeF3LdpLQ1apzQ8rtugs4YQ19pq/wPPol0Y0b
HK650mtVjCGUX3M8D/87uwfwsp9SBonbnU5eXgzVTqeNgSpk1B5exWOq+YoGlrct0Xdosejj2/7T
Ze2R917rQR6dcnbqj3BpW3SMAWAgaAxvKT0pseV0MjRbB3c0ODG2+KcM6UqdAmPCCcVbPIi4X9kq
I63rJmH9tu+ZevgBi1+a1hdQG1fZHr6T/DRXS/jt/aGk/FgYKM7fUb7vBBFwno47zZooev2aGuVs
3vBX1TgcB4VuE3kENpuAXHDdQbTzZDMxLnSzcAhxOSyoFO8J2CLFtkBEpJ/0WWs6/KqTr+wY2C9w
NwQpsk8ctu/9eWIeg42cGFqVfFT2DZLJpx5vmSFpxsEA2a6iJ171m2F2cOkvOdsjPVe5ZsAzvEGm
Lw6WuPcRpm/Nppb6Fzg1UN/Eq6mTrs7V0HoCcHsNvRplOXta0soU9koPl4p5aaexHZhfuWyZvF/2
LdjS0ItPnbghjIs9cgx1GyaYYQTOX3Y0RyRgvBtozD0+I5Op2vffVTMDy2OL9DbeEjhewup1ng2R
e+E/gYO0RQmEImVJ4HKVHV03chD4cZkigajfFDSSicGIKOhTcT1qL8mLfPPFJfq9TdfULNB9S9Qy
DX+BazSCHnPKxvKpm43XUz4+WddSbJifUbrbd+tFs542bsWMyrsZhNkD7LNtDhKwufqshHu5bbTp
YKBytzD7NmVb7+hCXaQMi0nhsi/D033P0D3w/67mbhNLNCMTm7B4lznRyqOAD2JmodapszJIB0Bg
u5LeouSuynK07K+hCU90VSVr5dBFHpMEgXVUDP1UTRH4U5nWjexpsB6oejJ2zWL4j1qyRTKgamJf
yhaQZKXI37uO7ZsiivZ0CBdtZJlHfmHwDQTQDyuL5H5txmlqU0seqhiRg5Kvtft6TrbURUe1SByi
1Uc1V8y6zpFzxk3QBqId8VRO+oHYBjLxwsZ5g3ksQs7toXSi+0zJSV6t9DdzGfu+LNxQsGxNse5I
vZ8E0KAQaRE8Gyzjgjb7+3c7y+8yHQdMi4aqhOCS/C4tUr7Jw8zxQ3zgH6ZVqgRz7ZmW/s6kKR9+
CoGpRpx7sHLhIpEyuDG5RmGne2vkAKxKL1QKJLSRm94Fj8UrdAXX9nIlzjf0a/rq3pFXLsoMD+bB
dM7dDw6phQFfWYGVr+SKXXhOpoLit/XolyK6VYHWfsLsFdL4lYlYVdPVwAmg3OhgCc9NMSKqMGcc
1cMWLXJ2pKrR9R7ZywJ5pRbeOFGs3Ga4GoHf49zTAkXjeNGUV6Hwe/Fbw8pF3ps313br5ph9z9Rh
NnQidkADSCJtEkyKAMfRWnkcYqoZozvgi0a/uVklPy5NcXmWiCnzm4PMHthYwplylLPlxWBSsprd
PZreFPos3rqn9iwAWieazPZVIoqsqZA9YPwFvYEUJ+HMIYwcdTkAhSZBPgd/ZJNXyLD1gOAKe8a5
BVCjfzqC5n+esFHRYqtJ/rmqL8oSLbp2dtkjQE2r7Wal+SLu/gZfQfzQcve6auBIO+B6xYUhWoeJ
2pkIWsN3aXkofuRyWEhfiITdt9vvQxOj15Oc8jQciKOVA8CtQZGzDgR/M7k6DAluCPGoFr7XYxhG
wmoiUoQvtJAH17ygO0OfnqZiCnLW1eE6I20g47LqinvXjFo/z7k5hciARMc6lhHVwMQpcbEwGwbh
o5dokomVGUHpveoUupQtvKfvAxRaoqTVj4Vvo6VCB+Pqm7l6IdRFjA80eVeBJb3hAw21hevnJ2id
MZDNYCZ6wG0L+PbXYVLuxVDwLLMtRUoe8ATYtPEdbylWm3xnn0jqgR22QZ4Ry5BznKnSnNH1qnNE
xykWfr1JAt/EXejnYYQfMj2xwgR+/BGzk1fqP3T5PQxnwYHkVQkypiqpmswFrZH59z6OPRACjuYU
lNKMLvdKdE7kxS3pxlznoWe6yrRLOUCZmNyzckgSB+Zc3qrFEJShk6KVqSV9v3+Oc3sKFQSVF37Z
9D2Wo7txTd2VYh9jUO1JM2VHn+tOiJjEd/raSYpzVlJpUlvRDYnjZzu15ZSiP4OyEFXueFHTmSLF
caSqGIEIR7vC5o4M5d7dqPUHEPjgIJysQNUxcUdk4cpvfPFsYuAIhCatGqmsrT1cGbvfPJyjss9Q
yqSiradN2bq8MACbzF9Wu2ssR6pTHKh90fCz4TmjDzLtZnLI5YuH74yh0vUgbM1NuEgXcVVcTeQL
+YClqoh28vPICegZ+RNK1y26wVpHqdy08jHdpVhvMT4eFTmWTIxQTYZvvSYhsp/5PBMhbACo32NE
mfR5ErjEg42IvPWKJcKqGOJH3WXjUHnQCtSXVOzGMpFmYL2fzQmKQZr9OBUe+otI1jCTuhcoTNy3
lHwmmPLaOgdn0/xkGApGz8dFYISTg4rAAMa8w4xRQDA7fCkCc6QDnK9yd10tH44+
`pragma protect end_protected
