`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
GtonvLyRIHa0BG5ascvXN09MZ3qOiFCm0qhQWasCekdFVRCizFoeirO1cOSD3S/L7XBtqzCllo4q
Q7pZwE0bdQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NcAWItlcyJiW5iNdkc1sQhABTpjXqZkOrg1X+Tcfgn7grREOKMnmze0hKfPSK2fx03p+1DXa9nI9
aDMO4y3pcvrSQRCRWXgMFS2qba1ARCCZEOEfr1i6f6+Nx8FGN5X5I1YnoGroW/YZxqunrLG+EqYi
XcxUyjBIkX9CxLSivhQ=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LPH3S1XGG8M+74c5vorJTX4Jd0Q7p5hXR2nHLPyVATbLKyNyCj3u2979H/5+r0KMFY+Eci03CiNr
huLATC3oqO+Ri3s+z9ShUHH0kb+eyBSFWWv4Vz/y3dKeMo7xd/qiF6cFD/jwZmVC699OpPLFZ+//
+v9QSba8dbzt+SXEN/jt0+eliBPMdqYocom4RnNiRzWVLRpczdP8jPK0iZ0dswvulkciexDQ2OOo
AH7xVOxZOGncQh6Vnj6rFermvVKMjP+f3wo5tFO3kt6qIlYJvlMl4+beZEF1FvA7E6pKL2F1zinI
FTyZEqwMwZWW/ux/d9gBr39V6BUQmOQXaUku1w==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XhsVvFI9R4kEmwKEMm1/ve3kzL6X2enhhJxnoXVsTfGBwYA297bpytmIip5AhwFQisRjBoqJ0K8l
8Pn3j20/SKo4hFrQQGF0dNNW6natF+zLk6mmfJ9vN5kjz0dnY6GDFbN+3VxaI7EfmTameGip8Srg
gxxI126PbwVBsgU+CTpGeuVit895aMS8BmBuDurrl1wtMGtV+dEhJIRJc0Aq1Wrns6Y56i0yfgPm
51nrGVg0WniIJHCwCd1amAGBP8K+XEMqgFg7Ax6FDLMI9fkEMpr36t/NLdEvEWInQ+uThyiFxWQr
JKb25unvEuv/D0FeWrozh8XdjpoKLAw1GPNMVg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
W3obImnatzWtWQxjvGXfWFuKaXr5FfPdOSZAbNOW8Mwmo4wQnwYiA7HkLDXfdrmslndHMaUxH/ah
zQFKiuR+SbrPT7aIULBLqqh72i8AksoYWph5t+HS6djOrRH3vsKtdR3ywmgroEjQ2QUcAo6U9K34
zqxoj8P9N8GP6+jAQYo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
p5NJqyb9TdyH8yE0AGM2W7x67vL0sjxs/jTTPTMrKPRWFxxZNuqsL6RAPf/W7gzVERxAO3iFqJD+
UoyFnOxci4budxkwr1k61TSgdoxD0V3HQjFvRukqTPnveyj/ep+eTC4LGfMpV/TPdXASgmKbIegz
1MyLz2/mIQLVdf6YMINHpls+EKIpYMQZpwK/hPkYr3E3OOOvzvQxNC9VDhaDMvYytD0fGysZMNYl
wnQ2rJfehLe6ywYzM95pSaORaRL+1Yx2J5fIpMdmGCqTlIRPg/vBGdEvfU7LTH681IczR8haG53W
YAR00ATaZUq26o3QwofFA/jZlZZYcN6rMAOtfQ==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OsRx87MiUvQMyOGPSETijoG08vE4+CeK9YRUiBEhaa6o5uSa2mSyUldHexlwxMR1rBWiQ6uyqUCt
nOrLjKhAiPGydi/JTIixYfKsNMv/tZTwiL+UoHRiZBVFKKOx3LAC8mgFXdUdYGwZnPhPVBIrRJxE
Rc1n40BeUgXQa/BvVgZFq1WN5zlUWx0e+VzL4EHCQl8ppq0b9oCO2dY5tSR8oDlWW/ZOlS5/u72T
OBDaxVQ+J7PWFUnUbY29E2dI2dNIjwjCjYqO+AssBOBH6HZcymhsJOjXSsS6xO1jpNeJMejZ9zqd
GqVBeDYMHSNvyuKhK1iLew/SAb/tdD8vIj8Gsg==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AYMh8vGmPAmkV/4T9vXCAbcwNUQ/U5Uw5Swerl5fs3AFaCZc0Qd8qyJ+58+zr5M2R7LYmJxqm46e
wTkAaUYx5X+VmZ+SG/c+BTOKZ03KypVWl/ISK1LXC/o7S+auCccud+8zMCxRUsKHuKYyIw/9r4Xo
hq9KP5hjv/dyE2FloIaus9WXSRmy3BsOrnOz34Y21Q3ThEHJzIUzPC9BzWKJqAiXhmZqFyQNpIPt
k/qfbsSvBqSTLaJSexAjyCb6KJ+cjdu04kb0KxNQHwNLCdnF8ejcSevf63EwGkmE+UzodGVDp+ZB
5rDYdmQGjq0EQCsB9QHiQJ9xNvYS9co+5Ki68Q==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ft/0b3HbGm8+/u8rq/UN1q9QtlQ7ydmhNvkUH1HFaaEw8IoZqW/LGV+djzXBf+a0L7Lslm4B8/ds
ZIPflSuox2viiVlo6Gu/oLKkTEg1tP9VJQ0SBlLuKdd+1Wtm5pN17pffr2TMr03eYDI2Wj8CqIF+
sz9vF9ralD5iy24MBrbk7D1MMaUjK1iYLEbGPul5XaMw+wCbhmYkQz1aq+m95hJ31EOKL5VFcBvw
0G1ICvealfGN8TBm1MOsgcXCDnEIfZlhrRoDLXx1+eTwJ9G46IioWqKUIgceTRCiJ0HPDdCrElbb
sSVKrR1ThH2yUQnQwI9fGdD6wpMKCSYrtlh7xw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`pragma protect data_block
ewowGykr0Xg9OiH+t3U9Urk9YH5VLt5MuvCS8SnVGaxCEoZGzImVQbazF9yODZ28cX/syNZ8QI97
ZgDvwSxrdZZoLHFnOHz83knxeKJHKN96YxgBLfa3ks3NVHgMES/8fidn7eZsXKvjlK5c0abpXfs4
XXQ0fpAi7oCYBd68ZssLXP3NXwfaQkOyutW81AdXIiF8ncXgBW1T6pBU81g87HLIJX5C8URy8PON
KywcFss7dSjGy2VQ8ERqrau/QKyZeI2R4giFolHL0DSDuHNiU+phhVdDYpPuD5JA/35svO74Truj
Qw90i/PjwlMagfmDrUU0Tpe0LQk7MWCGY7XHxZkoDl6Rge1izyJewzVujQBmrI0qy+RDJEj5z0dA
9LJtSx+6+CNbGOmf2MtIWXTa4fhK188DQZFYrD4LhG+4n4LJi0QIKDek6XcN3f1yAn5zTohiYFvl
NDRZU1/c/ZdNmYUDkW1dBclVlkXxP5J+elTF6lSPZhxPwSx7MhB4ZLxRlfVKePzflU6I9D/+jDwk
VYieiaoH+XvOkhTi2ox41yqFEygciykb3UCtLe8Xff/Er+mQrYc7fpYdi35vDAHuWiiI0HKPs31g
z7IkhCdFua9MK3JcBKLU6r0+oQeRvUn+dQBl9D8MDdByVXbDJxkr9T3EKEYKdF6l7d9GKE/Y8gUQ
6Y9tqjGIqN3xmKjcDLrbaVIdLbjJucG/qOuTmBm5PZu2tF3M1OL80bKEt5ATgd4SfgHgIPMaiJCO
3IiSRERpkyKTJx+8Tn7unUthkMSW21KDl14ktI2c74hL22xlaF/DJBK4bmpjfj3+bIxK+GwphtWg
Of44mcwMqAGfMzmzqMGHonqaUd1L17J1CdpEMUXuSKJcoX7UjIWhol0bzWE/zjLqfyeNjB9U+Vg7
bA+cXHI4emu0jcgdKAPzb3T91BV5OLMmbh3Nl8hspfDA6GXVNfj+lGbV9M210D1aK2zDp0YJnYrQ
czysB2IH8bCsMcD1CAb+UM8ZgyTiasgp1gQ918D7DKGZs6tuVx7oEts3pfDrkyMwP2C24Avgm0Tg
UbG/3zar0f2ROMTym9jXxf/2GmsDDW9Ax9PCfN2Kda2EmkQpJUnT+ck88AQdQ7AE78/oaCSoYETU
KwbWQ9BEbnT7VhYFCekGy6KA/6IQ/pvJE57eqdkobM5ZDUHbcy40174kepRvbgOwlA/9h+Tvyvcv
Cq6C4bLwYcb3BmRH6GKnGpNJEqQptyHyScllR+RIYWpcAyQEGMxkCAFVtxzrSD71ge2hm9vmIKsn
b8OrppF/f76AaPiAXdSk7H/Px7RaXuwLBJfg+l9Srdr0UTJ4DNbnEoFWiBShhD/5yQhFrsGt+a3C
fhaGx5x0eze/mtzl/YydWQ1qPPZfQoVXlBpuOVSS8hnrPc49riSI8nbNI4QTRqFQNSpByPhfioNU
z3XcIyqJrOAmRPFGgY83JhOFX0+sTiixNnxHHp7QxB2O7VbMPkAn/CM7rsD3Ui5HAzug01z/LgZm
0buiyV/+Q06+kpDf6rklXjO/wCZ7dD1+8W5F8ofFLd4unKgRPp/dFLcgh4txvZidy0yBA8sqDGui
JWA00SuMNO39Ifn7QbinAGG1muwJeQGAi4EPIxurDSiTYP/lRPDOir68dCLuP+IoG+OxqEg0iLNu
harUmCg1GinrRfHGC/eOjtlA27PHKsjVE17my7hbXG2i1s3uDlYubzrElwy5itowE1ErCEzxJGuf
YkXSMV92WxtKYRkYOS+afdgwEcg0WUY8XoiRE6iZBApHI7fg3DbC7BivKacV7oe9HgWRcTJQC/45
OHJ2/Lv9l64hMQR2Zmv5ZU5BzamxcEbb5PiDY1uNhlsX5jCBGZMGmUGfssyLH6edFYnZq4iZvwuh
o1cUTWkG5APWGxpILwaM1yObh7cSlrYAG6+H5LTDkkajgEDMbrrDyg8oItrlQJVH8TmfNwOkXDhf
HhwDQ9XP1cLDRsp2ds7VyRo1RdEeNsjwrF8ItZBMuHTM4K/Mwf6dbtEc88ZajC7EaQonmSSa14Gk
lcI4rV00exWv0tDVIZmEXY/AxIU/IcZtecndCI1wDRaw5FCrpB1i/R2fTtaJTIPGu/JoI0uTMlKR
dLtI9QpnV5KoFX40GqJnBvU7K4Xu1qkJ+Ll1RyyOg61XvesacoT61RKIlSiGJs38TiG9s0F5iW7Z
p185SgnUqwoTfr0pWs9FQzh8WNQ7K+bhm2SLgYjX7ErWHcrzgEEfI8YZvEePPWJFYau73F0uE1dX
FHrnIust/cuIfnmsUn+bqcHgPxLSdUyP4QvwPx1t98ansHM1tbMztFIaMThS9rgYNSf3Vo3zivy8
t5Mrsi5eZxuYYmcScnyg8leG8pTM8XemQ74aQ8Y2nnYwsmQHH6B2vpocFS6b49WX0ShR48N2KB46
Qq1mhQdRlbGD84bMrXxO0GbPYAhGy8RFGb+Zr9nHmOi9DPBwYqDf8409PyutDIkBLBzjc+ct7C3I
+sAJbnm7/f+p+esDXLJmZdfOrnZQLFtF4qMmBpH7/C0OAnZgMXgmOFWR5SsdxpH6VGjGRf6yVimG
BDSpw6kixaM7W/Ot7BYLoEma/5hBP7eWmtKZtW8OwvAqdf9tATYEQXdhha6/6YrHBXolsgcMnpAI
caz3P3RARzrC+pIi6iuev2A7ENZ4SSu2PdQEqTKJVKRLqVML/t883JXjFa0XLdElT6DuTys4urph
5e0MySAYy/OuD3cDMBDx7r83/n+UnqfIsN0jA0OsMtGKLJusz+0ZIz1bwGEsyemBw8w9V3um5HLp
61AIL2O3gOvf7O4+HfQyo8m3B3Pkdh9BYDMC9MYP2TYn/v7Tnx6zFDSntDNato7+EVSUCGkFu8X3
RYd4T7xIPjTpfMg2WwQUNN4zdKe8o6T6qG16qzIwR+h7yjR6JE1562vgMi4mpz4v2KOZtnXgwDMp
G5gFr0Egv5GvtQYy0GRmcrvybU5HijAttkWqD141RpHEOdnZtoVEzAhtNj2Lcz68z7ywhuOYPdm6
j6fqzIkKKfgmkdy66NfvSdp7Yj3HcYAmNsIfBJ9p7P2BnE9tNOGMR1K+qvIumxpxc/0B27OZpgHD
aBRDjPfY/21fVX5g12shnFEK4ZfkckvdmyuDpAmUxRHsAEfxudUs8xuEdEejs0ciTjTL5MB2imHf
7B68g2hpmYVfaQwJycXbHUDTc8vt4D0hzggy4j0/8IdWlypFVry8ssYGWlcO4VaWKpTVoG9n/Z/D
sVLq2zmcTn3UARzpGL0F2+/+NZGK11fZwFFmdmjkCTXYnGxo2B+46OpnWniqbTR4v7vvLXNOa9/A
FDePeBBE3f2CzCGDjeUPmFMVX4kRj0LLIaOY1P2RF6s7UN0s5t3lfRKvr6a5/S7wo1TLyMkk92iO
yTaAW8dv+W8Yx4/H1zFw/r4e1JcmZ/vFbZvT9hR1NVu+jY62mMgQrph2iX22ACWHuTsIzJ8njAJF
hXgBWX9WS/IJlVgvA0MfvW+/8bIdHfgoSCqVgRQpDxoLsKaS1ucmp2Gi93L0UMIMCKoT0AnuZ6tu
As4KfmTgTCZGrChhGz/12WhnpN61zqzZdU/4CynjHMiCn4oqdjOQXBE7nhQfmRf6TJ/NChebR9a1
Uf3kirNLgkwun7BghCITE76QvGvCJlkUdPblbZgJkKWvHWEJpyVz+f2cDSQkDnLxaLpcQOOdPR0w
GwmSnJFciEJZISiaSC2Ov7CXVeO/iWwykj5prbSf/rCb/NT8KHKI1jJnFvOk716eRH/NPDNr1jtW
kqSDlhyq8wHA6nPtjLBYYjMZ//ZwHJS/eVmky0SkXO68Oh4sWfMqkPDuGfNDkcZ9vJiRPb1RBuZE
CFj6GXZSVj15BH3OLuspLmBrb3zZaqJhDNV5ERAX/c4v/HTO+6+hJa+ir9j+hDnr5bgG4kVhtTxB
F6oEediD6s8EZXQNZe+u0Xr1NeTJ8qD/J16J8Y9GPpukDFO2X10F3LVihIKPAsW8FNdBsbpabXa6
GkEDELcGqimZKA5nrks22yhRHwXBQ5NF7E6FpRTRo5Uq+VaF6h3ZhJ/JsNaSoHMbN3AovsH93Slo
UYjghHws9wbDdTUyUsiH0IoqMHTEPlS7+B2aTpc/ZyvZAs8XHXL9TmmkDSf9SdO7DDvEqCtsrz2a
JzcqaksYlJIPfIaHmAGovbSe3bzLBxopgxZcqeMTZRE0eZUUwrSxs0LVw5nGUw/amkvTFS41PtSh
ZRA/vwgwDpfKbixCxacIodaIBFojFZqYrcVJRvsljTU8BKHK7tgpqkSCpour3FhbcjmWib2yXp1S
Vs2+wbZ/rh8hx21V0vfV2mEC0+FqwZTcV6CZK3P0/8Wi297Aiz69+YIhgz2qP4VwOaOcOSKEyWDg
AkqigFcaNLcddChhVG+CgsXE1Yb9YZeh7hVOUpQW0NGklKb3f8SELX+/64mu0cMSNfuIVz9uvaCD
oXqDvPZoLwW4VZqOC4jGZzvGn+PhwuP3RM3CkFWSo21kkMJo7cDSuYHS9FKAxOGAU6nZWSpUuIGv
X2YjIuBLdk9BJDn1Jz/ek17c6EJWK6zgJVEBfgYLga0ok6xDFRYHQYqtSC1a2/KwJsSXU/5WJ0Wn
Y9362cWe1Z9klgrKM0CmMqOqLXQNeHwnUJe/yrXLXTAVa75dpRjp5lvnNBNu433UTDcU/tSx2M8j
TYltN/tfsCpg9QFQ1rBaDrr/xH0ucdXv1XFzg1Q5FJ8k42ps8I/CA7lwYouzJPaIzapQmwINytFI
LkbJ6A45orG/gpv5bcn1tOPlMVFxXn6+ic69Ps/k5cG1G0vXiTHmtoWKw7s/U1LTTgtL+SXj9u2F
F0C/wj8UdRBBfKuMn8NscynMI45EjOkQL02vXGrluAg7tgt/GKMxWV4CgdYlRD/NVNZmM/pL7ZM7
Hq8fWKSeXkQAql4MNShr++ksNYZ7tI9ZCiCAJoauaAA5tGwCnvd6IRW1H+kQlWi+1L6B3Rg3GBew
50yaYlokokDFzqVH6RuNr40BAGc/3xPkG8RRd61n05iAxmdWs8ZVVj+2FNz5yLkpg82e3pkNqDIE
khc9ywW8rex5VTK1SvrUk0i/HmpuUhSf68e60TBKlIF4rzcWI+AUMRZieQpUAdofRdHzPlvVGq8G
Do2eSNlLY+5Wpv/8SXHJ8McaP/xOm1Kn3VvueXQ1dUKxKGpPBAJoUOy3sC64yT/xizERXV542MTN
goQwX3JSmU2x56+OF9w3cppwovkQc6y9KD7mkDBZMcsv68m+OVSj+nPYe72c+ZVXVp+Dbl99Z95I
/ADAR5OflbgLmWOtsdYB/fCrhnOmV9ke6uU4iUbi4dGWXDrCqj1JXq+svQm5bOAvc4ZvHw4NeE4w
uWijpeCHT+e88F189PuT0DJso3qzyduWU909UNKfiJN+fiHGQFDpE2uiv88md92Y9dHTMUHj/Qlo
3TG/DSErBHS/9cwt6E19p254yZenb5LQG5bbvuUM4bSpSb7kGJlsePrS2foa9CuNOF497UWy+k6w
cXi5oEIFMhQvtNH7+z41z2awcSJlRvzQmrL+P9/YlT2VWK4msn4msBddtN+5O0u+lC2Wqukq30OW
94CJUMGJ4pKB7kbHamUxAt4OwIJS5Cf690w5a3lSvLkbDCjyGAD2GduG6dXrQUnxWTp4r1cCJ5eM
3f2lQH5xF29SThrWKeyabqm4yEobeCN6Z7BSJzalM2o3l6oLp/lGm0w3J/xewaG4c1Gt/VR3hSyF
TEYjx6ZmxZ37jYupnFuh4BQg0Ym/ZAoOzsOMbFayMEBBzlzVVJCEEZY4ppR3aX4/lheVldKUT1Ar
qQsC3ULvH/oXRHHTsE/W7TGCpSoojvNhqWKvG21Z+fCPUTICLmKWIUGNbUOvsUt0OTgs1tM7fSBW
eLq5PLt7nqOzB6UoJ8FLUDiSKprnvrOecOx9HceEoZBeeFkRpgT7oAcx1hEsLtrGD1ILOXxz5RsT
DA5a+3iKT4UK/JHBRCOjCvC5Hz4xgH1HfffSzVe/DWO297IwVJa/VEgomloOv9OdMF/2Kg6K2syk
8ZrTeVQm+0XooD0Opp6jJK1vs10XCUHkOXOv8EIl4PsHplOSKDe9PwmaDAY4LL6oEZX2VtRVchlt
E9EKKheBPIAsSxnzVqVAslD59XouUdV1sjhrAafp3QfHwymFxYRvvlDA7yxFcrZ8OP6RH2AiT+tZ
B1gIzLwTOftzgPEGZyJ2fCCA0tAjRVZzPyFraYNwAcs4dwujgIX1nD/t81A+MvJlyJ0vOF8lsvWg
N1V0JkVoHmwspnikAEg/hTkmY+0x4j+cI4+mpPZlnTJmNvDLuXNc+lRTn2Szp+8MGSLO9hMzhloW
1bvdJCyOcVArEruLGoOASuyixA5LMGRUqPwdPFqEvDexMCk5XuWWOhtqVcvq5WY+FcGyODstKfAN
FT/iq+51wZJbSE+EB645MXpBmkJRTEnScbwIC2+x3bIu0vEy7ST/N1IhmzOldpWMOO7RuemEmDrL
tyoMd/rcig23ENjjcxQJ/Gt3BgcNQ5UjYwWJtVTaQbE57qa6MfGjDaBlWkTO2vyR9P/TmdLSvUm1
lsBeBoImal+vknGKkH60G4WS0Jm19OrBPtwuA1qTlBcGZoQC7G9rjbnHboJQZFGxPmfsQcSU8ZZJ
hUD/B6H1/nS653WchXXYkqYNRVwAklRGE5X9ZLk7z10kFf7ZpTS3GFloI9EknAGPo/1+RMRHCR5S
JtgYxvLafH/FcIzhfT0bQbWuRTxWD4Okb8RRJMwxZeUh4YnfD07OcIU7GB1UZbfJmTfu3Pk4d5NS
hrsXZEpRqHPZi1IWBDoxH9SWq8g/e4tb5omzPJ8458T7NTxgcEI99NX1XsjwZygye8iqb9YpoAF8
ozl9dmYPSu6bFl0e4U8NBxys7BJiTWW82t/GbFMLNVj+FotUhejybt1HA5RX7ePbhr7T8DTHzj3L
nGuYHuAWO25abJVmv4GWbxwun+PurOHeGVrlfMN1jdOYAJlujRsqKYNtdud3ZNahggEI8eGt4AXy
bdM9HQATe1IzN20DpuouS9ovA+MqMC13xzyd9uepYCh9+Lof7mozjiilbahAgZfTZsWI7ILtJ+nC
ZqEDn3KtoJezXuamNaKmsFBrvC4ZdB11479m5NTRW7huyEBTrAR1ewLcA+ujSM4pCEuG50U+vbK5
LuD1IyxV3C2UBK1zZ6EUgClvelhe6yq+GvmL83PTIM8flMCvVdn0ysQqnmk7NpSDMWROTHfeY+C2
TEqxwylnt8lGQNE/0s3ewwhgJsDYl2TAMO3sIbdA3BK7e6BKm0zk4LoUqgj/fwO9Rm7xxyBd5GZ0
SGBypMDPlv6EE7L0v/ZoN9FHhY3DqKRTralcxRD8+jkA3g2DRmeo+4Ylxax7GxhseTkKJ4TeRgLn
8wge32tbJEyF5Tug/NR6aB9AaI7izOpCNOCG9cAKJF6cfBN9eiaGdMqZACcwzu3oPd85LD9s91zR
zsYBzD+HABIm2dxdOnyIq0NxkMuZYkfo9MQ/FTe0r6EKKtNfY05bAaq4GeRL2yK9nJxxixPYrxj7
2b11rAlae/RMIGHhJb8WINxVyaWCOVpfPfVbMIOKAI+h/eRdzPf5nmfVtLE9PMgouPTo+R8PqJPn
qpjHxYTtnfuli7Mq0ImqdKI8ctUv5O4T1ZMYwOLn8LTrw3X/2hwBQ14YRnHVUqN6ti8FNrXGUL36
a72PvNjmFqppWJzjmZ/zsxXFeszk2sdn22cH1fN0gK82KQHQVDTHrD8tAsoKY8qaTcpG8ugfd58M
+cgKUuu1G+kxZ5W7b7/bgdoL0ERvrLcdqqFd3QVr/srWRMWXd1ws90PGqYtVZdpQ2Z5TWabNM+aJ
0B+4NPDkvj+v6qWEYot6trQRU2Ngh+fnqXNGlQiZcFRbp0tRgAPIavKE9kZGLIAyWq7HhCzPTUOH
5B1hFVS+WKPOnTa986zXsaprWAY1PIM/YLy3WgHvDh6pZMRLTlwJ6CGWkSIdB+85qab3L77GyMdG
9Jc4l+fm6jxuwuO7UV2ZyNfsqzAy0KpK/aRbjLBi32ZjGT1TXsoKiVmLlal6GzzKaTE3+hW2+3kN
1qCw1Zwf7q7Yaemxjw26sljxcxWnjUUZWPcbBfrLyrB2miVjG/vMzhgNZxbIzZH38VTk2oiJjanO
rNE4WeG6u8qetO8QwcRxZsgBOni/yYO2NVZAvwqiY2KEUMe4uO+FNJeQrGz+Jt40tSVGqcSTrsi3
WWYSGUAmlw5ws1qeFh9C30o9b45iaRpOZKralf+VPM2CUwNsPIZJq4MaxAR9BlRSoM7q+pUIL77X
pRCzS3vawa1dHOLVOWAC4rXhKUbzcQuirEXsFBOTNIkBGQ==
`pragma protect end_protected
