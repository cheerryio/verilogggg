`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53408)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCTcg9EscIq6lRv0lzTzbJat7ShZQ6RTzZ/gDdseVuunnnUY46w7GNolk
nbUaWOx2hoq85Z4lpVoWMlCDDyJnndUlF9UGaQOb+LUQWkjdYQbycRscyzxkE6VoR7A+bKTGrbGS
TLrzYJJUmxoHof6hwbPU/reWb8xawSmBqTJ2HnI3nXxZnjgw8Xhrz5P4d1gz0v9gX7GZ5an/cXbP
ObN29mdDqxi4kA7UamB9dyhojvJ+HC76Xn+D5MvwQznahunVuqu57NxmMoy3wAVJNbanBD1pH1H7
ruV4CVvcMyOywO0oUsP367e79C63ORLEchJmH5SqXJ10MzmBL9Gf1iJsRyUDWRMaqYO8k+36GkCt
dqXuq328Crz6Z1sYvAlO4J/D4x58fAiS6F+/kPoQn/uGjHGDHQqu7/N7DRqUKTRk7afptz41nCWq
cuvwkLdNgcBxRAuNx5tMg4y4/C3gjVGzDrjS2I8hW5NqrsruOF2Lj4rY8Hnm/w+3oXh8Cx90sqWp
xBP1eSPfB7fkDe40dJOadJC9rNP5txnNsJdQk3d+/l+xDD4eRLBOigLz4yR0p70D7wMB2YoY4Ysq
f8xMXT9VM5JrzHFcnWHh49854ltS1L9Hc0JpBKgpwbmaIQi4nlSZHzkvA6LKFtLIgFDBFhiLXvBa
oR/OCCPt5BigoryUm2pWue5+RHTxWHHdnJqIXGZFtZGzck23hzlhA3BsEX3ccf4R4m+k7OqKULSC
nQhiDgElhS9dOMMK+S00y74pnkzzt5TUPjdlVVBRLSt/eTiEAAASa0xDZWUvjx4480SH2GwRr2oF
D5DOmQj7YGGQn/3uhDpZNOWKB6GZwKPPpccavNnC/ZXFP4opzTzW9Ipox9offvkpqDaJWM0Tae+C
IkeUm9PtgWKtT6zTg2U5PQACgiljenj6qRI84R0wRYXsvCYv1oeanr5TtI/bTF/s3erNB+jsUX/P
B+/+Fkqdv5BMPRcvWNpKqBPNf4kEu5x+KCfMjtvPNAvf2D9KCTf+qovvysWj7XXrr6YPd4OO/CcD
j1uwt0EnBystrdIKpy3WUh50HmTZVhzSMBaDb5eYpWJvXjcGxTbxtOtsCEJuQm7q0xwjjiJmeBpQ
Av2NO92gp4cay68SLkfMaTTy5VDliNMWvuVj43yD9tCIuwIu+XQ7Um2/fS54ZOvFE0W38A4QZtF3
h9FzNz37Kt+wqBJFn0oJjuZZFOP1J4VUUkpIMlNflrfjOp9gW48RINVTYXpCzYm2ieNt+qlUCRKY
4qH5zKWr9pOlrASZtVZLX5CSXn4MGAhH6rmeEvXvpNZScATWEVYi2YUfJ1bdcDF58nCiruHbzSLp
aa6HjrYxxVDXUcBKc6uf011JVeZrWZqi+wMxoheIlvaGImUYIT3/YBzm3QcQu/KuetcrYhLnG0C3
LXalnit6fU5m+ahC6izI+qcFit9d4NKRHacZvb9GY6ULIUDIcel+0MLOYKzflcbhPwPJaxq8wMRU
cqcXI8exIFt8R4j7lss1faJ9wfpIRrQ/so/oacDBkNcxPtTMLMd7XcYlI2ERuNKjTdBQRa0CZSUM
6GrDSGmoVllZcfnejUjbN9WV8CbJba0x7q/DIRIg/Naazv5DYO4oJgz5LC+G/TeKOGYkiAdsRTnZ
kZDLeK7wAR8kekwtWFIWx7qG1jlrdUnsoS3LLvekx+MdCZJUkoCDv/T4LS9Uy1Cw+FyTk/wH40Qz
kduBhl1Zbo6RcmqXWhRELUzw+8HWz3YCHcAzEqFs9hkUNlN85/so2ZpqmTYgoJAwg+hJlK5t6rRt
/GuUfsT9pmG+or86W4+jOwfYJ8ql53WUjZcH8PhbcbA3TvqJZafw629dn7MTrm1Mhk4BKho85qn4
yTZ1REOHFSveFrQLbwV+WvUqMuT0dRkpc7/4XwciEjXvzC/XAgdcYlwPpf72qc8BAUkpjKXn1kxp
Ju3dy7D1qE0/c6AyLTKjerw5D3UiBjDrpY92PvttX6CSp5biY9fKdqUyIpsVRYsaToj2JaiCQdjQ
4yRAOVtYGnjl7NRvT2+pXLOOjHeYTOf3uat5X4hgCcEUJ+cctMQAyW6j7PsLbOwsoeeyVn1pPq/F
tDYZGGIRdey2mrJ69jFAYG1/re+hTEpJsygu5QGheTO0WnXzZ8Sa3nbJPsbaBkXYw/Yn0urtr4+c
kaETPQsjLUIBRJZ21SAV+tuSpc/gd6BZMP2oqMrP8owxzP2S6SU0tv40aIeJ0zAghveAQoriiKdp
szI3YpmPQsGEUtr+5ZEJnRawk0sjDABMlWWVUWiGiib7Tu18ZUkuawSZ+qr3hYkm9q8EXDd3I5Uo
J2V9ne8+w2rJ4rrHkyrCbX8FQZQWTGyqUcbs0dAdi3rg1bZmv2Zov1UKHqclWBsHrD8v1YNYXB2D
KPijlDpBjU9MWk1NGsLUJqnL9hRtCT9kBczM7L7kms/jQjm5FkDF8Ydej/oKQpdoNaNnVH1Pcitu
vGLSeiwv76ioXMQqPHWoX4r3lUEMj0qXdp6ytyawRqOQBRup1Gw/wLJTa7bIZbt4o1Fnt2TDZZkC
JC37Gm1zpvMfpOpBqx5vzEQY4F7I2hji87u2+3YXmu8Pu9hf6vnuztfIdTCD/Yaa++3A9MpBoh7l
ZpuGQftjr9V9Rtgzigjox9dlSypeYrH5L5T3NabQEaTk99c3KobAs5CQfmvUTUyHXsg93mgoCGFn
FhWdXbPTasYCFQdLSFBG8WDLfBX1rRxdzQ6SOBUDzRW3XFLPwXyT/dPpWwplX9mn/+IWOOtKFbjM
QiawJUIks7hKIYLMn1q3lAPQWK3GcEkSVgu4qslsB5eFdNn4b3BEZsYK8qPGKB0Zu8Oki5VLUiLu
Z/92CKgdZuLwZxJ2RRVVMxt6g+YCT3t7wWzYDPATgQJ8vY7IcY3Mtl2YsipDaQiHFlp9Hu3nm8Ch
LK80MJvJUoKHB0VbOE4lsYBMrxm1FUa+OSv5PQuHLPz8sTwDKRON8sCi7N/6stE6vRm4KoF36G1x
D5IDDNzMLgImVyOXUk5lo97PodbNN93QUTwqa4qCzXr5K7YDprHar9/CbUxQJEk68apHp9sTKo19
Lhz73wc2RrMAFHOUsyOurYU4rQ+RX9re1Gcr3TiJy31riGfNehnPTuCiKDe5kNQFmp6i7bRx1or1
pzT2m+SGv9//RlTnClIUzzQCmyg2299KkkAgVcdLiXJW4HnfT0ZjdgGYjBIalWKFWVeU4NbqrqzU
covEdt28jOcyGbTYI2cyeym0Af4+0r6A1MzfBSnp2M+xNV5gtnVzJkTmAUMi0VY8HRzb2HkNvnEF
4cXGwzxy+m4fKIkJXfZ3DT/E9UAthLcAJIIdOTDKmV04Sx/bZ8nBuX+aZ+JEbv6hRJoquAa5MVOZ
3HJBs+FpDx+M1APh5g5iGK4GTlttUMxEhnQzmkLmHQ8uvOyyOjMRX/Y4QP61H8wnQK31OZbmeuwN
W5kcaUAYKoEFY7hrXUxZynS7bX9FzTyjmIfUPqWT8fuNQUEdoaD1mPnaieMBwR3K/v6fvYXQf1Oi
Bc50WT6UrlMnguIFuhswLYIZ7qS9JPLGDCLy0OHCPH87wR4bv5Sd1SA5JBpdY1mZz93AYXz+4PO2
shgqlF8TR42R0zdYJBxtIYisrWRVl+cWNfwWXDsqGnUFbt+FoLqefjM2X8221RhQv21Rtcmniqhp
xYyvrDAhGNqsgrLcvzLXlq6ESm4iTskPsjfrUzFF3QWqQ1RWh5JcGVgcdsG2oNk5RPafs5liDrpl
l4/mXHWsI14CP2aCfBf2NwsEguvH3uKCmz0IpoTKaXXRTt9Ie7V5eAl3kwJMpOjbLSFI6nZOmlFu
ClYsuqoLmrIivJrKCBuVYas0fE8VboEfdj/kK4DKnikV5I40yE8Hr8/1+6bx1SMsL1wm+uQKEm2R
GPL0ujOKAVLyY5Ped4ug7ZUkp5luWEYfjwcIYxoy8YIWzq5IKumhT4KbSByKy+qO+Fd8bUMHmTPE
Qoprb5lUs5xxvJGwcLK3hopyQG8FLjfN5s7QoF244EyYojthhXq3WQjrGEk/dk5+KFGLIg3BA+aV
HMDZTMCopKzkNNQO1duyIVk+CgYGG7DJ98/UYmAcO2LkG56t3AuTiahfWNyyDtiqwRMp3y4MEzsc
co5uJdqLDTbF6JzWtJg+BAciy5gdYvhzLqu8LMxM8uQk8XAP7VlNkPGS1Z5aCRqqgl0sTB5romQE
d2GoLAQ8rss9gCr1g3oVpnvRE0B6L6Dtql9ywi8Dx8FRb/Bz/VS6thkbLEU1NDqeWB7MtkdA0S3e
z2/OAr4bTl/JIBKcBJcir6pxlgJOd8Ad+lc8h4P9R6WMJ3Tqt+B8MgGkhxi8Od6p5qcjy2Vwlmij
AOJRhjAi0OhUHPjgdbWO4V5kwUdzpJbdLCgnx8YAA5eEPmpg8oyRVC8enyjLrpYr0x41OdgIB8yU
4HoQASVtJxJylAaJqLyBgHJV3X6vy235H8F/Cb1zM98GAuRO/+L416B5FppJgJ1xvNNWZUSgOEF5
SLi2fLEZwVnPpbRNvg0DdN6cGXmXJH6aFpxqbhrBGN+Nx3nlV/RDybHM/yP+km0FI5GXzK+IIieY
hynJLzV6VFIQzq0n2ZX69gnMMkoFr7QNNWWetRQi4/shNfu2L4elT7+0mk0669uMwlsGT5iYNQ8S
c2TwFf5G0SEv9HJ9bcD6MCniqcYQcgEeXqA0CScGnu+TMTqEm79ty0vlg0gpbnSiXfRlr4+5ryzL
jVv7Vcq+vWnRVOUnCHmGZNUOsdrSvkoOOeMY9jj35XFN1VO8arJb2n4hwpC5uprvCmDnpIctC8+t
H8sWHis93dkj/wSNmMG/Rt4TYC6CaKHdYdEUhV0OGO2720fBZvAxAz0/JO65+vvGMgR45DvIhXXQ
sLdg1tVYs0+f9DWYdWOJpHBTkkENaLRV0gP6K11F+C6KSeU3tw+tlGIMuJi1kFg7m58gBxPgMYSc
E2sFftSsEi/CpaxI4/z+oKeBaVoTLaS5UKM/paXT4jmp+ABdkA15cFm4Guk7CXMuLro627DbiiOS
2qdb6NxhzKM7857vx+HJu3mZWKRNXbZIALEU4J6rxBTyLoh/QGX2xY7MM0O/TNE+8zfSSL5QG5Yh
0OvLJYVobu5wN8oac2WqAkblKJWdfUn7YyYGvXAlEX+veVGj9v9APZUZ15de/gev6RvZ+e2F8qQ2
oNwZ4NgrpFzvU5hpqQE89rElnRK+L3bAofHf8FmHBUPw4+KkYAX3vFZXZgk3QiX/5FHX0eCClr4n
VHj0znKNfC4Qf4CuRN4cHjgiWNnWWt8DdE2aoJraZGF0h1YTZLg0ppK8cGtuVnQXf35IJp0T1mVD
CYcGImlqUWcfoafnnUIc8X9ssujH2ntSEsRBLtrn6SnmE/3ME3+eDxwkFkgckxfdOZ8PnmK9Pqbm
j9x7o/gUGIuJ3ONRTo/SGLlzxWOQS4sDReXdk6M5rBqizlYDngRRHXd3IhVgY5nhivwCOPeND/pm
sN34C1wVAkmWQuCdLqKZEu9FQey2+ir/Ad7fPeFhEivRc1uxFY7QGzJ9P+kjBstVYE2Y7HDZX5O8
Cm2oda8cu8TS6Uv5CeYj09WqqX1zUfCwVOcBcbzhcLVccKYOkXiEyEIWxK+i664grZOlB3xRve7C
U78hd4RyU71WBBIK7mHX4LfM97zxaxpgaHyPybB9Q2oKLeH/qhnHr8IjMFxNcyx50spiMKLemnin
3U/nWfUUdn1sOsum6jAsvrIMVd0BJeCEXFBZISZ/B5o+sy2JOznoSZmN9M8Ngjjmwx/dOXLp/eGD
B4qojbooe6q3kUPGGEQjkUit9EKOfLIC92MUawvGJJigNLqnJ9XtTXJm5srr/PgwhqmigIntP607
MyxI1S1AEy3SzAYEIv5e6EIjlOgsyy1WyO2aWHfTwhWzZhkt3D3MOwy+tLIcL4G5D5r27AJLhLgU
6ZwueLB3ueMgNpTOi6WycTjhH7cWZ1ReYDB4NnZYqRQUqIhQBjCGoYuhHLNGD+ArA3eEcd7UYDua
QCtpqFDWhjVlfdf2aeSLuTyNlwui5lwN+OvRKTfJEfxhvGTsgWBpIdVuM/nFog90B1oXW2pLSWtN
ahrtXkjc0Y8vn3bylzSnL/HfCwhAkcoRTQgg/fqW4dK4KEKSrFI/WyKXEPhipaQR0Wry2iCJEPg3
ZAj+kijUfgpJT+Cx9gYtRhzlw/QMiHmi+DAbzPM+0M3NOZ7PbLIHtAYF+6bXjekhZhVT9OuEFSYB
CGVpZ+aFic8er4BXNf7U2p2KNVJzw6AzjDV8d+Y96Kxw7KazJVcTaImxetOHXaUM8CZQenUeeREe
MzjnUywnlEi3KAKMBBbCRug1SAhjkRAHoGzdebFJMw066nAKwSSM8u/aHPCAmFeFTnvWT2YTpeIg
ANsf3tQi2Zspeuj1xRxpQgHfJOkJPrmObox+uTvYVsiknC/VyoPatdT8F9SIvrNbo2R5HC36sh2a
iO1Ak9nEgBVAS0Xup6mNfEtAwRevmiGi+H/tm335d8JZQm3wILYNps6nG6OZ1O8fCNjgv0GydSmL
f1yus4ANhRw1FOVH9l4C3LAY9al3UHrq+NXV46kNjjsRwjs/9GxQTa1/W7v9ylfd2PSLzaCHZ8y/
GNLcHoCwvOFww0iWfxY5dSdmktsOu65tMWPuRr0pflenk5lV7uoHYEmzPB6wCIL8JGdDlamV/23x
OcLgGTxVdxZW8JNfbg941Iebo4K87p4Abjr5QLbOESlu1TsI6cqpx0Ca3lwTbItRtQuhV9bqwTiS
PvfeIaxI+LCvLAcgDGwOK+d7cQm34z34WJLc3rEQynCqdxMCuzCOsjldeuNidIsJnBVmFKOiCLwq
tdS6E3g1RfkBvPoPHzmJwq0G8OP0UODBxabhuKWrv9kMpHz70DlzSZlwzT6CnkrAll4+eCTS6EHY
h2e+MwXoEMe5QB7QIobs07r73JeF/KDoNVTIjroSZfDq0Tk1qhdFnZG/O9zwLQHELKd/D4h3WvyR
aS5e9WBsxL7lUKArTyNyZNUn7fSyfRXhQAiRhw5BH5zTQ3CTvIV/shHvFJI8qtfwyonIIOlEOlaV
kxf7um8s+q01b67Q+SIMLYYBs+AWp/IGQPN04HK9sOEJQDQwIyZWUyFNvBybSA5EMVib6ouWd1Cn
nJl4xf50eIXwN32GAE+F/Nm06tW5MB3O3kK+PdJwUH3/QclKjD9O34ZzM/lB/GfcfV8RCmN6+ljL
YX3rlRYg5edpD/3GMxA64KGx2mvY9Notq0dGCB+ohole6e1OHwsM9ayuZsgNWWMROP0hrYB+MSA5
TV+gGFeFV6zVJeQLHmGCF5JzCjUNfSYU2shs2auFWJkRtGfLoL9eTViWUit+k2CEDLZvVZP+hInl
/g4mifPlqdym/XDB934KAVO4vWyYNZ6P0f8WSfBPUdXwgCeyzogoQWVlUydCY3tnFk5swhRr0HwD
qrPOsgr8CX6UTULhsfpFCK8q4qTj5dolggkRppf/emp2q7JckryoJsVhDoEo75738dckRt+QzQZq
5clKlefRYggleUH16vpqdfD+Dy+sgIbQtDdcwuKx2ral7rfxCFKRmmZKXAznWzRMZHSxWJU82Y9z
cHvJdi+6bG1LcVocWGndSX0NDd1y6DpXdDU+WlFUbxgNkHGji1x8B9/KxyEXFESChSWR45vgQvEP
A/O0Vl8M3M6JxdZiJnuX2wh/qFW8CXmq+H0LPpxwjMbVPegnp20gR0lN+/+F8tAIug9c5O8gKLin
H+3BZ2g/8idvWHrMu0TFSqQ/Ues3hDX3vIvSc2TudBU0IeMXhbF7WYjWtqDxPr3oYSTtUf6oXvbz
0QfNSDtMZxVF7jnnMIXNKtKUnvb1cxTa1t64ysZhR6Ps10OkqocK+VeXnmb5Lfr1FBVOVZwLkBCn
zgyL6V9XCP+LuQ2BQVeq/cAMLp/iWsrFs5BiknS/i0KAfOVZTitk3MFTcylRGydRnKRGmuem3qWz
j19UTFbagoBDrSyi20SPncHP/ik08QsGVZ/Cbj+j4c+481PASah6knmItzHkIWe0kSxUHZrCghQ0
yR//GNysx3sv2LlSdlROMgyYbd7p4itKtrLGvM8Zv+VN7HlZ0+7c/qz3TbbLhXytPQvMYNIliJl6
5ooMajtimao7PwEDjblOWWegDXktrMqd/cYAUXUqcMtU+HfB4D13ebiulAtlGHP2W/C/CHpQlyWR
UBCNBDHRenJbdN02j0/1ZKLKmZ9kLRBKEMLNpeOOXvN2LJxB2mKDdBhMesy1paAPmeWcC2KaJ+WO
B/4qrYY8aLCMiiJum2hR+8Jjb5iSBcg2xpggCC0cyA3UBBD7yOgKYxBnCo4ObjcGwqscFG8Z7sFP
83vVCuQ970YiCwfbHcXrvI7n2EP1nFHd0HLJVTManVNeUwVQudPBWVWLx+xcKirlDjsxWHgExVYi
Gc/Yy68Dsgvp4pEKOIrGqYbccr5p6EH540n1k4gRlc8I5oweJpIfkdOYzBKmuKV3HXXXSNeBvIxu
LXv3N9TNtX6jPTkkJKDMXnayZ407xFE+DMOrStzRLwk9zDGKO4hAtywevpiEJT1C3dCiLRCkND+a
sIHRlaqZN1EAWnvG+LZQtYS+r2bBDV3OkjSXzPih9AGkDW/B5Faw5vrp9SY/DP7rx23Cmt3mqwWl
nKlJbDul0QFSBRfNaXyZAbBngqkDdb88V6IEGQIzjaZjueEAp7tzbxfMv2nntTVCSZ9m7a+ImgEY
I6WpVBp3PhzWLVJu7zXRCqwwbfX127P19lJuvr5bvggggs8jfJ+wCMesmYj0dTLIIhtPP0M97BYg
jXMeK5IhFQM09Aj0yCcfMDXjJqOvBRfFknLqsFe+EWzzrCD7QLg8+VTBsCsgrw8MJfdv69I4+cr5
S7BoCxY5fRrYQbezwFF/YyeVhRV07NEOvhniHvrPwJG/YTn8h3xuXEAjHKu6xvIm6e+ygUvSeDzs
dCxdwjGLkevSeYaL8I1AEtvLjNAJ5fwVdXjB1FlKcltKGrKZSIwfLjXDTYlrR9pvg7/29EmmESoR
Vsy4rdUCuObV3USqxzu+XVP6IQQzSv747LTK7fP9Gf1XiWJo7zCNVWLWCcZ5intBE1SbNMrXXcdI
dDLnjNl+mM5vplmhA/QBCk7jIrI54uX8crB63zquHCqfhBUpF/O6EgOZimkpx5cMUUakQFirOv0b
ZK39j/k3Qcttv+NYwebcs+QDlAc1PcY9OkqslBmq1/bTSyA10p0vryK/UdHcmGtXma5jPEfeusIX
3/xQwh8NK8KeDsJVfO2jB8nSSRI9j5uiPWgJ8slycL0tfU1SAqAheKWkORjE3vYhPMQMP6Cbk0nC
9yOw9etnIRvcD7/aDFj5swmi0XSWyiOnj/4hNdF3Yo0fJRToTRffPbTqLupMQz8SYv+/rxG2G4jZ
cIp3F/cez4VwLvl1nJC93KCmLqqzm9yUiEJCPw5Wc3mBlb5nXn+UWek1FxxGbwUpfw3dnQgs6Ftl
mNBh3BkR8ynxbet4QCPEXzFAR3ODdxIb/IaGjmuDNv+OLgCeAHJF5tyvJ2c68GpYrMM4U+sD9DMt
0XSWei2qgeFkoafSLHxU18qT3+43atUkTqeoj22uuPH4FCTbLsIUxZZ55BXvrS3z08TyzQ54krXJ
gAvMSM7aIvMWSJ4IrOyhM9lER5fyydqohFiyUoYgx2zxs/WgHiMsdc4PNY3V42HFNPWFwyr2TBu6
AKVoatkqU9ejl7ThSWx48dRsqtwle7AdcckRUhoQ1CIl6e2bAk9p5dQndfHSVwzqYnQySgiBZOfT
S3tYYssnUm1F1KntQBaJnWO6t459/Y/SB3SoxuzC3lEJroUwp5kczyCa6TIb14PbGfPVXJlxtWGx
P7cZLy0z09kaYFp8u53yjoDXYrCvAnHfMVzjC0f5sUf0E36fJUJknLTfADLT33j/2z1N2aZAT8Mn
DHlN6+H0AcXPfy5ajNDf03qJNRVgPySWXRp47mfSn825QBp5RTW3TF1hGnacX/csWMyNwHHMkbxR
4qdPHF15HIQ9eQKi+GI4cIR0OYDb5ZM7mt2vwNFuS69r9SfaR3/DPoocPp+nTM4qc6MLLPnwje7l
5oiVKfchjV+wh2uIUn0pru1KihpXIpC/SBnBZ4ubEW8lQ0qds5N8/JLU7LDkmD3+9bk7HJbRSDOs
bEs7GuLQhhjnk/XYM6tTTuXMEgeBrCLnDcJHvRFxhT4EPTxlyKJIEVo3GlQZd9OGbsTzhBsu7rjh
CdtFyT0q8HoEXpR/R17WkSiGxXYlI6MEBCnSFaG/7kGc3dSzumO3RsvQOYg9pEYuQq1vlr2bPUCB
VNofLCsGP8COuh+XXz5WN1a1JuipgS4A3DWgpesjINZyAUuyl6mlrTbAIWXmwNt5H/x/uZaNQiMd
joBrTUlkAozD343ZV8NDWias+AJNTEQpQGlSIdRwwdx/scL/lvIj84oQsn82mDVW7Ux2/DT8b5yM
57djP5m+WUrkItSJLHrYea8iUT4ZrIoLwOlRvyEaR1ceZH4s3qrFQ0gaY4m/CSQjftvhnQRNE+zt
D1IqgRDeIVSzkIfKg+THPqzfSCIMDLONDDE9OvgfefCTHO0tsMSJWOqwDt+mQ4/RnHex09Bv/fXq
9XY2IdFQ402UyaQE/3VIM0MEjdeo1NajY+nCH1blS6HodN3yYEfYNBLq2EW+YTTS+ojrWxYWVq65
jec+jai4Z09U+R9lKW8nAW/0Tw4OS81BzH4rbHzSWxsx86DCr6bkxP1RIrgqp+euwaOC06t98ovY
Me/gp5vGHasEP5aPLmiPcGUlhM+ZC8/ZhiYxYtpVts8j/9LSQyQMttk+iovv1UYXOUC+MLTXf24t
aL6kDG0/XbUd4lxtVG1944zwMWKYY6g3mxYe1OSoWMKWjULD22wA9PjFHXpmeyjbv3TXDx9EsNpy
Rf7zD7i5Hc7WoA1l+x3MazzxhaYdMTToMvTVQy7riBHpzJ/cU9hneXkW2VSFOvBv92FAFPE4Sp9g
FP87FKpQy2hDlleKnZcDuzXSySbkkrfA62aOC6TwkmK69Y2dNPHa5OyiplTWp+NPCTGxD09Z5QLX
q8s3dwUPdeFjIHhbTwy08iLxFK0x42dl+oTbmk/SxJDI3BKoavtB0V17c5Yhyrv2Z6c2jlTr1+fK
M/XQiGxnG0AnzPu8RGy+oWNZXdPrEGeI5OxmCC7IwP6HWWBHvx5NCP22ozedfx2NSJnL2lckpyZM
qfnstP7lQxIpEfJoYmigrCu6N9afpSbvDodsOut0K9Lpj+nVQpuGIRs6Mmfus2J0Yh59NBoCCesL
vSbkP5N4tWk0lf2e9H7bQgzrJfHZoKbcQWZ/9N52BIttmc/dDX3q1GAYhxeUB7+xRTdw2xOJi9Qo
lpu8c3AR3W+vAtxq6Uwq37OCvY5xjWaNzT0rmyi94UHSk1OLizukgTNuJyJdXGJcThM+F2z6hGOu
5KiIhJ3OmYjB5oDphxopfEfb3C6jB5qmzZOg58woGzgYnwp05jGgoDLZdAKkw+5M4rM4dOfm2930
tGum5u1hljT0zzjwGtC4FGvQibK/43duHJfnavrUcKTVAnr3Z3qxTuP6G9yQgnUqVdU9L0wyRxWQ
jIbLW3weaNVNfTCaOlp7Bp7IKfMcDeJ3qYd9cIkO7roBPFgl5HaKMDSTrKWJbryggwoCaXar3y4D
N3mf+SaVkaYlS6UohXs1qldR/hsFadv8JkWAyDCCzdAFzxVb/Nvo1NQcLJ9RF/6uNiiQVlH1M+Wo
yuu7KW/KFnC6id4WwiuIqxMvryncXNhkGlonO2hF4bQOkMNflLVH85dnfzX2bv9Sg4ptOw3OlGhg
YtQdcVJz4QAm0q8kuZbcBjR+LzTwKYDXRCyJCbK5QJ9okUEpbQUCe8mX2JCAKaADlTE+ntHyZSJD
NQeumrUElAm5V43CIY76EUdgOnuq2GZm9pzyNvjEY84v07y6446Zl32/yVVDk13Hpo89iO5PRJx6
m64x9AAhQtwJmNoJXIAniw9tpPnAoOPngQtiO2oFpBpuHu7M0oWmW7kSgouWgt/O89HfTiXenvhk
mExxOCST4ha0ezWQhhcbUtGTtX7MxmyzJch7TosRT4VbXPcTX/twj47DuZH8VsvOgk9JO4UVDKeq
nijRJ3/4vMWI0MSeIdS2T0ml74G5Q9jXncENVT5AMCkJCks3UdPRE/tC5keOS8N1xt/HaT/uggaQ
bS01olgOHqmG+Tsh1xv+uGzkKBJJbPVBKz2YMz3Gme/pQqmUssdccbxNfr/sn1tlvEltBtpUNtS1
F1TC60dgT+msxxyVd3Nz0GTmSHfutpcprtiMBHfTBjFuVCcJ6jzBE6Sh0uApFqKS9/EYVWqkucju
otxoNGnBY3POKUhedtKMkCakDjnKae2m7uvRLidAV4q46H23MV1fSftnLMHY+gmrgEx7TOtsGQJv
YpxliZ0BK/4dYVsqDExpP+FAOxkLIc7eXBH4+25AhgPX8IchQgjo96XOV0dHufvFLMn5RcbjeoPa
g4Vwa8gBFXLLv4yv1dq2P2DlmbOxTbJV8OLRYA+stumb+7f5ibVZD9SJMMwHeawS3HQ00glikNjw
i0CelwK3pvSRolzPoPOkOA4qwcCjkbWdCxBOPg09xBmAg8bLqU7Im1FSgKwl3F6ZiTr9eCiqU/Oj
NOw6qDQcR48vp/JIBI2vu7EhjKpRXibw+AhHOVTiG2EhrgtPHHdHUQ31ZiIUjcSMzpgvRZrRZijL
UcgC1Nmf9ycFdFMBfKC/g/1JWTxiJ0vFkS2JJhG1sCNjlAr0cOdjWIFNyJXeoymnAGTMsv41pdxQ
R7hpzdbqaP2BVPlpL9kle3CGex62rBtrdYXbDKmfoaCJo6KwVR95r8hK/BfavNFgeyfMjkmSDpbl
QgB71Lxcosu+IQ9ZM02J6x7Z4/qUe04JeLpqucvXmDk1zSpsB4tD/BXydQKN+d4hXq/F3xblJvng
FwZh7dXGZ7Sn+HE/HQZ8CP5kvnVngmQKPthnDfz7uIGc/glPeamEnw0ZlbhmoutYctynVNRSeL4Y
Ep1tOYn5VaE0qdUyzuYBaZEWXfoV9VaKTsTEQf6gLThgP2AS/VzXVoqwHynZWUHjl3j0Lafmzgt8
S/V/nnHcvuHjHGqB3qPWAQsh0jazI66wTQFpMGRno/48QHKgVuuX1wSbkiu4ffYAq3/hiddIPEz9
TktFcsTeXsMjBUOJ2KbgyR9aDLMc8qySLF5sOXASRCkHM0KdKCYXugAffY/Vjgd9Abet557YfOr8
Ro7wijYHdVWDvrFq9sULtLxTxBb7DurDcxj3MoKurEH6dnXAYU/gyrPsLfIyTGYQOq/xFS4HLDyX
yCjBVASoC4h76q5lkXzD8OSKQcJhPzKia1jpDklsv8YkaCaiUGi8FdzFGCnpqp2moKTveEvsABrr
HNA/5mVh+ka0VreyEhGV/VjFvxdWwjWBTFwc3JGvOcYjdsVTy5hV17stB1LG1RtDyZvVjOgmRQiP
l4s/8kA1An1WxuhlhQblXwwh32z82jaj0uthEFHIO+lFvM8IiB39jYG2DaeYP5PuNXSQLBERiv5c
efAZDQ6pWLK5xeGLFm3QpKnirUdE3dg/6mBxSREmk+/6UtAgmYgn3sje+gTvChpeu868JkMD3dIv
9rOW5NO1U1C7qsPKpUVMoYDKqW/Kuqyk2U4cctSFxNY9MDrgR5qpXTiyuWJNfYd1KGX/7Nf2xL7/
QnNX6SCwzfGsguxEHNxWmMXmnyoTmznB2YLjWNYXgK0XP6SUXBlbpOKvA2v73B0Tyzx1ZBogJMn3
6pqmzAsIDd0vcJAG6gHgu8PETqztV5Tzdk/QIqsfMyX5oCWU/rQ1MCdraoolFZjGzhd+SZxfNbha
GdDHEsxOhkW06/8PZfnuJUipmCgz5Cuug7wsGvfjI4MyiWkYYXYBDztLXeu92RGhZlaiTdk2V4lQ
OhwYN/Z2fPBGjq0k3EcFaSP/OQ2tyfUWH62p/bSji0OVuEeDR91H2jU+zUXBWuyhsbP7jvw2UsgG
wYl/n7kjO1uRy/wFpP8WMwRRL39QWJB+hwxkBthlhGkKZ195DBYtMJVDRf9hY87aURzrF5kYm4z9
540roNmnWvNkq6sg5weecBUr60Ux3U5HaNiLlbVG5AIaSFvyUl2RcqXk24fgxeLpPiLUtXRhXozV
9vUz4FvMa4YygSxXaCKbYhqm6soxUMzT31+m9+iOq/TnXN3vgv9LIsr6ECp5pxnmcLAGuEmUEWGd
oAFFYdYEM5c8wM6joUNpB4KYv2cv+CebvkN4X4Kjiq67Aly0vPdS9X/1j0FrwMKFytj/jQcfQmbE
il/+aCvT9SHcrmviB1239iN4G8Jffn178YHDOea7PiMlTyoSr4919UBX//HYA4KK74+LLBHAJJUY
/xKGjG1rBYY8GR550ggkLg7cqTPBk9ny/X6Nua1YK/adBH52oH3dy5O2THRva1mqJWdno+cbdUJ1
HUeqz5Ai6wEcEGq3CcbIiB3kUIUjp9kk78OjsWy88djZ4UVp5ZJFJw9Z4fpyV81OcRGrkuHEGjip
gR7nGaK1D/RZS0DwYg0Pp23PZKAcyoC/vB92uvo7DOkfuJ6AVGcgTZnLvYTpLdZkUbAh1CvIWLkS
FGBbVeudtmTWWbQ7cyzrjSotJ6wbWgdDn0VV7sJMJ/BCgnSUoPJ3XLUd9SPfUi8CBOKbweIjOUfE
f8gdhAsEQVvkohrjMU5gEmiAQ2gsBDPWLqkx077Y9SvNZpMHNf1vgpSHwt0qgyxxr8sfUC48YHD5
EH7Nl6Y8t36XA0BaHkFveGzshqY2BJvg95oI7SSjglnLjFKxTNTOC1ZCBVi7rzIn+IuofUfqU6oE
aGuZ1P0qaJ4XE7z5urrxGdiAZbPsrf/SEk96bMXmjVyk0mvL6gDXAF+0DCi9VmLAtEKXZZ8t+zWR
NlDYCOvowXtdR6m/uLiYcSKbl1LQZbcBJcnpUwn7X315rpQhvUUOj/s/4N7SLNIbRJPcf48hcWK9
vfU/jv+6jJjJPpZyMEqbZ9ti3PHfgGQxOVDe4XJoA6FOcXviVOLQCFUta4lhWMqBmGxv3xHlLMvo
MWRPJO3rDirGcD8Pa7d5KZ1VPvrVB1F55s+9H2UVWnaiRVXGI5ggEjUbHyP3sTIcB2wK/hUFNQl+
RLasrbTA+9AmGIEODsyXW+twxRd6Y6NHot4yarljuarQMJXsJFn08mG7WDjhLalNR3NDDhcEc+FC
9HSmLpIgFd3F6k5TNrPeiIRnoVC34Lm815IogdHridz9MXzI6IYR61VA/nTMbXZaq9X6BsV8Hg2h
WO87OekJhjs3ULxTgnT7u0jPUOGGUqe/2hFAHWAunRbkIYJj4dOylQTGqPG9biUhVQBfiZPOfuIq
A6z0b5QLidd48f1gbroqrs8/MJK/rjsswS5Ok9hF2KMgkd/jW/GWkHxzuB4pXrcRMfBqYFjCIFC/
pjwcW4MQlkr04IPjmMnVZU8rHy9/2eDc98v+hN6jLKJxi+MQ87geukxc8mbCs8x7QKP5rEWJ0PfU
Iu1ssaRBC896M3ZAy1T7WaiDfgb+3IvtXTqZWzSChxpQKKSXDJBunCIEQtlvGwdpRZRCyTVl+lPD
gThkNaOaWdHM8FEtm56ANLHgVAvnw06WOy3A6XoryAzcUgFVmJja+uLLTJ/VQh93cGaFVgIEGy1+
1WjlplKMnZp6C/I0SKGp/zxpPfwRfZ8DyLk62HRX6SadgYgQXCcZwNJ4kNaAxR4iVbRdTqjEkQ4P
5S3mSXmenNXgDKfq2KcEwri8L+3OTduZblwaaoFDVEmphnTKv9BCWWBZGPcMn/LHhW3jycSgyTrI
8OC5peyZ+2EeeI1nbvaCt2qhFeRtwz/ukgVtFk1O0l3aWpKPw+l48/PqrYHf52Ia+IIHyxZWMHj/
+8rHiikXm6Z0zFj+RgmmdhmVMOLxWTqgZea+grDBBWzPWSbdYK73Fk7xm5USATiEBlkfTqgNjOv1
8agsDLBb6zB2WfqYkaji9qkJdhSxfY9PosjbMw4aVUti9CkcbLYAKn4GRtRA/6qn+urTtAvL8wjB
XcHr7Fw7T0xmBPZ7wWDTai/bRNRvZOjnXlgAanWIBQTLZcvYu6rpWefzARtS2klKH8EcRAojTFFk
d8FHLG2nMOUP8GEzXI4eXmlNql3bLnTzJwGgzVV/Joqwpp1zEW68IuUyVUmgcADeW6R3PfJ4LCmT
X4YF1BWBMHFwb5d1ZE+DhVp+DHEtVwxZcRBtu0CEE99rpq5zmc5i8K31SWw1wGsEUJ/gGUlqYA6U
XKuYAxbKCsHVPY8T4F1iyvkDi5srSzUuL8mCoPsBeRu3J/9G8d1fBpUQJbEx2zCvt4mzTzA5ichz
sAlFyFRjrrtgCFbWToLJeyu1tLNDHZyyASLn3pwAwql3jjuvlrYX1XQdEeQQVJLmDaTXhXItA/f9
OOm7aHLGuNfuBqLOUTBglxPSeijDgjXDolEJIu49p52GWpXcXpW7hUD/8BsCP0OdjksF/jPYW7wA
AiQ4kP0dPqICT6eG6zIw+3VP5LCqjx2awyao//6wwJhPoBQbaiHzwfvvX5IhsyNXqdLxm1+Ff7z3
kmjCwsP9032MNMqWvnJVQRZS2mIvG7P9OZqVGFJ5JjqGeWXJWNft1+HsAruMDl+nrEGCC2iJTr2V
SwdGRtf+LLW8RlG3hvJnVjnLaX2Tw1TY90Jl4wiPh21DUkAuavoh29u0LKJRS+nLeHowmuFZNs4m
tptXIpMyTok4+RUskkAgf2TlzWimn1YQIvDks9y4tIj704EKaqih8pklnpVIJCEHk0zSCqQxWeDe
/chzCdQSgE3Le96vgpsx//sV5HCE+CLPd0dI8YAoj21Rmc7Qkiu+wSsWgj6tcc6Ob1ytKO05iHul
hVH/K+ooAsiNxOiT+6nDsuylTCpADlXyQr5fCwedyc1PeU9ST5CAQhazl6Smf8DkpWsf1sdlHCBV
YivJCDxsPywiwOx8H4BLliyWL/yNzgurZ/62vRlAEdk1xYdQcl/Wj3DqBwQQ6unEr+/3Aix6xMV6
X/Dl0Nlrstt1JJNNYXxGD0qSgMbk3hCOu5LyILI2r8Qqr/06AWpcTtDXiStQRtM625cQIOsKvwjQ
8v16Jw/h+52IBJeZXh5p2ozYUIge4vc6sbuO4w45gX9sVunRokAoMJYg4ij9zZQySLVkCxTZe29n
JZ/AS0DEFZGUnOhptSrbo6jx6IKYQoIh2BUz2Vg1CF9hfBozHjkw4C8rHvHG/2kAtAACpHwB1c0k
11JZsbEusWpv3gdInGnWgDmfSnYCBE7N620jpH2SI7MtNwYsqI144jvfh77Qv9ivkQuelzbSPdJH
1ZvNyWt43JQvilTBD93erq+x/xliubXPkQP6Gyv+n9V13TnzW7gpio+Fpr4i3WDXKUuEGVP2vDdi
JZfOMgTfPsuZRisWH6FUsEB8sfL22Xdv1cXs3uBss6mA6Vc46QSE/YxHGIr2NapMBAOjx8jHuYi+
mubObhIgYirq8lTfpxr3HfT15iWqQeRj6KjtAekMVJqdlu3gwDgXWQPkvjc1hUo1v9vJXfgJjfYW
k6ZAGhhbdXtlKDABgXrwo/+7+UH6Qh6PGddkLn9ptj47+tB6CaECpMSqaKgUfq/4YEMbpc3HdE1f
YuI8UjRFcpT8UXAPDyVWeILLfWnohOrkb6jaRiKXdRiWG59fgDUdj5DH12v/qczrLn4WFg+yGDzl
O7Wqnfei/i+tFZ/56+fsSqzEmryERH7tWybaTDQ9fDO4XKp6w6G2cHvIuCkMguYbMCdymH/XpbTr
+mK3A2Rj3DtwvIgmpkNDP0zXXqidxyYLa1Mk8XncVjgaNNZ3T1DNvD/RYYc831BRISL5voSXiRbb
hCMBkQJH7WIQ08iO9e5F5sVK/WTsWzAgHUd7f16oPHCAENAlCz8Tq+XGa1b4BPqFHW0odotNq1oM
vc2pbt2GgCdvWSZR/Qfnl/HHft5Aj7AEgw1qmyAQV1bpl/h977nvZdM0emblJhlWYdKOvGA+RWQr
6cNM+To1uumIEpnDtSgoUS5WoWDkKlIdLdsZtp9Fv8vPAPzcgt/raJN3cuR9IVMhfHDH7dRtghL7
CQAXv++umi15Lo92R2Q1e68Rnzd62WVceuI7ieZYUa3SXx65LKkAGhCSarObEr/KQ74UweOVdqzD
X1ZBK7PoJgkScAaX4lfKItsq//n++uC8zR4DLZ8wLwZF5tuZTfkzdgTnMIW/0axHQ2B55pm6Qfh/
qxSUAqK69E3Put1gd6dTXIxzKlhSlC4FTq+bdU7A0rsAtMJn0NUg4DWTxz6VAJA+XEymOz/sXRD1
cO4eiWpWNWjCF8816cAWuEIfA0ZZM/n5PDpCLCaRt1Vj3sy7KSJYuZKBs+/1c0w+Ez3AovMNLbzg
JeUaG0g80aOBwk/qvnSrXkNS0m4lVfuxsK2FSZTEcMuA5sqKxdYNJMESeMZWdkFwOc9nkABc0M+o
A8K/DIDsFWoSvCJwyQoDpDfRmL6NO52E3jEBHp+boaNgWMb3ZC1/0yoYo9hGnNCYuYHoF7zKRkLa
ppwuZ50h6JqA7znJ4u/yNCMQxVMsTLJ3xKOV4nlsiDGGppBsK3xdXpqEiAauQ6DkM/DalxWGkHFf
FoydSGL2zUclBYGjMaKcLfmYOcSDC2/5Er9/ZwFYr563blqqqE9lbF2ghzcLglavyJh5oey+7NJ2
EtsxK33zqPatTq/jr5wu99vN9V+SLna3yIPkhQHSROhD7RoIiMHdP/LK+BH7mPGPx283VnfukPa/
ebOCX0wLPo8xasPMotFqXk+4cirLqDvu1UdG8Vp9ef4mBfTmH1oNuPJDrcIWLxZ/sfbJT4qIMlNv
leIfKPHDnE+OHTR28lRXNiLwN3nazAQ3xr8qqjSpnHIoKAGN9CzN4Ii7ZXAt1CJ9gCGqXJxKMAPN
kuHETKy3rmz1VKYO2l4Dp+6aL7kRNVNq0hOeDytq3r+Cfs3SiPuMvtJkc0qkb+MDMQ5A92iGiXyd
xWRunegC1Oqm2b0cK7H6EOBl8qq9A6V+gQ6J+aqKF9RoiQYnzIvafN3vu0b9h7On24KvZbHGEsZl
5nM0aeRv2U0kAZ4BHMHqn7hJzGco41HlZGCWtXgDwG0pV9w5/Mf/Ve3zja8881THimyDwRbmpIzd
PX92PBOP1icRhLX8fNKTLTdeHMMm4vIuefmrlOBamzUyaEIoFBqQNC3dd/kOIuf63TjxfQZiBkD2
KedZKVTsmt8g9eS1Xyc+q+dwVv6sov7t+rDKQup1kbbs3sLi4v24+iSRVbImrDpm48vgQp95luTc
Pn//cE3SY4SIkDT2noj+VsKzAEio3lblsoMGFnMbVeKCElwUNisafYDRiL/Cl4g6kWqxzD5x2Eoi
mpGdgZE3GhtRYqxYHy3Dj6Y1MW1VIh3EoSFoxGCW3h9ziOi7gJmrkeoOuby6BdKtY5lc4E+lSXR0
t30k2UvUBwuh3hpTskmHBBRFh2HB2ZQbW/FOe1ZYJivJtXpwRCNMG4vw397vYxNs6CSOvwNqC4CR
+90Fz69dIbreXMbRgDmjmB1f7Dka5cb3dENCpLOxEYnuQhEMC6ODM2MNi1UMUE+lKWBkKx1nSnXP
eab+2bitCYltQTBZQcEWbVttBhEjFBQiWxZMdlhEFr0VXQmhb5aVWUNdBHTe8a6QCI9zYL4/4TmB
y9kK2JJlNaaF6hvl+NgpRyioGuYsz8NrTw1Q6wT4W9VRnQP8ABMTGUC64CTZqoDna2vVZZMrTFYU
rPp9xcE155ebdgCaVAcsii3F1tsvuxc54W/liaZEab3p3KpDxuUFsLtPxZwqPeSdylBOHwIhpP9Q
wZVnsDvE9u5w1OIvOqydYo0V0h6/Vz4xNQTh0UE3mKg9VQwBSCujLP5WckwHX+Bw3GbuHP9iLpcc
ZNknlWWYqJg36sFwtgCSa2DyGe4wLvXMC3TwHAXypJ/luNxqJhQn4V5muu98wuQt2KxmBkq5cOwM
W82nSL0KAgEQzKu4c/oX+M/xoAVZ7i7B0RtxjSocGeUWC5QO5Bc9eeDafOnSiaXrcZ87M9LqFIrl
kuXmzWJkWEh8ujVwqe/eq0026OSqCLrNIcJQHLBWy94Lkr9/AboXBNoryr8ru7uFrefRpQ/zbKd5
rmdkbz8b5OLv3GCAdXW1GJ4rR60JZMzrI7OUOyz/EwXUXabZ/1nTVXLW/ZiLdua9Cn6UmaoZ/5GS
SLx2syzAhN2pF3GX3QvXC9LuZDoGu/FYi2+ELK1ib/d5gp22fBfuZJM6xpHwFjzTR+Lb5+cI5kiX
QXfwt5q77rL8Mu/xONFTWnuii1bnl0QumnalJW1uOH6u8WfNmrIEM4IZrc1gDfqWwAtrGHInjYcJ
gNIU5aijqS2zvG8XPgmsKwPQeQp6ZnXE63Q5vCEm0BW6lIoYyORXFVxM5CQdIRoyZxZ4r8Z9OOCj
6PvolEWH+F8W4SkifWABcTtpnkHdPInynww28/mW3XKR2o3s0laCSpASMbh+NnDylzLE4tNBROeP
6JY2V7k/32+ejGro/+K5Y7Ia3+Ch/PXwNXCswSSxf9PkR6UnNiw+E1CiaxMs0aNH7ASg/w9WPGrQ
+aqerc1D63PijSZW+5tgytP03Jk8jmR86decIb5ZqbzblvSZfyXmYr+saZTquL6Ow1xrNWSInGys
cV4HCOggnJtPjyH8fTz7x3TVdeVXhOvA7J+Hwh3IZ5HWkbx6i76veDgCbD1ssxwSgXjB2cOrvE2r
+rVTcmGW5ibmXcia3LSHk6DmoTpcIpVLKAe9nYHdgwBD6VRvQ9dSEt9TdL/1dnZsYQWfxdbNwWfs
TPW3N2ca02sJ5C9xUJBrbFDbij+YH5nB3ibOhyV9srnVpajv9RK3Dqf90stWcwh1BH5sRnMeEnhg
ZuHNQfMl4POT5ChJ+TB1Rh/yX6iMJut+HxkjE3PRBUR3T2wEKkljznnasp2rTKz2Az2TI4ZcxGA2
fPiqoYsINzzoG2YqbZ0g5J11yVh3a6xzfYADGkGg0DTUI9GZsNQWSyns569A21vuKijN7ubqpg65
wWweZEAPumbtLeNlmakti2OUO2g3KZ3lYJSSxCB19npttp4O4zUTaMCKcrEPd+te32cPbtl4YcZA
rYbMtqqPnRpTbJPECtW99bjQDDPpCFuLQF/22eDmZm9pgmnRYPMNWAsCZG6kJXsr3zhN1w5GTzm/
R0Wv1omFP4SM8unOg8O34gmNQxGaeEPRULDxYZIyL0T0sXcvMEP4w+Z5w6I/OcYn7VB0GhpvCZkh
JQX/139z1qOcNdc96mXSA7fuH2Y2gReYLutH6WI4Jn7jENeDaTTDuGs+SzamHLEowtrj5OiRye9x
4aho9rMga8xXAhUzs53Xzerk1N2EClZGU9Y0hlQDCVDJcTX01okNoMyrREGqC++3GE7uhBjwfsH5
puBuSiFJoO3KgHPTlEDBRsgy66rC9IxDrmbY7PNSL88/eI28VKrYBQ4gEXyn03Z9zjt6G7/lqFXR
nKbQKFFYvwEWRb/SoPUhHuSlyp7TlJ5W1dRECy3O2uyX3lq/CTIgRYoQnLsOsnIZryI/B7Wm5WbR
t0VnmHJiUpyG6jWlwxsJnfWS0h87U2rJ2xvGW6atYhRz9mZGiBo7vYSUWY0t5E2g9Ltb12kRPC9y
eNmwaIrRrtkdmv6+2dhqnqQbJKSNeuG0c+LNenUYMDroZx/QpYpZX8HG8j/v0wG0JE4fBc6wXoNE
XDsDnOru3xbFd9oufPbe8O8iWros8mJiPIvHuLYc/QUZhmYa7KwFQqbOOt5vAd5h/mbjRgtqIpGH
+S4CDgxg0lyLhOUJtdiLplqpNWoqTrj63hoxp4p15o/K+CzvHF+ANMwUQEPmoQtFPH6M9ePISVAY
U5G5R4ywIbasFkOVz3gTzI7GdrZ4XJEgrd0bwmueB70CWWZxX/3Uh33RYFVz3PH+Dz44cot81nM1
FrQWkYZfi4vHcoIHlrWbRTBpfvhSj5+Ny9F4SYLprGdAHLpWGKDd6jVHE+j5zsS5etbeYSayEndQ
x5zm7KEx/+vY9Sra9fAIFOn5n3G1Xl8Zzmoq4UpjPunq+FDPU6Lp9DeuOmsUcyQ17Lc/tQJnEPI8
xVh874spRvkE3h4Ndr16zdpLK4YKkGHZHbFk10eUbGb5FTsuI/DhlAjplxkYX5eTGXfsJjqHa6y2
WqwwE6xnctZ2hDQS6ljAcUSEpsp0J+CvkvZJ6RpXPSgXnLj36+89cLOvaAPJV9nWGUHbVatzBGr+
+o+XnwJmx+9WkNgC8SQAa7ZzIFoFKBIl9xJoRoLqsa1UsklQ0QWcLdtCM9g22iN1Shl7Xpq4+x1l
cM03U/BzVTC25LRpvLScvOnYyTTsq8skUFIPB5Ttzb0MLqXIdkqJ1y7itSozaBHeQ96Kf3SIqjh1
pXLG+xtSVFB3hWg4iMnkNf0nuhkAK1qzllLXMteZN+sYEkAsYz/yuy6ACisShwoSp7F6hjrJQns5
ZxpqxnbFynNWGdNs8bCWqENGnQYbb1ySBvOtpVHylVe9EkrPOo6MTorh15zAQ0jjB+sE3l7Bowr9
HDCkKSHM0zcbErucB9rpRclUuSf8W3gavMbtByUSDgIkCDaKxq2OWwFh84eVy53tZM6MA+HfIO9C
PCXi5OdAScMMxVDtgyMoL3tlJCIE3/kktydqFJZwkCoBIlHRG/zLTVerph446YK1pRBpEP36FUpF
YtZZtIA2nXCg+zCFs7lj5pihxGbrpuC5xLvGlBeZ0yp2YYP13NhJ+kYqCtc1QQt2+kKZKYmb6LO3
019hDFQGtG3h9lIuB/xrVdwGN1BCjfWWTUfomDyMb+tftXV+X7NNiTiFV4k4bLe7qAhCY4Whw7SI
rD/a98WS79G4iwZShDhT47JTI7jqHXafGCrqPlvO3zA9Zkm6rdBhA/grwWFJRmLQjyTFu/57LG1v
tbxOwFH8POZBUC82VwVCzBhTvW700aVpHkjnTeyEJcnrt9P2oVwKF4r0163o/GtPOOOxMmfnd9n/
Bs+UMA6GBkoGaXkgjjrjuK6OvVOM2G92QmVTcL2I8R4TQGTCKcq2GWvvR8YHOUvG/iKOy+ga3W6S
+qTFEzGy9Aj1fKQWHmA4F+wYYuUXiu/vVDlR1CX8ZVOMzm/En1qjgZTkBUqZztLX2gpW0ldF93Fs
gZzfUKO7HQdkxvT9xYELhL73NWyOoO1+LCve/qdI2vD6S0SUdNrK2ikNBfKizQB0wByp1pEJuWEZ
6SWDj5tuO9ByxoJ26HrF8wrfKLbsPWwGpJo2a3KT/rt1LYYt8jeJbTr6NrPvJZsXvwh3epyhRFGD
IO0FS4bv1QuiMnkDvSgPqnh9BySUJnMo5cALOhkp/DLDZae/xui/aS6sOmsUjf8qPBYzonEi0v8C
sj5OFG+1OYvv6TJQwO1U06tpqeu0BknbJFJXbdIlOI7s/78PQYYsAyk17pNwu0XO5OZl/VKZx+Ok
AKhoQLKRl5SIaDvcLWc9GFa7/3RUFh/Qsnmohvwunr/9Mpr/RUxrEaNM2iMEFHqZrSAM2EBhYtw8
Jkvd+ytIWcD4sF5VVL93/S9owEj0SXv1YE/HIBbeUTzUUpmYaBfnGABB8YOaF2p9So1jAUPjwGJq
32jfZajmvTaYHak/PfC6+C1Rp4MkHpDQ3JCnbyAFQB9S35/XwCGQUolCkkXgi+GHdzWsYvRmVvJ/
inyLmoIec7hUpHhPQBQS2arLfS6/bAW//lMWVJH28hG7+1Bvu6POzBJWU2mYnmf+nyS0HP6Wbskj
4zfIQdtCbukV4n2HpG9RFCQIQiyzsAZJ1Lq+0uYqpDR9WwptrX7Z8l+npoZFT/pxq1Tl5wBOMosh
6WasgIxlJkd54h7RS9fN4tUZAeQz98WznfrtmPYLTCF8HFTED6qy7UL8MYIw7PrGi8/BJK2mLkbW
ecsXW7dnn7iwk3ES17n7719IDtAMCvil/CElzF+PQW6dHZoPCKmRf6z2QfSG4gZqmzVTy4KMGvcb
jVrCkf+ofyuVwjGcoqI1YhqSAqAZT/3A5VJmuhUkxWmYLDtmiMzbGuh5JfLxbNlC7bZeAl69ybP0
OjAn+6Z6iijaqfrUlD3naLGa1OFcF5oStZ+VSg3tgLg+AhLkBTo1UrGDx9iTyJUubOOMRpvUJJpc
oOvrFAqlLjVNfMhI5z4iJIYeywYPJqLlGoHZC/8V9m7FRbDGxlvmGEO6dWD+9tmAGBEtNVshLumX
vaJE6dk3sLoYh2fOmLA4vJKjDSsnl76/oQiGApQD8nvsWiNWTNs66BQlXQZ7cN8DyTJt5uEpWmt0
XqniswrjDWoiyWTbvvpYQPQVoXFkh3JXLwOa0JsjN66QBs6kSCmyLsbA2kQGOOZ0mJBQy/DSxcDW
RLarPGRDfeVSSk6v95VcyPlxaZs5r9W1U7Xi0CtHor2eNSAixZ1cmF+lJBg9ieSmUoM/JX8Hc9bw
fld3yRMMjfitPTz/X6gOb5AGuftDylcdNWrsVzXbzE+OoWAUAoTXtBatCnL8NayRZFhR2XsnSQNP
Yg5lMlvY4JmcZ1PVLEqtcduKfjug6iMIpxXqkqX/TPst3Fb913FPeOess4GMeQEhKNthonLdQPA/
knGTGLvksRmE+dc7Qf12aRaYlp3gdVzPpQZ0x8kAu94pVzzo+S3Amw+IqWGoBPXr8laS1FhtyCey
3g6EcfHCnbaj8SgUjmf8fw2sXqtV1/2kZTMip/fTYgy26yTau30xSIbFXWt9CIswwPzAFPMjyykS
xp15WfyKgDr7ETa3jmrr766ILHR75C3GdiPOGlqlWAofrccoIgt0avK5e12/0Adc9Ihl//HOpoSt
RIYznINiLtIQULBU0/C8Yol0Kk6dyn17WN95UXzX5bZ57K6kGPiKKbgoMp672ZqVflxqx56WjIsr
VycmMDi0IP0/TGaT0PIHRx5rgbKG+jN0qAl330WlrYsDscTJDLZUp6zit3xEI44IAa3H5vdqW/eI
9Gsr9U09raU705mWn2RHn1T9KnElH+ArbFm930VUgHLaB4VhEhOuXde6HrN5Oy8TTgCzH5iyg+h0
Ocns5gKFAyXQnHjIpfCV/9kYjCbbBihylD2YG9V6BA7TDPCIWqRbNEx4DEG4q1vn15QWGnMnnqNT
0bXrFB20DCwM4t+Hsl8cFILuKRcW5ZAcs7GikJptTCalCfPq+qIcGFDaQuyEA15o3MD7ycpyfeAz
aODVxN9omClnPs/SmeVAhddWM9nC1wYUYcpma+VuJeUv0lmzDIAM4VZYP57Klqz99sdVZbBVumKA
tTP8kiWjNCovGZrIgo6V5Nqtq27E/NMcju8ClGKU3QdhGCp/BR4tC7DUmWZmVZ2tCR8mIWX5dIe8
9zgdfWYOXyS4i9chHncOcZ54kM4fL64++T/1A56lhINPrOCj4ERVH/Y6nQvOn3hkYZckKteNpmcO
enrazsKM6+FcNhOsE959jDAj9BVDmnHBItp1wCWkubqf4RMJzyr6Dsw/GrNl6YnPqN25iHyiM4bj
F/MsYV4Yudoj9FLgLZBNQ1onfa8sf+NepMf6r7nyL5e/LLlPRKHIoHD/VhI9Hhh/B48q5D+cJP+0
v5P48OrMlzm9QM6hi9KEGSv6Dvb5VmO8PrJ4wh1y28cl+NmNsKyd6DkYduP1sW7HjAuWyLFYLeLU
oMWXX9CeSO//FYF1jxkpdWrxW34Pgb6jFgfe/wGpTyaU98C66/MkRpiBokpWRvxGFk7Znj3AWq81
G27PgGQwFB+CZpKTbdwgp1I2wU7vjT1jgve5OFEkueHwC7wmkYdU2FwzBhwcbokSnupLT6eHyP3u
in2IXAKDWHOtCmvlqpcS9YVvGK04jL2JgI4KSJY5nvdcaXjZpd4rUlgJE/QOHy47aMreove2GcOr
yMUhmQ0PHE7yZVjLwTPq3Wt2gNFMnStaOEkE1OFFp/WijBIIszFpFxa7A9tTYYvxcvwWQuvTAMnU
GsloITJ0RCYprG5WidmJZ46iCP7i1QS/rqAOuyDuGdZkhfvHCWgJpFdp49oZ5IICRQlqvl2LoZJs
webY6fGRddoOMIPoSdWeSsaamg6iRW4eHVpPgNfRi8Jkie+SEGQkTMM/FEKIVLEHrLOa31NZglRV
lt7ub0KbEOfivwxPMGWiDmi55ka0CUI/mvXA6RlsWOx7qczDj06Ak+X4FpJAeY851VAxz1XB017s
prE2gti8nYJvPL1JD8P/E67DRpcuE8seyF15+KmMBKfvgfkKVsT1cPTjbp5rjBdyTzUsYklUCEyH
F6n/CraANA34Qa47fGyuE+RWtfrpq47EpZVI0LiypXuOXPC5M2V562v+A72nSAENCainQLsFd8hb
nq6IFGK1xMVwzIt48TqbNobKd1Dg233JP/Wd3NusN9hQ5rdNQ7r/k6JpTwfALPytUikZOS3u6ZZW
t/Ch7GNRjH/eJkHFiRU9MfKFX8qi0enzQRY3K6UWGDoenM5nGRn4j5cFajNj9h/G7acStMFmnFQL
zCl7qhZ5+i6z4CxhPrtB1baY0PcETZHORr6Bm0ps5mzQUHDe7lyZsa0DlTvG2T0jwtgk1yJMqKMM
mwupUXaxBUwHR76lhaEmfjOaHLB3O/lZx96HcGaFtz6yXTutxr//WGWx9oeavk+pgpVF4yuuY2Ib
MJSGux+RZbx+fSv8QDYOZlGKIeWi9etL48yJT3bGFDgFc107u3CsuQHitD/iGjt6cpVAmX0K9AD6
c8aT5NzYUhLMHkmzHLNa2X3+RbwXLCFkwqCjkj4teA7nZleDPCDdwKeLcks6jPwmEF5PH1D2OXbi
xDfl1CvDxT5lGrquIu8dl67SyJb3EUXAbJnVpBZq6bKT5bG2Xwf30Om3pbMIkopEpOa26odW9TEc
45gc8tQiROUpfHBShks/fTMrPTmxrksbVKE6yR0/gLAPytgZks6voMGvIi32LL765WDWmupVa9QG
lxag6nVgnqfbFd5V4Ypt0y6KhAYZiMAKl7YUDE+7uwv61aI08crp1I7OQaOMaP9TbGdh/WXOORV5
tV2+e9ZWbYFYOIq08COqW/Ioyw4NTx4vj2YSnhmj9YY+z4MCVCrII9ImRAbfqCp7yCFJUsApkBVV
5vSTejDq9SlT9nJF04krxMaaZ5cCZnZsUn8hsS3v1/Y+s3VHMUi0EM45Pdo8wb8ARxGKCyTxSzy7
cawon/3fq9NuzGc3sUKtOu03LA65gqdKETM7+7aLNgeyo6W1GN8wm0Uyl2MP251qUYFLVeKTvmNE
EfCsqHe5I5HYKl0afXeHnQFLvIeq4UY3tC/ju/ogaBv2hz/Rqb2r7GU4AelhdwNGIYEP2kFgjWxd
k/QxaUnsMVYK1dWc3rtfIZ2tKglYlewE/vEDUEjlht/CqzppPfOHWrsz+XwaPWEOGnd0EEKAivTP
peIkthoyPFoM7ZMTY7+/C+W/lotC++CSQ1Wf0YtBQMArLF3LnAraBDGFw6yOQ+TD+f7QrqaQ/neo
QjMYncAl+NwtffPEzshBctqrjxVkvhpFkZqwLNEIydtvZfDcTJap3pzuo7wNpyPQAbxzDeZXAOC4
5r1uLj5hSnBdXJvj5z2v1KvLEYA2bDHKOatkSdmWGKY5vdwh+Ql2Xs0HyFucbexX10Eu40iRag5E
dbs/g8CnC/rfoLmVVdJBW/Rb/YN/EcAWgyK9G8CtG9PebRL3NJoA7gNV4xJyT0lgXldeFrXKqWXt
eYGgF8uPmlS6hOAflFuD79sf8ENcwuxWRetHDbxlKrlawFhnccxX5Ig5auTo0/lfdk2jflQrNRQd
IvEwM98JqxZUWtxhjKkBvK+JnZBDwBhMLWnNxpqyoU/Qpg0omrEnnBk/9xNF4hZqtASlgPpBo65C
7aqooNAmMtG3RvTffXnQbMWCgs5+UbHJHae+Cx5Zepix82I88PnOQcGpeoK92z7zzNKKVWp6HUO9
DxZktvoRVQKTqONHIPRp8Ed7GeKIYhCFrFcxBSfYGhR4z3LwN5oYNmve/601WFzEw/humHufb4Ht
9WL5Wa2RyGsLzS+qhVv8UOewA6TjvRAexkiOjBGA6y800WlvKc3oIZs6D56Zpdx+b20qsR+Y2vMR
1KgmXH/n94JLpK1H2L2rYrK4kecZD0sH/sUP4UER7MBkq+Cfyh5xTOAzlZ1ryJOAPWC5tN2+/jvP
50N9wgXQ4Ef2FbftpqKRgraQUP2BbyA+9kiAXfpclCcWf2AGH8kEpB7ihFrnkqpgjM3cMdiI2BUo
2OFjLr6kiM/ufKp1M+Ka0CLzJ5g7ChZBoKdZXeW+mpcvcnCOfZMdFhq0LD8HLcxAmSuEDf3HI2dr
rJAM0dhk1BL1WYPAP75KqFwkCSoKGgCxyjhzT3KJrGt/lRYGYcuNB9swv/FA0WEp7w/VPH1yOzSV
bZWYoDdgHYbmZlSF0oCMi93kMTCwNdu0/vqszir+6pas6QOwEv9S6ACAtkf7g2v7n8p/ax/c3OVQ
gUrxtugnnHZ0d9OXy+timVBvmqn0NCyiIIuD5bfYp4r+Gdmg9IaAq5RJk8dhBd4GTVqyRGcz44vx
8FEyLrI0LGZ3yaldu1Atc09JZN9+CaMnsL6rNt3eLvcDnBU0LUDERocS5YavDYIht0EZkVIAxFZG
ITJopYqIYezmhm73yFZRdkrdRKWSQgoCzB8NcF+H+LCzBBICx2qRvQ/fEl5h/Ny5c8ZeJF8y90ML
RhQjlTxirSBR73xs94AFz4FeCEhgNYrwIB9IM0wZvLpTPgiDJ9nfyEieIq2qmTsk0Qw3VeU3i88x
6tXIXZJzR+t0od3bNx6yho9DoZWYsPBCpU39PH/nA+vUcUcryrs56LMEqBdTUjvRFuodgcuqMDg/
PjBliQ1x2CCidphlzd3046IhTvsMueyz33fa/3dLFLIkZq68CsNqDO5HBhmVWpb+NlMJ3viyYopy
mE4fObGl5xPjEbzlGE7Z8ySADI6tGQrw4gsmPNakFahdJnzxkWsKxIEB17YJR/LLaM+OgRnxZush
IAflQFE56O78SR2H96kJolPeZ4uvWcsB4lQZ8K8xOllU2hu6ExHDDUymTRjBPAcTb9Ve60uSVdZP
spRQpGIMVGB2qlljDxZopxnJqLnUfZPAYAiMmNTpC15dpBJRSsFNH9sJADTM+lOzPoS5/pjJImsc
5uLPPwb3AOeGGvukjz3GSwOmVBrLqJN3nCuYyU9rPd8p2elsCgJgmMq0sCWZCO23Fa1UGRwmfkCe
h3yDeVaMc17jleIeWAwoY+TcDKnJujucjZG6WzS2pA6nnjcGF6vc5rNwLCvoEvwslRgaYb0+LmDi
S4IiolzGUyVW4jj6cD56N/qVvhS0KceanGj56aTYqbtAN6TzvJ46krzQBgdZPbxjd6m0XP4VA1pa
qGOv4MeG25pPI+clGDedfqsGoYgm1LABWWHcYbisImKEACckDq4JgyEHXpQVybcTF4stkqZJd9ZK
nXDsC7siWbmn0viOhA7KgljKX+ZhGWVHPF1s2hwiy0xt+RL3yGE4zRpKfodCkwRvFYoE0QnplLkB
opcKakVsaZuw3G1dlvvJoeR0+H3QtIQLeRFaw2qbwvxRaRiJcPTod0p0J/zU/5VlPJdJQxdLKJ3j
nFng5wBUBM+hU/KkaXizWZP+QiAeoIoo2/YTokdot5WZdmXy6U850DIdwxduIPtgKIU9F1PqPeTH
fVEz8xZQLMUhQ46533hAuyZRw0R7Q13+Z2ujzWlsjP1ENiZYVGBeDno5qFc6eo/3xXUW7ev65rWy
CHhYU+f4w5rT13XC2P/CWsPppYIyRL1f413XaH+wGJzBjLO48SHiz9rkSEnl2PzKoQsfFn5yXIG4
WjAS/pQ30KfoB4mFsnMij6CDt1+SOBolP7NqcTp4tStxrymV0VjwH1L7lJp6w1y4vqPXRnEfpAaf
8T21/zNzdLktVB7dXLBSadcRO631s1iGMjSQM6vSW/Cj+yr3SYjB4i8/8JITnOE65VFLS6w/uw/x
7lh735NHlXkT+1fREwnuHA6KevPWjJoVztvPMXYfR2J63EZtvXfyIVyIJ8hfzk0Oq+3zbiRvfR2p
WQ6vqH978s5ST368W5d0Ew97/Lwpbb+RgSqCG/JR4ccR/r6+EzsQ+HkLWgalgkPEU1FyDWZFHPpL
h9qgnn8VKzOwmaSPgIjJP+7GKNs0hBVzduUC7mjvmalXITFvqk1BrutG+3MEGU5Q2gCIWEO5yzUn
0IYf7L9yN1n/OfWmKqErswSmy6dz+Up4Lp8XedTaXxwzR4yRrkC20j39WcoliIJHKx2q+FLjLpXm
NwbGhYGO+1mJNVfHny7Hi/DNoW8LNtoUqDMfgokLzkrI/aOuSP6D/60/0atJpjJ0iP5i4fwu9Yq8
WSVE+Ub4epuwqRk3miJGRueztT0XCtNxkx5Hx7p3yJ8gv/Qq4m1O92Rs6SWBrY1PKxYHZErg6fbR
7dHHQnFBWM35xxy5g/713wZ+gNGrmxrumPY81ZJv+J8OPoryjLMrYiJ9L/ut0zXcGFV5FhcYINPQ
Q1P1FR4NEyBFZskg0oCscoqvFmaApeF7TG/JjJATkrU5pSoG972WKkrLHAO9bBTWsBgr/o5w0gji
QBNh0Kwzxws8EwPBSZugJItNJ3RrXHz+sQ5Gz3p11Pcjub4dn2p5aotyu1c/QbViwvy7rU3SU5RQ
SumQmcFIe1bgVARyXwAD0mgpBJaxAls85VoYLyLOjnJTZsvpAVHV6th4Mu81nDj2Fzo6KpYHT0VW
7RHfHAQttrvZWi4+Z6+3nlrdpLUyX/MTCx8F8QFmyiq+eL0kwRQwHZyuxI88dJvJJjHOwS4M3hpf
n6/5sL6StyOFDQOuG0qzBkdjRBL0DMTjTbo9YF8YsSS8IF7Qe6miyG4hHThDRyPLu6kEMyqBWb8d
pXBvRof2ehPaRi0VpyN2J1XmC8tWtsBJe/b+9ttM5lcnN0FYfVOdb655Y/kqUqhodQrA2vfyJLte
VI2LsOs3yb50372RusYH/PuoNgMhVCuWipNMN3I91Z27YHSE61WkeBnWsB98gqyUe/l6da4j+KSP
ZH0p8xN6Nc3ITlKI48zXo+TSiK20uiTNZphuhiIVYYwp8kVGuUl5f7fcTHJr3SGMCb05TojDCa+z
A/jDx3GMV3vrW3jfG//ULVUxb48ubanZ+QsvC5eMws6vR8EdC7JKSEHN7D7sHUaVyqn6Vz7pY4/1
cpsKTTe+2lF0JHmKwSdrUrZXooYYZgullQ9gLqceeQZKAVG6ShYsb2GquD4YLggz2Ko6tZrPHtbX
Ad5wCRb5h60xHdtefL8nCfeovGOaVr6iQt6HHlhiomQn7R0tWZDGmCtcMNzfa0Pk6BdbTn5s+2xL
m7aGeWMwGEmBhxjpSbIkEAa2+Q51CJuwk2kz1nJuLxCwokAmZh5lCb/MNrFcjH5AZNKT4ajL2iAe
46BsLg2DMF2T4ZlKIv7c66z63MpjNF66N2zJwc6zlSg4FnSax7cDoZeyC6oJ2KShyuF2mt3OLE+3
dNvvrISmHmpsZus12VnHH0BFq5GClHAcgwpIaQ9w/honu018h97hjIe8lOx/f4I7HSVVO0jErV1J
qxIsXi+iHYXMGGpCJxxUim8lJF6nEAAwClnKc8PORjPLI5neM/FLGE/S83rXZfJnqsyKtbGSs/Fh
SAzegTACVJTWV+OHiryvq+0w89GoS1ub2KQ2pYHeNrKj38Y8Z1zS0b7/NU1bvcRdoM3RBc21NlPX
DtSmZfp19q84SaU0Uf0cwLBan2H04OuU8bHkDnBY44WZKDvZMpPZxGISN5xUku0/sZIxrShYxPdH
42V05cOR3yROYn1T+aRNVeKfVIDhTmaXxKA5/vJKSLvozhtsGHpZKQ7WtLPXmPdPBy+vPlVJJXJy
BZHbZAKxrksFCf2XtBg9/JcTVzDQWzXMnRaaT0F1Y0uZ+m42upAhQjesafg2H75UwCNFVi4PbGFD
LXHd9dhI71EIEOFjTL34QjCKrYg6513PrVojcDEKTMpuAVLsqqqiTAdLxKZBi+LdIc/XtndPyek6
twrQz+PzvP8YIxBRldJnQfuJyfw75l08XXWeOrwIScekcdRY0ruwRMy2iWC7zT2vknOa1L+GJ9fw
uYzxAUjNwWJV28IsKEI/S1ReIXEF/0vF7cH90krhlSItGaRCMpyG25H1jwgBg6Aoxg6Yv2qoHiqM
Aq2dyhmJYGXnMRPLzaON17+4fGCHVWZ9jtM4hCj6aOccR5LQ54yt/SgK8vNI6d2WgPpNpAfCU+ec
2LSa/wnE0iZhK2WhU6mMMXFHkOMJwvQQaCs1idSNZwALS9eA7IXk/4C5yzP5k43Ra2Vj9tyRJQF2
EaCZNLaUAK+n9rG1hiqZ2IajhR8vSbCK5GzpYz5eoyt9DKEsBH3H4t/bErgJJv1iJ8sbToTx+gSi
HthgKYfy1iFOBcUUDMzLafrMU/J3oBFc6kpkCvpa7hFY7tQvuI+mwDX/azoEk0whki+WjaxHiINk
ITFl/YkPUzRyOfLBirIftudKagqv+cL8uCRkv55YvDZp5qTqw9L1mN7pCFkOfWZUFnQPGKxMrP6u
gtArhpL8gaRjLKQYtICJHIumkoYLn4dZ+gcGqzWEu3vFGPhcOGSf31j81Y05tu21CdoiWNY81GUg
MaTTphIImbST+QuJGsNAmTEYOCajCBsF8jhro88juOlhxJ3RnKAjzlomqdFFZxizh+IQOeqp1Ybl
qIBP9KRHSllgHQtsxv8tAnY+KnCRAJHzPaFAsvByyoGM4T5c1/UZ4yW1FtSh48X8JZNJaGgqbTnl
dBGilxJSjzdyiImbv5d4WG/95knLGHzMGz6Ch1Vvi5QJlVGsS+fpH2mz3nPUr9LsVPhMfsZC9JpI
2mFlpiLZ62+ZQvv6HEfJzyHMA37KU9iiKZ6veMKgCiZMyR3KpeUmwGCkBXjB3RpO8/0KJmuoICoI
ugd4cackyU8kcGAIm/oe4sFwj6LX9lC1URQEErh6ZrMqhhfTOj2C4HFfEh126MrqL8zECIXHwrdt
H1IYkQKEc+FDNqdgGn6oNjSKJB6zNHaflV1bsW3Cz2IipWlgfYU4Sa/vPP5CShthf7NCh8X7e5hc
w4sNFTzsMqJ6BTp1SJHRi3XpL5y1TeUDj/d7CTV4Xiz0VxtmZBNXAyMpjbGELqnasQLS2XSIykVs
Yi4N0qvIhYcsuJX4hsXpLQA0AwSZLwlmqHCovAVwQOMLRvAd59tqHoHN3UJrZmsP6eL865Z/QnEC
VNrzRMTD+hN4N+h4T1EW6ebMUGlzb+JFB3ov639eEVNlcCaVOxs4pl7hEdx4AG8I3ea5plQIQCm7
bnK9oNsAQ9n6tpOYpKHRPJj+tiOTU5uz7HE5Vbtz6ubQ5SKb2q+sYR8Ma57nRi3oV77Zk1rBrmsH
dvUAQW9tVeq625SeYSOioXN4mdTUx1s3ipB4HK3KxoYg4B3+Bk8+h9uR7lCtU54QhOYoXd6ATPuZ
VmehiGCYmgXMde4Hue53iQYdVSVy6X/KcY5ndPTpeNsuW76v2WkqUUgp0JWK1mrogU1s4kv6ybNq
m0Uvh/wBdlGC3WtlKWNuU5bateaGQYHPen8CbdtWzoJzLeOTPDhfB3OEkFZvQ9QV2o+JWxSvfTlG
mMUumtMDZZT7YgQGz927MtYXbWwoAlrH7mrfO0ktOZA0brQMEgc/UAEpyqVgDQxSc3+N04w6VGsa
CMG3ZxsrmNZb6g2KNCbb/v0bbV3VqCZj68RwHdQgAwuaPX5cdXlN/uUNwX9BMqbqiGqXUwD5HMf0
hMEaBDw3oykxkwDavOwIuQ5epuhB6iQCJNszHvLSy+Mkr9V7xu+tw/HLOnHJ2E6j3rwzdtpH1dxI
4Akb2ZwnXVSCEiLSgBUBNi7h52y+PkUQp7pd1Y9hDeq19rq0Aihn8ULbn65uB7RrVKKXQ+qlxvvG
+74cE+kINIH5Et69IYTUTKKztKO8JCj/qz9HRmy15CVv4k+7mXvQoAwCamWcAmCCxj3Z1c0BTUEe
NdHmtmkbvHK/X8WtsEgYZUymVbgHOx1ST2td4TpNe+K3aDHo2634SkyFcMq03FMLrb7MNah34nGL
4TcWbtj9TEIIZJquRnhY7Abo32UjxMxmwlp1GcFouXcCM3iQVdC+tx6j2qDzDo+Jx4s392bjK4Ye
yTLKxr/A3oo8ECVA+h+Cg95ni/dumXFIgHrtSeJMhaNDOCNv8VKPfWSCGj87q8QWGt7ZsR44lL11
pN/arkLi7hRsAqr4lwIc9TEZ+//oiJlBm4rTQSKShO4B9/7qh0ScHpZZLigEItguqeygBLBrsfz3
2SLaVyQEIFJKqpqbgMoDCygPo7q158Gx1ceVuJ2BkHzZKwSDOyZQvrW23Dcp5s5vcC52Bf1dKQ8R
1PiKi9BwlX3uG7gLJ0tUUbo1cooecxWDw+b3GMPIdbdV+Sm4+lGYmsmNumFMPMcmE4XTGvuzEtAI
QcTZhpObUBAIKCCMWXMhmtY6lt7xY7C5a1cbJ0ksXVua6TMZHCqT78OxzkaHTVJKP+vMNa7mh64Y
ElV2vrWE6UiM4gkU40zVS5DGn+F91NOhvUrl66NWVSLHfL+To4YrPoVz9wuRfdE3ZEFnwehFw3H9
UdldLJztjB0rhifElRsUu7eZzTZylmTG/1UKUCTxVLZrTBEUG1ugCtcGb/Wp2eYqVnqMFEitcMBY
6BZ6qxvqx1fpCUovwQ4jZVEhI3uI8ksrSMh0gDd7IXoCLapBHHDQkwL2oXqDTx+ULXuBKMYxC1E4
FXsZdJbasj+rjudoJUMvTMTlrbnQVyzFRYbMRzT5hI4XyULgpKsAPavwou2jMp21bl1kZzgGHgy9
a55ughWKY0oTD2yR08ZTk9KAyqG5OltJSBD6xqkHyFQms6xefb7+sRx+7jc2j+R8QShyWEq8c35L
Z2SB7gsEdr7JH2osdQsJVdyDgQBMJq5wMw4lrIsGHwK/aZfTx9MgpZHwQXXiGrVwkpuulVJHwBG6
S4bqo66fcQscwrsr3rNnZVGYEB8HO2R1/Una85ibXxnDY9LMMYW3/wPACySz6xuZSmDt4gvXnhot
eCAD2KoBNfHhrcEoneJBkF9d+gBOkKWGthWtF3M6oCC445HIjOn88Sxv2hgb6eJGiFNfK/OsGvb8
E9Oyl/4hbuTnjmcyBU9qqu4ebjELiAW9tj0C9TKYsyYHM0G59ntwPNFkWlBHjnzPZI2aXIImIeQf
72kk5fE3zax8TDTb+VGa1E/pf4Ob9lLHWD7Vqtn+Q3F1Kcjd/7geEQ0wdWqDTPFZgi4b6mSyOfOm
7d4BAxjIvSCgYXvKQlgkAINe8iJ4CdKjCyOKSAm8SBMrTDYuPmVeIyN4CglcaamKwnLCvYCuqQsF
x+I31qsCBmrbfUWPMGJDeL82+GNc8J/L1Z8pz4WCok0AeozR6MaOE4/2zJykxHNSUu6TgoI52FqB
o0VYKeKnldmkNdlQZ+pLf7ellJexPielSzNiS+aNvOql3OzjPeFReRSyTJMo2ZzoU8XUMzeUA6H/
KVMyV9SNaJGxpBz8Uv34K3I6jVU/E8PONPWN+1HThR7iusbiOE24Cr3yJBkKQgacc488ZTLxg+WC
YyCFmvUnR1gYZeXGobKRkA+nBITfEfc6tbJGn609X69ZJzBYFlk6la+51cpSvBi6UNSQ3eyGm+Wa
Og8WZRttyG+NfX506G89AsUEMcgLeAfQD6uoO7HTGaVYKuqUGzbAToKXrXK+c1OlMffJIU71glLZ
tVgAmM6nFHXmXlpJAH16CSVthIJdwKWiFd0YEyqcxiZVl9ayPHKdD08cZnHqKONn0+qZRLsWBJ8n
Qc1z7leHpRGX734p5IRu7hxQL+I7Aak5qL423H4m/s+ZEY4F+2dTO6xsCLp/2Xr6PyNUz7XpTsqz
Nq2YyGclqVgP7likXsQyC0Pic2A1tYhNy588sc34EEdrIpUTWK5tlsORuhMgx6TAF8dIWwF7hSIJ
sm4eYFv28gZsN/5rHT8czw7lTzLLwltgDiS4tjlRug7ZRJVPQxT1if6ao06mLxdnJ6edPl3vz2Mp
qQLdeO2M6W9DAtCZ4kskizSTD3nl7dpEICPcswp6KiyDwiuHmDS89DZOzfuJm/3eTB/Ow4DyxY/9
mHd2alhrPlcHgvdxSLK3Sovy/Iybje1uc5fYaqVxkYKt4YP5pVGDMZypgTI0g7/hkOm5PLPLqj7t
X8VZP2kYj6v99TbCWznDyUbSOmCFVjC4WKFzxCoFlFoiB3/tq+xj3SnnG/Ca9o9Jpa2/LfB+ZKGb
mp9LPskcvOZImR8IaXSS4s+9jNQ4RcS6W71kH+5gph5yL1ksNthfjpgw8NjW2rygyULXZtIq0mmu
btXfVrjQiH4kloNKEgZywaAgdqxzEbrjBP18cllTMjmD38FSZfwQTEkTKUQFIlOYrieUM+HFFdwY
vYD91Io/R7BXcZ0Xm5dqseZRwpAEEUjsyXhdCnrFDH7CO2KVZ+ekJNT8HGQ0XkcfGioIMIenE2fp
kmGEEL2Y9wnbV7t3ja3p067AoIa9ZeNT4riFLvEtssGR6MJGqXiHCYXzvB+oVeB1hjPe4PTsCqvp
DIVN5ri1V9AIhZkmy2DYxj3rMjZMzWS0Itbn8QWxPmmkv6e0RB6U3nefly0iPdovgqkAQ10DEvPM
2KeW3VGL7XjtAl0RyArBxGl99G4GqGMvZkG1WVvGlWBI9iYTy4o3+EwWpVWKOAYds4ShcBUMfifX
tgwLbDihNFM8ANw1L3L3NSDfs8sU1ZOUxoXRCNO3aHwDBqw2Dxc9XjZeDUrlQNvIVaXpw4s6P3cc
s1NdwceRUPuwg+d5xnMpPQ1Sjz/3XlSNAhvArl8c3p0yjRuyv1+w4aS5ibUUnmNGhha1YznUyhBO
cfHAjgJPARXSjxRdZxMxXEeF/Xgkm5FL2rNlEOhab4SS17QKEIm7VUiMkahv9Z1tXLBmjmKOjAH0
4GhLlNSY08TKAOJByGr+jmEWFu3jx7s4JtF/Ci91bO08DubKkSWX4tE3u5xM+voIZLNmPMLpwGQe
xpUzT2mVrarplgFZZBcaEQkUH2d59/TUgy/ndxjTdfdFKp2ARMeWn0lAOt3rDTm10rLzJc9tuy7v
YFwLOio9ellmu9RYH4SfN9+xiOH39uBPygqvqH32kKaPd5MXD27cvsWuLMHyH5WYGLROxN+UaXrs
ghiLWpmJJC4s+QkecMhXEw5W/9mdUQTNAs9I7EfCkzsk2AEfxzZBElKhUoI7SOP06585X/cmHQ8t
fV99oEtl6tKvFNX+bwEPjotBVwaeOFz3Kmq+GChoXH2DVKpMp5ys8vZWMJqbNFuWO/HSzNN5b2sK
eg8tkKX0bRm2WvNTxQmdkjxfJQ9QWTE1HW1IW5MVS7Eh/T/M16zeSugHmZvfDUF5fl8ZUZV71gFG
pr/95g+vcuD9XPelF2wh1WQtHLjGEYsPMJdNmCNSpBCT2QIb4hKMwxWBdyiYtaXUL0Z3DXUmwe/1
PQk774wI/laGTGTC5ACT44zDzpPqIGLix0G3u0+f3wg/8V5C/1uTVSJZpzKVnerGbs1Qeb3EHCap
GSsc5jLBJE3Zf8oL0VXYxSU/XpQp0HRwI9WghPBmHO3RmKnYljo+82F6GOtJDGcdnSvXnYYW0P0j
8TiedVnxUKuzCFBv8waGhb8gjm8L4sMrcToMcXf7THZeH+8Avgnui+UEVPuP3xNfMQhlBFWjSqzc
Gp6xbqc60Dan0V9hNwc47rjQKAq7QAWyi8GEg1KG9SgsW3K+PwnbLExYzGPdkk/+O+Xpm+rC5bqL
7vhFWj3mDu2ZJ3/laQTvcI1sO3UNbsNCU41LHSrxkmpntU1kmiw5wdSKQJ8jcvAqw7OwekbSeJUW
rtcqQaTwsAIrWNSxwnYZfYTgVJFypjRa+pNLGJ7o1G9bjcS6Sf8u6RsM8JHnOfYxkhgKFx7ne/BB
G1Hn9PdxH5OcOVyNjcuZjPZxnn4s8aPsNGLBfw4t8eFeplAVc/tWyFadMzmILBh/5SBEEeb0TFhV
RkqIgZPhBfCMv22mNJGwHM+RH0IPv2uy8oEQgT6Aev5j4ge6ZeXqev6R30mHjsqu3L1Z7ZIaxdzR
qzMga9o+bJIUcYW6XYzgNKvGRncDKDnC72XwFiRtHMZ6vxPkaMSeih2vV6GBVAzdkN1x9YWblppU
noQ7Evdipie7kWAPPjUFcRLsKDjjEsFlLdJ0r2aWot2W325fwGSvK1Rc96HPbes+sa1LrDu7oHXN
QRmBKy0UaLrPQNR6dpTkK32F5UiBIIgTmgAMJDc9JSKuw/R0KvkGm2mGPx2EXiOrz42dKwLga08w
5pOeAf1OJz1l45iGBkG8t2PKQbGwPoxbQtY8foi7R/HdcPeg+tSAtqJ9DSYnKB5+Gp98Z1A72Scx
YkeHToOu/9a1csxbyHM+wpe7gwdlmPxCh502t2JqC4LxEnocw35yM1g+glZwTDyte+/T0QEeLbr8
uNyk0ZJZlZAsZ/2PWNRJ4p4rX5WhDrHyxCOC52AwllpLqURuRiahk1gOjtllhLHZEOVa6VQRLVeC
Bc/Lm37Zmlo1xoK6RIObSCaRs6gQn8fNThPVUVmMJIHlmNsrwRUb0oyoOM4mJBNjhEyddNFe0mgy
SQjCASv2uPvWXlsFcQliNLUhUN5ldX20hzXJiTF2u4UbRVoCqYzywRHv4y/xwMqsqZ5KyAfRIdhI
L8GpHuJwSwY0Tb5wNFmYqDVoBxeWlcknvYo+Bcs89h4l2Ili1f4pOamMeUO9rTujRGj+GVhlBGbD
HWx5rGUKAISLimSs09if8TEn/k6d8Wv3dX5ZvT+otSX5uwoq9NWjZ1fGfQOI2bpdqsBnSVGY87hv
3rwUUIqHGPmQm8GAlkiNoFAsRtSg9wgTT42BFa3OnGSRT9aJn0xqiAo24C9ujEny4MnGr+hGKL7q
Hxr3lpNbUeHcScIvPV/6BpvWue06iPy/PB94C7NB2F6Td2xQVnOmW24MVLNh2Mf/rmGRFHOyWoUF
TFXi3qLk7jrUO8zsYBuMGEe+h4tRMS44aaMo2W9QzK6ZUlQnVnbm8ibCKdoOGK/jSb8qgWfDxtW9
nNB8WAfvsLZA/ex1W2OKv7CIyMkDBcbt9+gh7fBC6IUtM22KtqWFyjV+fz8Hrt6VQibrwo24oEaY
gKsu7CKa9R0SSiS/EXMCDUkwfJkD1zOFOdxQTOEiD8x0fkrqHgly6P4LYcrrt5HLhUgi+uEYUfdf
l9rwl7EgqWHpomTnIXm8zSq8DsIhHf/1gC/IJHOk2jNwQAP53Bi76TzxMDGlQmLCcVW077v8oUmB
DQGpp280Y7PMTmH1B/W2Yz+6i+ki0VEFGWBnoiRdevdrIWoYIfhdpJvERYqYYpJWO3fU6/TE4qQE
BxCO5//8uqKUfHZrmK5vC/AHl/O51jCNQiWwVyUao1uUW4ELj3qL2Bc7LBbyGUFfWRfPqyVa0t25
NALRW4y8I9HUaiVRONbI56nQTDgXuxio8IGkTpyFwP6a3BeIPfRD3XCW8Vzv4kJNQXtfRcsdu5AG
wSHCnDZn0azWRF1scyOHG1DrttFVggxVJ1YuGv8JaXCe2uqpTjXJqhLmRT3jQSHm+TL+oHLfV4UT
/b5k+0xGyayTuMdAcgkUvmiGeBmulG/er9M6byiCPQxUM85KOTTtZvpEyAk1/xn30K1J0wAIISA2
LRz3I/xV4lQk9QveyMNBG0REfpWo4ko1O3Y5KEe83Ma/aYSrdHThPsqOXWr6LUGhHCJ5LXhilGie
8FvBzZaiGwBP3q5/qoMoa+3chf/10KZnFbfUmppv1dWJNzgAy7sYtZvEGbacaPCClRLA8SASeNwX
xeFZUdyhWEwFllVFvN/jflR+pRa9TGHZKYmGPJEn1zg0/DncsrvrA6uxJMhbNBAUE9Kz9umHHRrO
iYabcj4WnUhst/56eJ+bNZDn0+jFoZDklqJjcu3U62JKKO0fJITsOmUweGFUkPtAJqgap4aYDbOD
nlPr9uK/FFvQiK48Qf70dHK60NGV5xPp8+/0J4D070sES5KH+eN8ol9Sqp3n1qB0zcelWI5Kf6xQ
Wn9RXJ5bMLMh2SZfveCfARb21DlRDPL0lpWD7PTL2dFuz8WXZ544xzHN2ReSbO2st3EgL27VY5dp
7OnDfK0OHsZmo7+kC7LqAxAJGFed748vOfnhn2mQBF1mZLXWrWW/iq0HbeMORSoMggd9SAPjN5iu
z02CJoLJrIplJ4F8nEXNIw7roUQlT89goaOtvNPDqxIr6dmQvqKv2kWBBNsxjFBt5RBQj0UshIz9
8Z+928xr8nJTM17vmfhapJvkhjxrO+s/TJ4tDA/gn7BaHsPgF3MoGZkPp8t+ePGRQ1DYgxV0nW5b
NaTl/Q/WHPa1/QkwoYEoRf4jb3MiXtAUj9ZtQ5qly5KcF0IXzpeIpPC3cJVT75Ra4++tGx9zFDiP
/COh5q3gryPYYAHadgpkTMcWl0S3vn1LRxFsfOMbaY6+B4gNuUq+MRmK7WdnSENCx4JQ2pzYz6cD
f5x9+FGxmYzVcCQI+GwdVj9YpdohSmnuNezWYDNokTuswmRhKvcMahbPgLk/Y/untO3Ua5ey3a0a
HSDUS857lGJa+3iYjuTaQDMkO1DShAhM8k3zdu0rQfNlxnYXeP0i+kkfT9yHJcbRwVaLqyClAI66
ov21QMciftGVS+Rk346rRv1EhdLPaUaCo52hYOUXfZmuysk6PwZygYUUcPEMoI5znkjR+PLo6zCr
dWgaaSLvDP5+UHdMXPmEKOhBUXYZjeraXTK4CMKiKYIRdsxZUBdqKX47I5TY4lV2bTDq6svfer0z
JZ0KcyrAzR4obYaMKKyhTqekeVhEJdOtjAsJMseB868gcZGTtFLErEvmgkXn6d4IpXzfdo+RuOYH
KgvGaifYC/dKWz/1O6kcFWcPlbvhAESgU2qBcemhQ0WR10FFmUH8dP5O+CQoUfd7B27zupU2DSwx
9cGCjOc/YTFXrSt3cF1SfBvpg9STuYFWHjls9Mbyfug0lWaEo6VP7xsNbaQ0YofdEARRP8IK9M30
qt/HtAA70mZmilP7dvpx0BPik/0h7gh+QWRgk4mt1O/9eT3j9BU1nAo9BPSIfg2xlfw6IIawipVm
fhe3fEMtM+RapYzE7bsUBDU1vPo8WuccJWG0bXSSui+ealY9v+Z8oQpHN+6CnwVyGv1gIunZIKcl
wjo+NegvmSOB3HCb8+idRXD5zH9cgmk8YUVwHtTdA+iDvOo80hVS7vTb3HRpAgAODwvco4wDSUHm
816aWC/BUNflkWuMtH+AwWyUpxtLC+GTbX2LI9daR6g/48bMhfr7yXcOz4W+SB+aXnKeDB9fINzT
OjbFeArvbfBzYoQjfA2Vzda+gjGK7MlQ1nA6n1idUA0EAdaBGn9kMRiA5OVnW437YQwE80vHLpsV
VjzRmxm7RpfDGIU5jKi0tgghYaO5SH5Uu1ptQD2m49pfbDYlpKaneu8cmWGe4nP5gM4o5iLVvspa
XxdychTZq6hcOkNvS1g1NilG1DTlGXDRfqfhk6im+fH0nk3pgUB4MVlnyuknKJO5r1taiecYX+PY
kvjG9o1uw4Uo0+JitRdCid7mTcVMSP5i+rnmDjZEd6EUqaIlo1RnyMk2m3h6VmObHPgadq1TYd7p
BNp0bxni308lbHihXr8wQfN/4MGG0i6aasnrjg7q3+dpBaNc15hVeyE9tLyBWN1SJ5yo8xaGaR4s
lTdaSfaVBwCSW7oEB7Hlx/22GnyN4rXG7IAXEqDHIrTENKS0AgKy6W+WmoYLEhOgg0SSMKnPT5Es
L8OzdEU9K96tc2myoQ2q8HI3F63bN+TP+kNUJPVchXjk0gJznOZtYKrLbUYTEy/Au4Vtz3SDGFx/
BuVGO772r7vpCd0Jo+SVUgrNQJ3wOPhVtLFb1TWHR6NLwz+uYwemrGz79YdAYnHlE9nA2m45b/21
ntSZDMnIod3cxudPbwZKVg+xSftRSSxGrwGulYew0nJ6RYVeNsBIqwhDXa24+hN+gadyOvCRsEoM
BzwhrRbFb7mlqVDuQzhoZtpM3qo4bStX+Rlu05Dw8TyJj86lAYMpLlb+GSLA5l1TFiAm0BLE8q7C
4g3TZRw9cHMsNdCejVrc6dprRqCwF04Wytu5WxxPn3qv4L4EpqwQqTf4ATkCLPFDNq2mJ+4AU6xd
OL57YnPnV3JvTS74V8+LKcrJvDcZAVrfqZk+WWtGxNBdS6rdNGjgB7B2feqXhwuOgZMuA4Hi/XXN
V6S4eUXkv4n3PyuXBQV1KdCP75maZ62Kl7RjgSOmW/vXeUnJ+VI3gVwqXcccut7fxteWgvJyDRbp
o93OG4bi4EdA9UnbwqQQwmVKV/9knSVpF0FIjfd3B94qg3hooyl5scM5d4paWa/z7vmwCGQk7DrT
E5tqkusvAINEQxSqz0STxqXt5Bt4sikuzWflLQJBG97hlXYsBWkJksqqmXYl8Hd3aIcgi9Dya+j9
onOi5h38QvYl299ORZ+iH+lyhrev8QjZna0mFDZ3DPOPjnxj2vwHtpZt6C7ac71SFlyxsvz8eeNi
8CCc4ku1FF6cPylSSf7Lj8STsoWHHfBa7af5/7BMH0BN3Zb0drbSzgYNl5W7d0iS1+XT0bK8KS2S
RvCzLtzc8GeJBmn26c2/qG3TMvq9FVCTmMCvnPJ5pKld65xwm0J+9bfLi3YeR8s51EHWPuB3husf
2oZmfaoGsM8DUFanTkHCki8k8KtTSGMsxTz7Bjo7je+pfFM1EFBUN64I/CG3fq6zuZ2CnBvb/U/P
UggOuMMbwnZwztqvvICC1bDu+JxZgf7YxOcWEUpbNGarQggQMqKMDTVbQ0lpLY2OWfJbUq5DTNdA
gErwGbDZPNLY6vPIp/zPzBIQOcoXfxJ/CzQ3PdCKM31r5+3X1smJcKjRZmyKbd+2/gjvaQ+OeMKe
l8ybJhvNrlbOkWCmNyurkVCi9MEP4HKphohrdfj/Q+kQi0fzcHwipbg6v1qXQ7C0I6gK8qkJcX6R
Vwl1/8Q3HOlGdpMTU2Rl6CEsfGG71sLXOz9Hl4UPM4ei2yM2dvL4qjw0FjaBDacH+MnaWAD6v4GP
Mopw4KcOBgW3oV23qY/kU2MOFWfrSVdBV5b2CcO+taH9eMbAHTxkBvE2+ka4IuiWzwT5tLWovOG2
Nr/9DFp7Om5JzN/pUx6Jd7B4B07RMFvG+T0EZ0e2I8kNnuHoV7OLhGSzb0p9Tjm+a0p6PapuD76N
njPKMVngKOcfnNg2/MN8fykSn3a50+Rq2ZeJJ2ZfLUc7Jpkx3TCeqLGBJkr3qO4yRqu1jpKYVAQ9
fK1anq0SSvG2nduce4dKULRFdHx1MATeqDtFABjHZ7CiK2nlqbmETVa2WnGssMlpeyr+j264SAr9
ON3luAqJSwmNOlNgijIL5+ELlahE+Ahyb+iZlcP3RhQSjfCEFQrj881khLmuR9lFDHOU4hHGSVSQ
OuCz3/xCTuk7csArdcjkwG5TBhnY/PyDKCkNqQqVYWFTJKxGRY2WkVgcfIJRHqPHqc9XTydA+P/p
mzszBuz3Ck/KaffRiHrXCiGPpMdOQmPoYnHokMhUYf02b1ghiyT9H14G2cwu9L9P8JzHc57IjPPb
sd8ityGkdMTzCpm/NzHGxEAI7JRqzHP5dHjr68HD+4I+CyBOHqTgXdZunzfF6zD1QwtbU938CZJU
YxNj9g2xukqtA5ZWRPuIzmg/qybJydDjjWlgZT5xep8WOR662N4K3uFxg7MohtIBsCqTu0yiYo8q
F3fwkCs6jeLak/mYkt7t2cBXUsKGTt4mDQPYVVKe1d2hKlbgHKG8yQQpCBCubnRdcGxIUuI0qfvE
/lNbYMcS/vfumNxpQ7HTJgDnG9tRKKAyHnq/XO2YqRfWScAZTNfk0vcxugGhOYLbtEQhY4GCuWHc
4/fK7qjvthfabCbG5OQKbznAdg8pitv5X75u6tQnVyOW1/QUGwzZUVZ9tZpX+fuxL+/z0Pq4/W/F
FKvjsfTEHOAVbFF1Tf/Hk9W6zSC2yYb7bd4rsHYTFdjOy9C6yc9LKH+jDCSGogWQ4AX76Ofh5scb
EUmEEsDXt7nHsZo3mGNfUshRZdZPmLDOuxGtbdYhmHKqfGZApMau8VWggVD5Kx2zEfb099QmTa1J
kft1s8GzQ4wZpgPI+tUM8bXQNMdXuaz/8bn+VYKFol0BBd4vsIYba4jg7hgLDRG2DVcGgiAae1WN
E0LgQ6fzUG5Z+sC0Kx6QJmPreXl5sulILhX0cmxq2jF5DzyO3YiHGShGl4TaNWYDzGMu0dToZeak
h+QWlR6POgsxc9Xg4BEXlJ2l6tyBM9rRY9Zd8bXZV3Kp/SJMN1rV9u7T1tZ5s48/guj9c6x9MRH0
NNDqI1P3YjNRWULvpg9NoYcK4Llz2QxLkaRDpRaa2uIDPyPVGwZSS2wuK2h61r0qgT6xd8kJbrTq
xlzD17BT53LVue58IyWXZX1WCRqclfOwipI+wmfV+W/7572Gfx6/ZZwH+2y6GNg1J/RFwEWKK2L8
Mxg83kC8hEA9JvVaQbq7dSJw/qJdUVO6TRCemAUESFOdHpoArcCk2xKAxtuDzlv4gb1moBfu0ehk
kwws+4tzljTzemJtmhRdjDJlDoMzMnVNc5se4jUxqFLQ/pOukSOITtLggi3QuOrpiwdbWM7WFknX
HKB4Zm7aml/HSjoDtoq7Hd4+jMLSDXDVvMrg0fpHJIz0s4Ao9qazaGtozWsEF4aEAElXXLp//oQ/
Srkm9dq9+X6EpO0ZMpWeKNBK7/ZYftneLmSY3dxO2BPY3+KoMMIxzmFIEUNnpYnR6gNfQvNACDec
aCBzEdvdwGdIihg4XkPHsPql2/Eh63Mn4WIR5zBIUrAk68itWn+NPmzM9EYhmfCYnmFwRwcYiGr9
tYjOK4uG5AZLXyLR/9Momt3TJIw2ynY4tvkiA5tbgp93MECSfBtUlR8oA0R6f6fWNZSlybQTWL5+
0DNrtKqH15Olr6OuYkaJvQGjkDL2+jt081VvABp5sPOclUUTDkRsXS6BkxyVHVhXIMEKunZCv4PH
mckg0jFR66Hz7ISCQyrws5gdHBjTx95a5QAukd7WG8l0S959KzYDOKnV8Us2SplkmQAxHLMVvCTj
0m3rXN2uMiKTTUt/jYd2+lNHOWPkHRtc9nDBBAgRUh0Es7WHTaJ833XgTq/R4rzc5HfF9RCtiSfc
HJbuKA8B30ksoDvLLlz3jaVDuLQhgp5CsW5XQNuwYFw8AUl4sWDFno4TMhPZNO5ZYrjlaScTH70P
/a1Yu3lCOxUwLw949tBaTAwyfoCc+kakzi1MHRDQMUDjusxUQYiKq+4lLNDLrf8RNzaqdT3pGjt4
PoRBNKxqfb06FR7vMp1sme2b0NVUTf8fWObRgATHGaC/wnSqXdqrw2rwbb71dFCLZsn/yruZeva9
honGWLE9oMp4nEk+VRhZvVkF4j9x/ae5cjymb1KwxEQVoVH56aRmjfOhOnnzde/9RcdK9R8SJ8GP
WvhsEswuD+2OGB0nThDEjPKi7enzj87PIh1RfZawFey3EoUrqG5ABm7bzFMUKieAc22T/hYxB8Mk
BfZq0EcDylXTEV4kI94RmBRUJ7heXm6mEdRg9kZXhxDxnQ4e2ECKtjKCxxzSwKYfS9EfE0vJ7hpT
lRFgUyyOIvq1YEspxBv93JgtwrKFfVuhp/kFTebL3tY8dbCXTvNXEK2BZDTcp4lKO/67uQBwa2pT
r1/Xtv5xx+E8Tbzdh5V3e/4tGiGWX7CQIAYGiZStERbGivmkfFMupXVD4If/iTfwjeaP3VgirYpR
TwVNkT8tmBjaIu9S6isuBCLpImWw7tWV771u0ihPA0Ki1kNzikx5ATEfBPVivQbGpzkUaRKDMgl0
W4AGpPk+Mh7aprowvJD9WMKxNWLIQSziToDaf11W3mWB9NGZQVimqqj9CYG3DXVGRUhORBjq7pTr
9eSawS0W2BwV3Ds8JU/wkJ5CWWwXmO+70I2LUI2qVgk3xIs/UEo0gsNQTiVuP42ARmgkPgcq8Ul6
qTitsFuQi9q/KPqujYuDoebhdFTMh6reqOA1DWZPh3Fyc50RTeCxQam7RU+R57YKfJJ4k6GRFjwS
lSuSe/MTOhC4w1vVSBM5fEYtZLxgIM7jV0bL2F3Tj9NDAYe7/GtdGW3DjCJZNKcX0eljk5hcMfbJ
+j+EYqj63pmgFXdmWlgN6wYGvi3X5Lt/ZHuasKLCMEcby519umoM00+iIc5iqW5j11gIj+DWx4jS
tO0LMnBkWz+WAZ63TL4OzGHPcO8szQcFroQHToGLOFq5YunfhI13HmmMTvkB1Z0n8DtwSRZF207V
7klcbOPfifVLgqbGVdPeELM9FFP6MlbgiuzCrxMGFoyGMZxwnBUlLXn3P9IdaB7ZODD6LJPEN8rO
nG+smmG9JizehZih5uU4g1w/Ck8SVPcfZJBzTgZijt2N6vJuhnD2lz+HAO3hqpBcnsg3FLF2I7E5
5PIOxSPKa67hqr6T4xZxr2JObi+AUUWIiIg5RVuWzZsOGjYWIENQkO3D5yphA49aQqs2Bwei86ew
LEbX6wJv8IQo8JiRPBSuJ0Ziw0fAy64zJvTT6ibZgnz+2Tj+7hO5/jP+IgBy8NufdnFHMpT2dCsU
CjaCUkHJQdYH58PhCSyJQaEqjkOHgotM4Y0VKVTuBMQNGCoroKA5nphfQt2Ja6IZy6/0qRMBuq0C
T+bwX7zArRVb06yOcZKSY16aKKgH6VnGBkrawALECR51W/2PLPY4dNpOBAxEaBtQ3af4k/iERSCc
A0+/kfzrY3XsguFZBFvRCOyzCLA5M8ckAOq+gfokSnN1sEbfMDbSwxOYljrU1MNDW5Ko2vooW6Yw
x28ieYFFCX4Qtj/NclvZBXSPen8weahiXwY7ksjL0yjq6aRLFTwbbxWZj1A93MX58wrd8xWqCHAe
eEBV3m4Cjh2mV0SygsG2NXTq8OVEj2EMC0giYinEf9JnWOtBF/az7qU2goEy5YYCnQBsuhTTN9FM
ZA4c+3/ZHlBMQdP4soWT+GnbF+fJ1c+WnDmymMg7Asxt+M1hN/XnTFUMsKzWrdTW+RH4n4TV4U0y
PB3Vj7HFuXhREaWKfoXoT8sK0SXkN2qIehxpod9viNBZZp7rkutaVw3jOgVbFJ98vAdONQqc95bZ
4YOgmkmgLlsg3h2oqwTeox2NmMEjnYTjVAHYlGWpPgL7PzA6cYS8F5gsT5cwRQg3C8ND6Gckon0j
V6pzf41r0lpJdOxtvFh09+md2jSGJZQqxax0VJyGxww8Ho5oZ4ZAKQvT8zC6YkUak6v5KMYOWZcg
A3a3vKAvFUja+rWRGfXzlCqXiGdYlwAheZeXkuDVcJrXRL31oXK2gpH2oBRvlcBOvTVD1J/uXbBq
crVhPYHt+aD6WUPnQSKsLsa9ihUZ0qCJQBKfmgyh/uvdD7tRsudNSfgTRLHqMiVDGlI2Q9JqlE9c
Up2WWFFFv+4A2KQCBdLCTv3Z0SZa4nLAayUK3QAFpKkDcerkhFoGXWLaXe9joeWJd8KXjdEh2TCD
nUAU/XqbXeoVipuTBtbegmClu6gkmfZEDKh/xRgahQJC1PpYI1pg9tyDTNTQr4T2xm3zTut2a4CP
hZ5QnEvQzGFiJBnENi7P7zTt9ti1aDrO+9luPeXn8x7B8ISe7tZOtgrrghgUh0Ob+OJ4/IbYLnw7
SZX6VHrJ8DmuMgAA/yZyh0iHcztU44HhH31HLl4gKnhLJ2JurMgX3jZgthcYXRNvVPYrfoFvGTbP
CG+zOB0+mLcX5M92tBq9UuShD4Hm9WOo9EskFB6a9X2SBMc4WzTjq/kB1i2Z22YxiKSlv/5l97q0
ML4qglT6JwPQpPmunnlon7svvDhQ0RZYWZjkU9gLWhgCI3EWEERVK6zFmiciWGLNbZroOR/SsuIJ
8jnwQAMiA0ic9fhwIzuNB+GOWuxsWwMo1BNQj+3O1t4mDUUXIuPFKZ0WqjTcpK5enB/Nl/y9HbTG
nzGOa6hrvF/tw9t5sVyPizB7F9yRtY46bcYHhDGf4/SwviEFnBuBXUxAjQSEpZ1EcPUsB/SMyGZr
sjR++owz4d345m+aj0ANlSZteOfCftC7R7gLWq4PjnQjKGZ3slousko6rP2wVMh7hYBPX5CTe4Dy
WCHeLUmnk6ZUlem8mWk0OwgnA93HOV+QUDqPsyvJXRYfPw26BRm5LHNIq57CHJ7LHaIKaaiVpQpE
gHLk7mVBGrS4KvsohSGKw+O4ccdAvhVXoMg0Pkhrj67eJjFWGgDZUiqc5syQFMpLNAuxdo3KUk+x
ubWmeLav00I1UYcVBVtsMbzPAzGAgx+K3ev6XOyfXkLt/T6i4/toGEbp6ewYG4E9xZ+X34oBptk5
+oCvOTwhL24V/xF/7R8H7nS9fDBx3mgAVwoA4S2ZvCy61Ff3SE9y9x6uZ+l63EgiETJ0PwOtKdRe
nCN023u+eNDmxkgjVg3Y37unFRHmLdu0Z4fiXSK4WQ4vQq7x9Re6uiVDDcEtfa/PRM/unDZTvOaL
bj98ZMXaFO88dLqzbo6SEgEZaBsAgeZz06n85XCf9GnQxb5s8eRreIEI6MsAhMGbnYDulqS9nWvj
C/9sPoXCFKDwLLwrJfwjaJ/Sc0gruxqu8ggYV13ZrnGzJ74US2yHE1okMMur4qf6RpAaVv5DN1zc
3fQoHh64hmG76dnFsGxppeD8VIr2zGwT4oO4jlvIQcWzF33QABT+ZlMMUMQgEVWIf0DaQpypXpiL
sFVzEOTWF+zP70KsImky/Wu192zjufR3SXJ89LSlkkOhe1jnhGDAPsY4NFNNZRSEARy9I8OxomNq
YoffnrJKTCYGreJKjc+RZkCXblbUSRhZzTbrseqFAa4K/iqmDKAtjiWmvISnTtalldvxzyzSCv0p
ByP4usdFiH6/USEYtGkSt5xtNIds4bY+vXnNmS6FYbdUQRege0tzYvH2ruFDoDc2ORWaAC3lKfi0
UooiVjhKCQJg4oMs4MDPockjMij+T7uJZABeKFlk+e20xAp8TknfzCgFyj1cSIZTNnXL+Tj3YjyL
GNUrcriUUNvqIgintJHlV9lW6QZ1dAmqabVMdN5+fKNC1Z1aJ0ioYJBvMxZiEMo+GGuD3CNVlpLB
gEWNb6cut2LqM+a7aawyz8aTSs0rJvn3Wm8Gb0puBgo2AQEC+BVvOdpuVX7NTgt6wvLbZHzh2M04
la3ZungI45TGE1KxcmlhnDAJqHz4FAfURAKDpsTaXOlbv2HZZ9+I5z6l27JU+a4QI9a30rr2SHai
n1pe3vFzl7tFExtyCNkD8utPn/M74STxbg1yzmm97FzJJuSahFs83ppkgc7ffb0Cgcmh8vHvLB5k
fAbyyKE9bvk1h/C2qKTQ2zh/zghJy1DHEfw3uUwPsTbHuAMSdI8XcdvahVY53daQOdcExSHK6cQQ
TZ9B5M5DstcnBIjJOPY3HELNYuzAdMI0xmVgAA6TUTTO4XN6Kfmg7MSJPxT3XTxFc/chN4Rfs+LC
gLP1oguyfK436pVGjQ7O15rgIvDCSYPHO+CSxtzhlRDLnsgx/3/tS51ddTtjodxJs2nJAz5dVW8i
8G7WAb1Vzh8HEP8eA9Tafgzj4mGK+ZN8zRQ6m1wUIOu8KuNK4JdqHH4xaqx72ue2a5dQ24R9UIyp
yGQCaHhhnT4QDa78E+rjJvK2TEzOsFjBbDaEKDmtdmL1CATBLLJHUY1Isw9c7COi/MRzfn4qQ13W
s2tfwflRTU2/6bXXVjSBWBNOU+fdinCttrVHNRdZIBlofgwZxTEKqKN3gVnZWFRXs7PZYgHjKGtc
Mcjj+peZJY9FtZ1cS0b+leEdjc1iNuGMTfDhYB+WNsvQHBwriyv87DZPnb05U9BSOyeEE31NG1nh
ZsHDHJFhi3HDF6a7T64dvmIDF+/G70d3y0ZDkYkadxtjGFQNsAvtXEnLxz4whEDW2nDQL+dxAdn3
6WATj/nsHFfu5xIjZwE2pDd0du9ndw+n8O8+kxSBQpMenfWzgM8jFHA99rer8kkbrKGwg38WVn2s
eo0gfw7WBDKOIVQFNXKmPJW39I1pRCDq3Do8ArRvOMryUk7pQVCMmNUE7Ab0OlJ9AVvYDwITi4DP
dQ2eWAXZAs2Y/nO+1+/WI/I6EgV8NsAymc9ZY0SYKwfay1BpaIk2Oj+GN3harPeC995mCZWZS1MU
X1JMyYQtlkfJiuakKk9OQQ374wdm1bI4VkcRD/zAY5o9ASQfEYivS6lSwdKn2hu9Eo5PlSqnbWUt
Xv6EzIq8qIRYQdGsu7NehDaFSnEaoCn6vTATd8vkvmNUVanOIFldQ1+0I+1n08QMnh9QECbxE7/0
Uzu7JxSIpcv81fkrfIKdwGhSIYWXxTIgaihsOa9C9+y5Vv3EhG55GpE6bFqa3r5Hc2cwb9HOJN4p
d5GPuzCHJc7JZ+8//4a2iOg3m7353QeoyYYJP/jHwcPLX2/B5c9InieFsncneLLe5CbjYJxbcBZg
qfiPDWmN1lMboxcBXI0c8hCTfpAUz3KYt3VA6Ov7TA0RDsQve20kMuiQZNDWmITFNM3L6k6iSPhc
cNLlvsDhnkV3wtdeyDX8Oqbd7wRrii5iV5hWatHyPRqyLMLTraOt4ZOi3TNIxMMT3EfvxzfcpF5k
zr7W7rSfbnTirg1jOEsy2ETxJl4em8NSPrmkTetuLOz05cQldO0xg+1p0E1vn/D/20gs1xKywsn1
gdfwqJXgsCpBfbq8vBDjqY/N15xCsG+U09Wh5Mh78VREThpnTJOHslALkUxQOw6glfuqRTKmxcWz
j824b3H4OIdeZoRNqp8IQCwefB0Wqg+FXYqW3vb+ZRvxvb4X+zFnthYX5PBM29KCsQm/yQQOOPMu
Gfl32mYJnVKn7H0Sda3Lexd72SxUY0WH1VbqUcR6GSEXxm8uTkdgpnB+eXi404jqrl4EreUqcBXY
RjOuabgmsPVbf/J2Ed16VRdNCsO3EzxOsQGxIg7Cw3yhA9xsD137bu1qsRVFx03tvVnlgxlGdPy0
C56+Ky1Ctx3kpRWeHw1TCYDs/kXloFIN2EexOONVW+rjDPysioGtS4Pi5N05UcBtyG7YYEYr1sD0
hVtOn4sDqCOLOFWZAJxqIGmbruISWQAFkO8CDTqYgo79hk/PZlTymt3RLiE4bZ/Vipj8P+dV9cH6
W2a/+OJrA3V8OpcyLfHTBpsMZ7X/4itagmM6l/lzgz7lHkZkf7r01PPBsFT5ZjklJMkwdOlduoTA
We32CfiEX8mf/bz2AONY5MjZrgncq4TbdEJmxUzg8ut6wvcM2U44H+EUt5khY4u+6F1nA+pLsEiW
gWiIGD0sInVU1slbE7m7HE8g+smHrim4KlJu1qD9sEqFdNB/jHIVbkiA8mQAUsIsCkzMqHihAdYw
cidoc7jFt7RsHAp74gwAIhi8laKhXa1WXZWRKHuHtzRuQIIcQo7cMtE6u+zLcGaB+6M2EyV5Zomj
UIVDW/Y5s88iT/DW3TMxoqw9PoIDqDXdIyjNTPZgjXTCUa1WnCrmcrIxufsS8NrOppI8cJZrsNDe
2jHM6VnTeuTDU5pjzGCaB31A21MNxm8tWH2G1Taz+0BGRfAsoJ85caikYvnKmRzFhx7FMotxuGVd
tUeRLSCe/WXdYcBPEzTXxOKT7ZYbPu7ezXO+Gx6ATFoYuOHfRkcnXHl4O2Y8UgWOzi9bRQbJQop7
GivPi6PV6cl+ahSMhd/tfxyZFut7HzoIbJTQz/ZDPOQ0lO/ufLPuNSJeGyT4necFxOhLtBQzP5XK
geMRdg66ceRXFbdvsm1yPdUKHIv12eK/jYMjtl0jKRk1VtgRHEeoNXUfBiEcN0UpOl6LGT701vVu
i6bRoHqgee1egEedK7cz+HIxdr6VPBnQGkyNwn4QyEhNF6RKyyM+Qv+8H55oJSQQ49Oq3Lbo7jwU
E0Pd1c3sKiPceObfkP3Prt+nQbad5kiuNfhmgdVMHcSmrZRP6loKI8+Akhf+ac1aB9FUACg/SveQ
QTaOjpICn9Oi0Y9IfGKpdB/3mbS3swAY1UXAFf9lmoqr5+U6zE3ctHfM5XggN5SI/HldmC3L/luT
rBwO+STqdpBWBkcOlQKXF6b22SuKEtKCn2SESmgHb5FQ6P48iuZRnumgJ1jLbTFV1kKkynsG4ljg
zM56k3R/hNfaOJk3NBFf0hMC8EiA7cS2lwzDP0RTkF3Bh3ZQb8ORQuKV30Ns7VpUuvTVliwNn6rs
izdcZgL38T4GEUEvBPu23D2qeZNjCbeHt/Apz9ZnO4pl0M/WlKZeTSpwqB+Vh1Blq5RlGWjgrrHv
HWHlXFYX1d372pUAuF9K5tQ3em5asYmq/nXKac7dFetq1xprtBVCXh3znGVkdcW9yzcrdPEwKo9n
o7Qi6LLzI8AiL7OQrt7t+HK3TOQA/kU4OTtyzoemf0BbKzbbGYPKkNAr+GejQGOdYppfi320s2K1
XG/RatWU6IdBHu8w2IEMwiUAI4wkglUsC/U4hsp7Yt4vpx0ikXUyoqCcP2k+zHulzHfHg4uOAV5R
XprDBJ4xlLebPyl2La/9MIIVv038IQmsXYf+gJtcOeNxnTEQqmopZ12hpe00wHG0UVoZCkBgUSSi
zkyabCHiIE6Yheey/yuCFLUiSKhQ60nezmWpKwj4Pw0dt9aTUtT5UlmeEw1q94/gzoV2Wn5ncrpu
Y2BfN78hu8g9BExOu6xSVlqXcOYMJ4LDoJmDiFUf+zU1rAgpnIo9V+kdn9GIQZD3k5yprjWI/47w
G2dFHeZHHeR6EcRUm/7UErtw6IQXH/GFZNZow8VgjSxN132u58IiAfaxqwl0nFyTPHanuMJoxVYQ
+YcrvzpxWP4TmaxR+jMy+fENC2kBqT+Jh+PVuR80fRj/3Jkfh1CkGiYMY5onm8Amp5e4JAvamONP
vdsCMOShXcVaoqMk2itiAo9okuZlX1KR1jZhKntyU0qX6wIUPgrlm6kFmazhyhVQL4Dw3vFEpeis
tMuBH0gKowOem+1YVkmSgak4gqhnLb+xPG8Lm6DSqgJvSBrK/CTsfxuTSyWJGi7atE0TANKAGDEL
u64Y9zZ9Iwfz3z5igIUz05TiMIgvJrRnmpU+MTtTdN5klmpf9vNyEBd+ZZs0OTR+j3Z3ohcuFeBM
+Q+OSwy27fBmyJeeHBs9XztuYcx48nDYNe+zpFHPSlbLDMr68uMaSSpoAwcV9mhv6G2crc231aa7
CHrTnS+Q05pZv31iKF2jcmjI13ECyEGdFb6Th0FpYbirQVSeZP0FK7O+VatH6alLzqz9FmYAeeAm
NoBybVhPWncUBRUZsUe5VmC8jIDXIjz4gpxj295SRvogw6zc8n8FBQVjdJzJ73fEJTuQ6xMdk0g7
1+bcHT9hpKByzoSEOPQ1bJQPd6NZzYUdiK0XypGT9HIRpQneFNBNNNEwAAOJOxPlMsRw0bYYOYq4
s7kD04w/S5OFNxCyMAn4H0467U9n8SLo4cSLsSxLQK7PqAD+lCW0sGKWHseBx9FFFIaEOs8djRaa
MpUEaooevlHO+R6zclRAAKoW7y50rUh1qOoWOh3NMzdNY6z6sMb7z4xTIET5cUfNU6HKbP75F7dZ
jSWLgpB2PJEoABhmnoBSqTH8PPjIGdMOR02pv5I4nySakaj8d/0iVhDwPpX6KGRCrx0z/l8HEFdS
7cQRfKGLrMrWhUb8k4vbjWpLPamNuhylmxVdDZIzx3CYtGGCqr1Vt/Ee/xrfwWW/HAidHL8rxL1d
Wz8Ly0gyMgq/SeiVwcFlYugKNdD0iymYZfYeXC/ZnBpprJYl5nPXLMJrSvD4macKCHtjUFSp8o9q
JVDwPvReAADZbnHsob2RFJlekFiKN18QABdGyUWh/AXTCvCjRGTnZfouuCBxHnHo6IqitLyNVe8N
RONmBlTGXqWQG3gVoUGjiWudVtq92O2Ft3zm+T3IPCc0dBQPJXhueYcGXbdELucIOdIYoB/Jxs1B
5QcAuCZZwUdiob8Slliofa3D+w3e7dfMTzKe7utuaFNCmw8VwfWiNyBgFHm8eEPQRqLqsrpH5AT+
4/7NC1/w0wnn8BI0rQSTsULoppnGIu9dpt7Zcx8nxGDBUq8LtxBzgFfCaLaGxGJ7N7NnTa7JkIyI
MoiNdJcutHlp0PR2XYBQ/uZNs5IUUC9lsLiMVm6xCpip0KcrTt9H06eQErmapwXBd3tHnH/DVld2
p/cRcrSnuYH3uoPY0QBmXjRMlvo6hcN/xdZpRxJL82SHvP7kaRq49LnQFjEjEum2R4iV01+hUp0s
XI5X5gp4PQbto3sTwpkW2nKj5nxxC5BQoiCQpj4K2F++9DHLSNJOSdGSHXY+EFNw7NaqnkoPTRnX
KFaTTnEIOjt63NJZMJ0YMQBtfOT+tbbg8nFLiu5G8SqikzNJsfPfYMw/NwYahhu6IXal42QRwuj+
7Aw/G/86E0RKSrs/sjn82C3l+aXdB0b6QoU7lV1zse3lbwEVjEdR0lKpyDhUNLlG3tjydgOnll6F
yG+gMog1gMoKwM9f8PfdVOj3AYZsxl3i3NIBTIxM73CTYuhKtqZZdPYw9neRMduT0jRI9J0cQBzc
TZuFsyF/nC0TqdSyrrzd5E9ZyBIzwn3gtUYv2QDopsaBClVj8RvXwKhrv56a26r8ThIeu2mkiKUz
8VuCPT7oCChXHDRh6nQRJUJnwIvcYO1/v0E/0+urAsfKjNnz81PXvlikwdDwDKhrK1FuUeCoFOUx
dINEqVPEM1vTqYXZRo51glTf9GnSR0Mbt7Xy3gLhAF/tMtmLf5TH5gEqjVTmbowV0MVme3NZ5Zlg
FOAjZhn597ZNrqNj5P1v7WYNk4vP14FGEe5LqT0dVSsjClsfzIqfDbGN+1qT84c0GByFan6VY1FE
/Y3xxsG6owCWv3H8J+CjPGex4aVulUaTr7AyZ1t0o73xrki7zTj6p/o5Df9b6zrsowOnBuERdN1x
JZM7xyVMIgNLLpWggF+gz9tGSJ1ryfWWfChWU1UG8sR0BBPtO4C99brRb4mEw3Apo9Ct7Bi/hvS/
QqjHc4Lt75HCgPzOSZ5FO0Z1c9NDOv0QFkaKDUuz9aprVVL84Q/VqLjla/LRUjUahouJ9JDP9DLb
6wBUgUB2DeDwi5iDAEQzxmP19QcFjuSauaexUYJGUt2nf6lz356f6HVSEAPwtAugbrYVLWQ8FHua
Cjxo52y5Aw3n07NDmsOzMX1XuD5Gy7mxRGBV+1JoobwoSnUNMiOkJpRy3N9ge6fWuiRQoLz3dqp3
KrkGobtUhPxY1LhHV5pJcvQP1lAol/oLnAuaGms1p1EV8ygV/TrU//RxQodv3ifH6NQkbNxq8ksW
10JDoFLsBVMU9DQvphDZttTbP/2tb0Igp9zW1bhM4w10NaLIe3KnPpLfyzJWlB2gEahXrjIpR08T
ryGZZ9JZWO075yPTlE4XB8SErSwm/ts7pXOJ949DCHY4Lzo3Im+Qn0TWRzXH0hjtVKAJGDrjF3nZ
zRAyldsta2biL7h+wxoWevx49M4grBcFjAv0mXou7Pv4QwjxURVCRe5AxIbWp144iKw79jgJ8DqL
wJKD/EF+BwUTZV9/IJMaC3OZp3zAS+8LbEHher+kGfjSfxgWIemHbChzv+F/lg/fpv3URS+PlG76
eqSJOc5aNjIkHtLcnVu6THlV8792aOhUR/JsZsPCa23SgSfluVgu3KARUcwehCmjTpXggLuz/Aet
OAnW4hP7F13g2VLy5mebC34mUv6ELp1Tv/zJa99QWCPCjaZZL1HcT50tsNJYBj14RqzOmiasGHf3
EG1PYbc17LeIlw644MDIRM56uMLTLS10kS79o/aoVpWhr56VP8VWPRrfF+e8mI8UdL9pP27HNFpb
p9D1OaX6vwgWRR1WbD2AIVCZmKMG6FyBljHRT+/s+YtLr5oAx5JRBeBBzLr25wXmSfRQ/ylXLRHC
CXwb3sHighU11QSaisYkSqtoWCclODs2eZN67y1ORqKJMBI00b7O/6bn4m3NzMo+ho8d+GIAClb+
nf9GHkJRQbyK5gg8rQqs3oS31rlEPgBjRK/FqV2JHK6r4KNpiaY7kTpo0FuZSW3avHs/236I4Jwp
nFclrp42UfEYQ5EYINtHti1QPDSm+I0H+HqFqmLAMP4l4j5yTvpfsroKARVY9COSf2z5+OR//JBH
Yzy36sEPdMraJsSpBnblZIPCYVVqCaHaRk6ecAEFrV2ncGdRVrVr9zpLgpMVhZ+QLHfhGt/Pnxwg
rS54uZ9kqN8KMEzDgiaZoBlgHSdhDjTvsmfeOG08vBDTlaqTL05m38lrl5Bv7TP4TL/iPSxGjMDv
4BIDdkYlV/Wgq+AFbK55SvOegA+z6yZOrHS3N2JijU3nEiSzwhc2PArNn5XkEyeogCPDc/HKOgIL
0luUOpZCQR1PA3uLEkUNOdB1EsZr4zy1SPxz+eOKmVWXqdqO2GZZQLa6xYi7tshIYrAgocWUhYbZ
xFWmxp2gMXT7QWgjWQsZ5V7FIy/VddDnxIkSOTbSzclPMZKea6ZW7N/SYiPyMwR4aArVOFJbilzw
DEREFWMHk5D2gZWDVbxS+Z/dbjeJPvZlbRVTsasy9tj/fkNpYdLgtWp3Q6j1suufEk0KXZWbgu7B
WiiU+cOEN+G487bl3O24WdSYVfQIEBcZiGSvH+dD6Iy/wrbqe0uDK1R+k2FK34C16TJe9hCNqwKE
F9B54gouViZ1WrrL6dHQCiUAL59lSnDkN/yVWTvoHGgHy4i8c83kAlQfPs2vEok9N36Q5cR/5ZpT
kB4WR7Dfts0CwS+rWaswqO3dv+u5ry7VIqirhEsAQFSWumuy4k5VVEjaE1BbTE4WhUjh6zCWjjY5
Lsj71c5R6CegdOOoIszIe76f3OcMabiCrtksbU+2iaZ6kUSGWObyi2FMOrwHrKpgGWYelGqK4dxq
R0RrHObDpEXTyx5VA8DajItx8cadtlE+i/7PFpUTjjzGqQr0LKmoH3k96tRv3KCy8IVlXeLoLozk
X/7dCq7nLGrRnuiNWHXDCwwhkF5BgPuEO02U7WcorZFMERTqj/Gm2hD110mf6+fygsW6kGADEuUl
ONTe3VpDdQV8KXnvSVcZpLNfxv7g6fY3DMds4UQ7hRGRxS/My7T008s0XKzXUKrANu3KnMNzcO0T
RxYTlBMcsYWwUliXN6qoO3RCRtUs/RrsLkIdsZPppwZ+cgXLxFDW5R5UegVzsbN4dLt5a71LxFVo
4TOyOxqPfFoGWjGwSvJYp17haI34kARa4exnUkxo/DK2A1tvK+oXPUp+dDhIm0wAVKml0rrEZmPE
BtE7n5Ii9+FK1PDxH37HnQjDlwvSCr4q3/vNwZ06d87e58gpy1Z/ymJnntG9ge2cCaSLtiwZx8J2
G0X9hQCp51kee/gHy+1JMmkkO1qZMy1z/zsCgGh1WVWDn3JmX/g2CXqnH5AP8C5kLDSmCBYq0/73
yp9tUQLNUJyWtKphefswJSaEBUzLYd3Gb9rpGfMlpLklB4jBHi8pNuHmEbG1b8Q2YGw5ZiO9FLuK
YpeV+CkHWUm7RsDKwygFwDl3Nj3xaC7WWAt6yYwTKpxP1/t2QT9M3lMK3E+rvZ6/068OJCNNhbDl
g2Jvw7tGZg5CVnyeBBlTqgyU0nbkz/rr8nc6/8h0Rz/4QvC6WVNgiFLFDb7p70hYDtcX8xw8qqEp
NC1l7soK9SPwNJxUw5eLLZbWX8wOPlcRlKqzNH/L+XlkBByQt+UoARTTqWrk2GK24T3OYU6XiD8j
xAR8pV7i1V21feK9Nd3iv/IQ81t2V3GjwccnRBaNZizLUYsJ2ME5952Azy1eXFCdZslBpBb/fYMn
+IIeIbkbn+G378JrXnQaZjyMnxeCJ76PLOn3NtnPxoYjXm2kmX5q9WytrcILqBcSjfug6c6z9X4z
E9rugu9/FHsT/tArn1FIL1PTbXJllpXYX6b+s2d4oDd0mkQCORpmMQ4WkJkAJZJdAUf0m10TboFY
FSiK2fLtaA2Yt2BpxnOQ2JeE8XUOwf2paZu9KtfQhxomLsgxqJGnE1bOiPkQz2gj9lIryf16VGJZ
UwGrLtjJ5inlXbpmSZC6zq1TJ4Egagh4jHEZ8z/UCvihns9t92uNyRDeEhx3cCQXCHg50tpEnI3n
lqQJJwbLyYR7ClqrSbyJUi/NrISbBiVRGZw0V2i5Mv6myTelt3O5UEdgRB39oo0im8CN3pTkf8Fh
ysSzJnW40rsSatyc+z73o1efoaY2l4gGb+wesqgI17gq0qSrdIC3YM0BSJ89JAc/cvxmkI1RmRLO
B1M8IhQD/y4X8wlap5HtgMWdsIG/2ZY/lbN/8lxqHUAma1PuPo15IbOOkn84h3Lm23SDAEJIX4i8
xU+1MB+XeImmrmnDDACL5KgcvxrVoW4EVDDnwXh7AA+zQeRiQ+3eh1BzLY/7XqSArVeDB9yHhq95
217wbTZrx3nhc5bmxXtazdPe++ff7sjS9BBzgORXfwwrIchI9crFiJLQe4leuxOQZoxhzhfwdU/5
G5b4/UifUr5SBpLFIMbh2Avn8Iz3/2qclxPukwXzMRrLYCWgkRzHIAR4rpSAf6k3asb5TH1IDq18
xJEvFQcCSqNBwBKE+93wUdBqRoH4Jzvul/VPoOKD4j6IXz9SRt1tdMSXhvoPjmpI+ZL7vd9jFHw+
mpKPVQbpNgtvIOnwjVurfuviWaeOXPqrESTgmHnKKbUyX5j0GCa4YGY3QOgHq32+dtYspCOzJEav
GDasO/VgSMA07SyPy8TPttt629t0dPbO9Enl9rqKeutn9S+AZ1G0r/d6G+gJL4NbtWKk2Yxj39+i
SibqjVmmQ6KqLBrW0ieHBxV7F1HMG6AfarehGWUrxkv/HQkmR3qSS7kbec3AYr4w30Tk6//Ah+DW
WT84OA0MM4WSNtnHc1KlQ3dbdONlH++CrOWIo5wunJrcBkMWZlCmZ/G0b+RPyVOutiDW5z/FFBV/
LvrllcgvB0+2BeQcL/Mr5DtVkH3cmAQSsNW8InHwLTUjJLno5b003C2xzbB4uQSoL2ZVJDPkeVuX
XpwHTLwagx4F528pKUMWXdqgEBJmiH9L0/z5JxLJ6ibLQO2iYtAZ1Ov7Xl/q3J7sOS6BZ8R3xycT
N3oQMGgqcx4BC0h07rwkTtcJILG+565c+1sTQZN0gu5sfkEQtPFpDi0PKBmDMdcaCnpGF4glMaN+
Q02mSTtnhFjCachDrQzh+ke0NdRiFcwwf+7B7nVwwUXcayXnEtOQhGsKmH5D+eaqE2gfDwOdC1/9
TQ2vy6ibpu9r6D3UUxgAE7vE9W0sfOz2aYTUgXfUZXgFQlIzGaAy8W/QQnsMEM52kPxIptlf5TyU
f28bdKMwXNK28g+95HC5elBOKShROIhpNou6iHlf9MiEoXcPBuZz29+b6rsDHZFAF6bzse5oaXtf
saQgfUCOn1eQp7KmHEgteNP828CeEl6vdwhCfiUVKr+VaiQGs/BDvJS0wQ+srF1LqLG239xLQmIz
StzElwDzHSPg58a7qSHEG03adu5mnRcggsAKbGZcK0+F8b1wHjj41ffHEsCUJNL1FXQM/yzScFc7
JeZVSNVJahVqWh786/KJQ4Zt/w63wnxJoF5TtyBjhcYiSQ5lLHw0ScpAP52ROJgzyN3siB3z7UQu
q42tjGi9rA8uCCDpUDhLegT0X8zS1t6OrWXKo1lzwO2Mr+MZHi2Yd+a27VssCcA4zSXR1jJrfhZj
D7JTLmafQuv+xIOAoCHERHIoXcZc48fZ/vRHbp9EWEMXl2imNkdGMHtD4nIx6QEAGUyINCh3YYIf
dmH9AoOKkWzFoBLQXa30+ziaUQXQXJiQ4F93Bg5yFqsBNQoQlzPamF7momi+0MWhulmgCBwPkpvY
3EDviE1DMhj3gMuBVy+3Yac027BEp+doohvl0HHQzsdeWty1MBbYk/jQ5GnxgspXdMPKGabQbhN6
dm2hSaiPx3AsKGQz8eF0XQ0g/lVhWxH37o0bkxjDP9tjx00TCR8ElN9xuWrnuQ27RUsuT7dHXZKG
sZtILi1gzXqtRyso0ZOJkPHnzD+eQFH8OLspYhxP1XQl1XffcSIZwSSUl7ThvvC8zZdyK+RuBYyP
De02DO/RXcj7EfpBkTp8gyPElMze8cvG+PnHAeLgIbvZZ9jx/Hcxe5dk0w7c1Wu1d0v6ctfsudrO
wwZaMh7wC8OsHFSzNS0CTypoG3cbtysj2g2oirr2jMubbU7blDlTWJBn0nUj340Kmo1NPO8ErVPW
9piT1YY0fS13RiwtvESyfKfrZk4X/F7Cmn8yv2mFjzO5mbpkoPu/bMHhJ+8lqC03dg1Qc3g9dxlX
fh6oBfx+3nuweZi885L1Kk4uUIwON+Zeec3fzA5p2xG5G/quTATSoCX4YwvO55BnLwOfMMpKgMF6
NG9m8w5PDama3YMk/VpKTKH9gckWI/692pZxmLngpCqFEAtc56hmr/U4C4V8jVVG8RP8leoTGMaB
UJNt/ezWRnhOdFk9950kh6KiOu0I5Yxipr+uS0zjDqK8QkAtLOdMNeyI+uXXjl9BcvkJiRCqQgn2
k0AzFe9U+AIVbXqkXGE2sqKFPTwiuIuZTwKTkgyUHjwWMhoWrSOu65iC2v2RY46CIvnu/QaPNXN9
a3V+7uRRC88dymJL8PTXOjC3E61FZn3+jP1vJvjIXuYsMQcrH0zzuPuUYnMP05lH9V0716k+52U2
VETP7zY7SVth8UISVIQUOBsVslbJOiXtfGN0U+xO805j2M6kdgMmBv2hL7GKEVs1qpgvy8wmJ5c6
3FhYMagB5MH9j/6T+fIQEw6oYmZUG02Ma9z+XPgPthyvOlb1IPcYyiRv5tcVUn0yWKhzxZGUioVU
lJcEDYwWMaD6BEZeppJB2rXsC3FaFAiKpC9QxFexe/kjKVnMwMDjStPb8VUOS6Aat3twr5EUtm/8
/zXvKlOK9gB0wsLxjMcaaWdf5FJAnZV0Uw4FTVPq7edEC06XLLW52w5iwX0WdLwA32K/gKkZ4aHh
fxbupOn3RheUzmWL5scRkh2l43U7qC8BaLMHStJSMkpqJ5uP/VYBwI14YylMnpz/XpQkaD09leJY
HXslqVLdvdah+rFTJEqNSDlAiJiBKK9C4p6cKKm6QplKOoJIsfD9UX8D+G+3f2DQgsniEY9xUNEU
98e981NBJvcT6exZDSjOfOzdLuPXFwwPG6kALFU8TVZ5Jgsa9MgD/S2i3Ov7ydWdNNUqgl9x3bN3
FdsCaBp+FNnCFVqHr98vHDH7qcgtLPKSFFQvU/Iev7HVw3HDXXCOUw1xvUvdF+wETOKwPSaCtSfc
O7ocy/SXaVpQ1TJQq3YGN5XpnLD+4EIQJ+4UyC+QA2vD6bW7aUUYUxYDw9WEfJAHlK5V5ym9l8ZH
cKyv6V9zugcW/JbiL7B3P49peex5JSTlpBbmAX931A0kNtSzFYVBm2QDEOyBVWFo/QI1OKhSbF0K
OhngR1JDkaRY9VRtMpMld+F4SyZjtlc64d3C6iIJlVOLF8PXiOAjj2gMx/l5pWu5ea/wCJV38J/E
cuOzVzmBgcx1hw0jyFnXYYdhBLfPxoTWaK8E/JPajTc9keK0L3Z84vaN2u0WsxG3B4jKhUBYaUNO
1It8mtOEPI8iHR3T79W9nxaul+Fd5ws1QRnGYYTPxije+l35JFX6XjGzulXuLFjuLGBioS4dYBW/
Hy88VyQwTUj6GeLddB4tUcPQFKKN/gh2jnSxiiPQfoaDQX3yCUt7tRGqAxxURlTp61MvkCfTNbne
yvpm8dpseibLbCA9GYhDu9lsnH6+GpWHrz41qgEi2FqDo6lAfAhvIZE1Acx9g9t2UUSEc3VQUlqU
IwJUbXQEPh3g2GbTMPUawuPe4HEIVwDdHP3A5KYS4mdVoShUsjTlTlKcTn0wzMOHpSzL1IphJ9l3
34ywycF4qfeVgaMLy5e2T+Lj+aZFwyxzx3FYg/ivx6k8oXPbmDPjsgaf2cx770RXdue/oR4SbeJ5
R2sdQLb98CpyjX2ueJeSvdNbZR6QqZxCZKYLvpcJDchcbhMhogrUABBf5SKsAJqOLl3Pwyc+um2K
YUtHtWN9yPuPPceJhJD7kNfMF2rqbN7BIozeSteMLJTVPr0B8zRCEcNydg/6iudHOMSR6hdly8Pj
imeCjfnJvOcq3DS7xD16h4QaCREBNudw3OsYD6eML6nqQySIaKejFDOjWSpo/CkE5PcqbGxxVFzI
uHvMEA8I/gFvEj1yWQSBfCcgySI+ci725/Lfd3U2ghmb9Kzq2BKmot5xmPPFe1gPHkxPOfcJexMx
rTRiV29FjYkQsmvqKAHZGwUH+a83wtSKP4hPKVbFnxNrJu9wmdklGEdKiDHff88jtwRvDDucM7ri
Y+rHg1bdlPT85CJK1ZdGgeRqXka/5BXs/hPksQc+09Mrjh8rWAF4cZUI5t/fVzfKMtq/RqqSiFEq
1RS1L27oRCGtPxoC2HtNhLJGTGr5BadbiJsQKeMjfPPPzlh4GWw7mdo6JXXwhu4dVtDlzbFfyjxd
x1aH4xwmX73kwhfBiCmW1K+yKgN0UxgfLW/b+rPRf6NFI4d+R5JifFzMZRwyqv4PDSMbfvOntivk
6manHqkGLGNa7jWQhqT60+vStapeLH3t0bBTbgJOpx1RCRJIZR2VAhZcMjkRYnnYAMjdwSChoAR1
AVAmYzkyAk8KneQ5pxf9MNXn46DaNLZRzAIuFppctQfIKZk+z2XqF7IXppm4CxREz5IJe5pHDXfM
l6Jg5QCK2cR/6pUjR3qOYhQMrPt3LWd5bcdMCy0Xdh3IuxvYOiccL4acP4OOZhcVucqFMTYozyD2
9WNPxPdOki/s7gNP6OGBjxqg4/LpR+oT4Q4MkBDbQke4I3t5iifve57D+EoUq5O4Nd4idb82YQCM
gsJ5817jH1p3BRwvgtuTze7ASKPn41PrF/UVV2yALVK+hHyZqhorA78ZFHVU4aCh0Hi2AmSkSmjn
Y09q4dJbBC7XNdQIsW5VVgjPWfy3D8p8y85LpS7XnufC1GhvSwtOaaM0P6YHLSCxPBR/OzeYsJ95
pmDV7z4vNFh0X5Qr42k1kUxghyyC489TrFHgKSMTZaSj07wg1sXAKcyyqOjnikVhto5XPZFmZaBH
5oizFAbAjQqh4c2e6wC3UQWUab8nENZmH2NXBb0iacjOfJ9jtTXvxZxUyLm1JOzEhyxvkVn2uBFJ
ZnGzyIdDNo48fRZ6knQMgXiGud9ilDgcorIGVr69v+gwu60BdeVstHUzsOyaVuEwVb+wzuNoK9wG
7zvziBR6xcl1ZYvUp8zl1EIhKv/ncmhDSlC9cPpPe8nJhN2jygWc86zu+kTDtJeUXHpNu51E9TT4
liPJbz8VvSJLVqrqwltd53z6Zbk/zgI0MATdc/wOpbH0tQIR1l/uc3OWnKeBP2pI4dcnX2/NVbZH
zgVoVqQECQ8hwz/NmRmCh5fQOfHyjKCLejLnVT72rjB2XABALFHDi2Q5lJotBuQH/xKNLsoP3dck
pv2EgMcPXK16l5YjgzKgT4A0IgebQidxNICMfWCWVqfqumrNX5EvmVpaXtdkFidSoSPOsxWKXe28
2P9KsuMvbcoY/G5MnzBYJFfwyoxHo6wQEGGSCrTw3ja6WQRrgqDRR7VJQoN2e4VvZSk+iHsmYpkd
cjyInFGcc6wLOGIWhFgDWfDCt7Qa1tKV5VtJKyi0Ai+IHJCi+vBuNZG2ReC8PnQkDzN+SvoStN3q
cxyuI6txZK1a5bsXk/y9c525KyEwiYRVIKcNiT+3x9rKSK3U280OYGY0z/YEjqksqeQYhH+lMZQP
yxXwGm4Jdu3sDicT19o2DB2lylgf84/wq4q0ERrDx1S7tfuEu6dCyQkKnuqAIUZnaDih9diMHhMk
5OVj0YEuv4aJ6HUnj9G9gnPu6wP/XFaS4GiJmbWr7ykFx+Yy45vJZ/5PBVduZSyrO+B765q1/Ztg
i9f0qwHtRu6GJr7+Sz3TYn812UWZmWXSgqxj22Cfj2BITtvUFiUtraRhUzkGPWaqzuHvS3z+TPsp
r4pmQGKaOAYrpsZxIfdarpyoTvoGRBASVDGLhbHuBUtio+SYM9WjvDSL9d6j87rz38PzcGXbaE4s
GCG71A7C8OG2A4Xi+Vf7cbRBwj2XvWvdzuYNh1yCxJ/Ct+UMxU8CaFE++LcbMJht7YPBvDRsQkwX
F4JpozxCtIjQu9G+nWt3O/0Htws5ELMtkXOwg3pIK1ctSEKCPuAQi27t2kDJSmSwEc4OW/rz+WWN
EpH010BGvxmRsY6R3d0sse5YRdFQefEEfwjU57PnBjvplJ/CdEqVa+21en1IS1nZFIDg9EVEB/l0
pGM5oM6BR6s94r9Tt5HgEeWk5YXwt3iqeZd+X7ewCIsDFn56O1mKx04ePLLLhSb0LbqdXk+bRXo8
R4WvGE3316eTL521Xun3d+GGQ2QAfVFmNe0gZbm48YWEpIKzU/z9OnjUKheUJskzUug+HsmhOhQa
TXB3EdR8aj8fsHLDSy87jyWzdm6vFwc74UsKXUuMlhSsalcUiGpL3b4c1XQ8PXuD/O3CLdoQ7raV
hEpJLlfxL71siHDVv9G0sq18I9sXCHk+a1S6jW/ydHR840TdoKFDSe7ezHm2oBI8g2qnbFIkjPwA
LiD4hK9GF+x3jVkcEie3fjgVEtoH4eF6MnEybg6bvJmq6e2oDvZV+YPO4+Xo1hPEVe8ajuiH2Rwu
F08SxyA/1x53i0zERABxgajUehzfcAgVIgeJCwUJBA/htMZtfcwM7RTTMinumL6Y/lqAW+mQizyj
ee4/H+6zcZ5pkBJtp+VOc8DJCVTOiUi3jZuShJ3U03EZbArASSaHfJqG92emVYoq6W6w28c4GhPU
Tu4SHDl7Dzof4mE4AMyM+tg2HomVq1qWhiuSgYDP0NVfG7FRoJ2lMJYbkQzY7CVbIxy3Spxr3zzG
miSRwe9aWFH942uU3IizyLAL+fVfKCeTGm7xNVu7+r2b8qx4HHTfB2BXjocKapmEXeDXlVjLocrQ
3Hbj27gYC9uqcE/DH1eVBhGxe0yiOE8R+1nulZWDbhmFqKl9oRIYC5EBtJMgtLc74fUUN2vDxfJ5
n0RmroKbJm5hITa5ffrxJ21nsF5hSxIO24o4duaXZ70plMxfztZwWVcyAisdqfZwhA/T/k+1EFIX
EG4Jm0FttwakgsZ1DOHn0JLu3q3xhxqGgpy6YqFINrKykzJMkgEo5272kZl7YeEYSgp0hoSD0z6/
6f3Ds8LniJ9ihQSlU04nkv3ygYS/Mo6g0i7SpydhSJW4yqYA2cVZxxsIuNyjXEdotovKpr/zaeHX
NiPnDX0/C0xpGtU+QOfKLUQ4jVxn9DPKM1YVazAHnBSEA933I+7YR8uSvNbJdJ713rYIcQruLBUu
LiULFoYW0iZsqfUmQy0ywQ72neCmmfEeiUa8bLLzSiV7FCW7aL/r9FJQXqPc6cPEfdsZFRl7T2Wt
ErXN5WDjiZpCQkioNBFOfvzywu33+T+wxuOsSA1OLzxpDfdUt41cQZ6wxMSHNdEWXSJ7EE3XlGRf
Q6gD7Xlzx8Hc5dX5uzhhUNISae1Si15Kht9Jd1EOoz+vEOw968gih86qvw0tR1+cCGRX5IcYpNX3
cxBG0QaqzIc9Il+YwFOivcvaXvoYOHp0lWq0RwuQhE4V5rRoTByKhDkt5yP6DoZKKoPuTTqsR9TA
/4KHV2njXUE24kfKNc7ztjtzD6PlK3pvhWX9Y2owxuHHOvlmaHcF6LdIiwCmPg7PHtWEQuF8LOCG
ffMh0JhEr6AadXM9lpWAEOFn0GYVte//6RAKvTf6hn+BwoG02SRQeNyvFYpbwKljsnJFnNzPCJhg
kQp+YayXdntvE7V5fkkksf3/1+afjhEKonksKsJ7U6FtmaoJQVp9y3GiUMmnjva5xYq6Nw78V9or
XxIKUegtl5WtczRm5a021bXmr+05brDuA/Dq/wNAi9cwCc+LUzZQ/ghlkyYuTwbpkBfXyL1wthTv
/+Awo9LEWx7GONXfzfw8z2McV6sVdk5PdAiwpSk/+jRXWcdJb/lTNL4mS/d8vcq/5L1p8QP7BMhG
uStDyNM12R15bRf5kmWDRMl/vRZpGHgVX7VtFZ1RbezioOsn6kssOqcwdwKTriO6WHwaCqU0KmZX
UleadLGiPnHCGW5f8Ucu4R7/mPP764R0sZyP6MrM+pFZXwWkqGzv8BnoT+HPlICgUh1CJEXtdt8f
2yjcd3ACgGXGRcblsaWaTey9MS/YEa1ml3veUowRHjyffVUpZrD53WH5Z4qosgebpiBWmVFu2YWq
tRlBBw1QY1iabB3o0lwgI+ZvjyT1F1s27uQW0V+N+oSYrBYExd5+VhY/7SZbtoMR0kY9es5wdzjY
aryIUpUr56Klsfih1D6mg6L5tEUe2TS7+XhUSYUAF12m0+KjWJN52jQlQN/iGX6VN0pGIi2N447w
cG4RVeuQFIjZqaHJEO4PzTlyVh2M0KnXX2XI2ZAKVaYl/wn3ae5HkTm++Iu6Q6f1Yt3GzhrMdaVj
hasIOYJpWLxWyPnV4CPMabgJbgIHr4Lnw+PeM0k8Aa4Bc1kTm5EipOyAVyl3KlVKwExH8IGts9xa
stOjQQXZ/Yvoix6CbcmSziZy2sCWMMiIYU+mvtX7vKu68Aiqf+YLFMFrf48Jzwv80O7nSJHGf8z4
BLKd9SAt4dvWndx5nwlaox3ruLOVoZ8pz/TisYUgxq/SlsL+JJCDihERQ5vlUBi0V/ClAt444Hl0
xusjY9hi5P1XOlEkLBQUjX9JEEoHeP2Pr8aH7uANdDqFc8KIEJ5xoKKCIvHR4YrjrJ96dWE1Z+rR
QWuloCpzo2HRph/ULkl5M4DAABFefsRC0wqx4S1facFAXdBtylgKQojLYGRzjCk327s2Fl5w5K1N
/O6AnyGRRuQVWYqzHliOEb/Nq8LWbVIr0LJEC0Ge2GGQSYJNLX4Xeh/3RZZa5UyzalVEnLDqFbfr
5CYt0KLYM6syuFraN8xqRxxGDBy0ejm2MUEGpdlQ9r6J0AHJHQ+UvgYHMIav/Mw4irMsWcgoPM7K
rM8R+m7/OOUqb4RfgPY/IqxM66K5rfuXUdKbICXPh3MdX4BAO1xrrOJCYt+FweXRJEBaNvVL10gv
QtWXowpXqE0uxrEcBtnjrwm3K/UyPGseVJqmtl1RqmGHhT3dbnfjZsGXsj2qzRGYP6hccXxqywcf
idbA5jCr4KqmSVqkqoxCgDGUDL7M6RyZTovhXXRC/rz4nnqd9vSqJPH8t8pQLL9ZlJ6YJOqcxVH/
AUza1z5H9LNwvLfDOIsrSnO9i+zr1/dBn8aBwLZlUl5jPZGScJvcLdkZwqs4NVZKsEjv1bAJjZbe
sqhTYpm1EbnFeuPffX311pC0TDQlUblgxdeheOCRXSmz0ixzkFfTp7HhxTocd+ci9LkUTySKWpTI
QnCmjBltZ15yqRfUx6Edqo0LwobgCfuOC3FDO3mHU7f4vTKBjqChiYBpVuI3DsqqB8xIy/CWA5Vg
JjAtpcjPLekgTlFNMqY/6JCeBgc4ltMAmfI5yieT1y1qJPtsssrh5DUPASd4eo0q8eeR4mlmSyPb
mvnep/d0vSl5Hzt6VZSCOcs7ZD5zBSazBRZgvdnwrFCxB8S+8FzhC1QftyzrXDjoRcswzsJKF5n8
E4kHmYdBcR7srbX3gkbH8JLR2r/KK3aLNa4ivjI1A6UCtnQ5bGkSaLHLjcRjP/D9e983N+p2YNO2
A98rM8VRc4idcXc9yJOn3O18g4OsP+ZzY7Ir05NHnT7brLIKtej+O3972MyDbIqliy3RCXAvAoFC
dGlnDgTazQIYZbbGJoxNpMqRXXN0lXgORDybMpi68ywiOotxapEVDrjqSIdVssNLrAP8P0XL2/OK
WznpSTjrYOTStuM3CHcqWOZduusInpAG/zJGDDCu41TdoYwpxKDSDu+p1ox3sT4h7j1cvK5L7lV2
H0S9vacxVYTgPzXnKVFg1DImslJ7QNkxnUETpuiUHHHRULo9lht0slXUp+9+hUeXvNwratVrMLcr
e/CRJLkFxTH8Tgx0U05spuQ7xyp40e9Hfd+tHvncrWUfx+1w6vNqqVGA9HyDcT/2fBrGh0g7+4Nx
iZlxBnTj+EacWT69aQGkNGSmIXtpBmoE5RW4PxDnywxtTN2U2o+U2O7YtBE4h8UEhaoLTlZtWYwv
GcAlMBPzAx0SLGThVoXq8y780UXy/AeSQKm1NAsJqsFZm5G36lGhrPrCDvuHJsLOJBnZnpfkrv1B
spJkPY61qEFz8+C4mgfYF+cTuNg6J6XUHA8qyVN55MHL1+rw4ReAa75MDTFvr432PoNZzz5Dsk51
1teCE6LeaogGndoCBoiiAos9NG6LqSnyIPYVRm/IR7S86tKXj+4cpiJ11NofREcCc7/VfFwsqSEY
+HztFVX9Fso//CqhM3GL8JA+fzD+G4IkCnLWdctoDwAxyH901ZQY8gQqOMvs6NG4QQFvivkW8Mpw
3axWqVIR5hYsjCB9FvEOLpTQUdim9aXfQRqlx2PTSROjWKFOwTsHus1DuDjQKSxk18DdyK55jOAy
JxggQtby3b4+SOA6UeNJwJ1XmYou3iNw2bFseSJr+z64P4Me5zCL0Vf4slk5Efp9E1JG006lcrJd
3Xo2G7Z5FlM8Nwm7WmjvVRY0YGpHxwwhQD/QWOAXM0sgXlYJo3ehsoPxxDVHvsvSmRV8Vx99o5Dj
Hzm69cmQOSfkZw2mkp/PFhUXSGzeprwwA8vynCMHSHPhnVG1yNTEnvzZxN8j2l1HOpctxPaPJ+Du
WGWtqYf3K7WrZyw/XNSjwTy4ZijdofsK6r/7LyJQ3PkyGy3cSmoJ6/Bfn5DLvJQaa7smhbrWQllq
jGnLyf+H6mvfJ7sA/oCI7guk1nOErPwEH/mH4a0hpbuMaMbToKSqceI5hGQ4lg7eJslAqCMJrJ8f
p3wTIko+bivhUFZDgWSyEd1TTxCvd2HduRgmLL6NwAro0q+GpsGJj9siCJ8V5acSRtVSQUF74pNI
xuc4obPxwq09V/yfXuFlBz6z5rnaQ8WP9tatjn8j/ew8rLElB/aIbl8dYFptczIYnr5LfW8VAEjs
4CxekyD+oiiYHSCR893mvYwH8vYjVFdQVDkfJKWt0Y0SXyv50ZNjsQTWaJeTZHLzRvSZeR9cNNoa
r/KzzjpQo6BHwlVVXh520PQAo8lSwF+qszFGXpHMN0s0JrH5xJNrhV8086pG7cBromO/OBSoFujt
6TulZcMRPHEcbW1EHTTusNGol7PAFlCszPRpgdH4QJ1jkJQYLMK0YaC+dI6303Uc7v0kyKSdWlCM
kdw+pqp81/Lsim/2u3EroBMRMtuCuw6O96n1D/N/6GFTLvgIMKCn2iKI5r8bohGTWg6/uMIHSMGA
QJEwfUgK98F4LkucfYRxur1M7A1sVv7mgBqlvbSOQJz5WpM3T+ZiSULj1D1kxOFj099BqhrMD1fH
C+v7XKdEYIgoUp/L+XZrgSG0H2V10cDW881759O9ohA5oaRqZMjIUpXUTYp1girwNHp8s7s3khNP
HLaMl6H0s9KHqkqYOjFTD2V9S/hug1fGWbZ6rtprEOjaA4ypj8MHf1jXSqlUJe/3EhxoZJtdrxJx
RxffmvJbJYiPVft5NuRrxlpqx08t0yZNgeWhzt4wOCbPvP+rDptfSXdR+6gBd2XOMQLD6dVVAsQk
raPUIT6mBZHuuAld7eDnrkeWwdmDujRc+v2jiNjJMaTQN1pZn6UUhz8RJD8hpy4uvyB3CgnN5/AI
c1Izyiaz7P381sGNBMWJCSPc5p9wL1nZIwMHbCMMeUAHQBiAKOrPLlKO7L5JAhYAGwthO/b+UsZ6
Dh3Qbd4DntJdg44Xqs7iWJIWHAepcxS6l2bC8g1wt07yntGgcoklP8cero2/Q8VuyaroHcGi7R7d
G6zK8GT5egdMVPcHScupIm5PBonFcuLRGWX8wLVYa51SRfw7fIm/aEJWioAciryrFs9iYmBl6tCQ
i8C1devy+wk31HsOPA+RUu1LSWcCJw4ZkAJD6OzaUAbxgMb86KNahml66tKM0Lggb2lXmfVqwjQn
3vQlmVJu1aJWa33y/a2gSyBiz1wUUEq4cFzXynNSjmvjiHLMhjuRJQsQ98WxG5jzdIemEE2jB1pD
QZNg59y2/sgVSS2eGm0wSasPd9AMPC/eAIKYzXaCgIcj29BVJbMZ2QMDvSu3fOJHwtcdpq/Xziri
/k06XSRe1dJx5SQktejwZdk8u++/P+HasuS//haCVW8SSeq73u/V9RLRaQtNxCPTVgjybAYfUpnR
OVjBY2GLu3cHq/g7/85RiTxzs6Y27n0NN88AZCtJJ1x7zWha0qY/E2DeXgVfCBpHD98hjFsdB7cj
Vv1VUk5xZA96Q3QdFGJB4Jcw9NlW6+UjJzCGU5e3Mmo5tIDnn6C9FSDK8Q219BXFsqPFNwzLb4/L
WVRLE34dodI7/526w1/DJyuM6lpWs68CkQF/2PfZiS5aaTVME5WdGTds1tDlRSDEX8Os1ooOTVs9
okYdhZm9el0pYloBE0THWVNJxHPYCAc+cnhwop2z8oLNmFTG9TbjS2KPolzKoCdIFf2EG7RrSZNy
I/2WKv7qs3cGRj8E0lyO5eAu2bbhDmEPmtDmw0npv9p6WOGK75UFOoiGQsXopiAPIkl2LF63SeFz
7jCs92bwMnIwedspjyK7CUrQvtfmNcvzQiE64IbQXgldpebhujhaKVSGL05UHGnLW/zaBFHS9IZn
IRWj9Iyb9iNRof352rYdA6n/v2Bxv+L6KMt3pfU4cbJhZyiVEYJYxZ3roh4G+W5+W9ODdV6ACdg=
`pragma protect end_protected
