`timescale 1ns/10ps

module pps_generator #(

)(
    input wire clk,rst_n,en,
    output logic pps
);
    

endmodule