`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
GtonvLyRIHa0BG5ascvXN09MZ3qOiFCm0qhQWasCekdFVRCizFoeirO1cOSD3S/L7XBtqzCllo4q
Q7pZwE0bdQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NcAWItlcyJiW5iNdkc1sQhABTpjXqZkOrg1X+Tcfgn7grREOKMnmze0hKfPSK2fx03p+1DXa9nI9
aDMO4y3pcvrSQRCRWXgMFS2qba1ARCCZEOEfr1i6f6+Nx8FGN5X5I1YnoGroW/YZxqunrLG+EqYi
XcxUyjBIkX9CxLSivhQ=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LPH3S1XGG8M+74c5vorJTX4Jd0Q7p5hXR2nHLPyVATbLKyNyCj3u2979H/5+r0KMFY+Eci03CiNr
huLATC3oqO+Ri3s+z9ShUHH0kb+eyBSFWWv4Vz/y3dKeMo7xd/qiF6cFD/jwZmVC699OpPLFZ+//
+v9QSba8dbzt+SXEN/jt0+eliBPMdqYocom4RnNiRzWVLRpczdP8jPK0iZ0dswvulkciexDQ2OOo
AH7xVOxZOGncQh6Vnj6rFermvVKMjP+f3wo5tFO3kt6qIlYJvlMl4+beZEF1FvA7E6pKL2F1zinI
FTyZEqwMwZWW/ux/d9gBr39V6BUQmOQXaUku1w==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XhsVvFI9R4kEmwKEMm1/ve3kzL6X2enhhJxnoXVsTfGBwYA297bpytmIip5AhwFQisRjBoqJ0K8l
8Pn3j20/SKo4hFrQQGF0dNNW6natF+zLk6mmfJ9vN5kjz0dnY6GDFbN+3VxaI7EfmTameGip8Srg
gxxI126PbwVBsgU+CTpGeuVit895aMS8BmBuDurrl1wtMGtV+dEhJIRJc0Aq1Wrns6Y56i0yfgPm
51nrGVg0WniIJHCwCd1amAGBP8K+XEMqgFg7Ax6FDLMI9fkEMpr36t/NLdEvEWInQ+uThyiFxWQr
JKb25unvEuv/D0FeWrozh8XdjpoKLAw1GPNMVg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
W3obImnatzWtWQxjvGXfWFuKaXr5FfPdOSZAbNOW8Mwmo4wQnwYiA7HkLDXfdrmslndHMaUxH/ah
zQFKiuR+SbrPT7aIULBLqqh72i8AksoYWph5t+HS6djOrRH3vsKtdR3ywmgroEjQ2QUcAo6U9K34
zqxoj8P9N8GP6+jAQYo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
p5NJqyb9TdyH8yE0AGM2W7x67vL0sjxs/jTTPTMrKPRWFxxZNuqsL6RAPf/W7gzVERxAO3iFqJD+
UoyFnOxci4budxkwr1k61TSgdoxD0V3HQjFvRukqTPnveyj/ep+eTC4LGfMpV/TPdXASgmKbIegz
1MyLz2/mIQLVdf6YMINHpls+EKIpYMQZpwK/hPkYr3E3OOOvzvQxNC9VDhaDMvYytD0fGysZMNYl
wnQ2rJfehLe6ywYzM95pSaORaRL+1Yx2J5fIpMdmGCqTlIRPg/vBGdEvfU7LTH681IczR8haG53W
YAR00ATaZUq26o3QwofFA/jZlZZYcN6rMAOtfQ==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OsRx87MiUvQMyOGPSETijoG08vE4+CeK9YRUiBEhaa6o5uSa2mSyUldHexlwxMR1rBWiQ6uyqUCt
nOrLjKhAiPGydi/JTIixYfKsNMv/tZTwiL+UoHRiZBVFKKOx3LAC8mgFXdUdYGwZnPhPVBIrRJxE
Rc1n40BeUgXQa/BvVgZFq1WN5zlUWx0e+VzL4EHCQl8ppq0b9oCO2dY5tSR8oDlWW/ZOlS5/u72T
OBDaxVQ+J7PWFUnUbY29E2dI2dNIjwjCjYqO+AssBOBH6HZcymhsJOjXSsS6xO1jpNeJMejZ9zqd
GqVBeDYMHSNvyuKhK1iLew/SAb/tdD8vIj8Gsg==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AYMh8vGmPAmkV/4T9vXCAbcwNUQ/U5Uw5Swerl5fs3AFaCZc0Qd8qyJ+58+zr5M2R7LYmJxqm46e
wTkAaUYx5X+VmZ+SG/c+BTOKZ03KypVWl/ISK1LXC/o7S+auCccud+8zMCxRUsKHuKYyIw/9r4Xo
hq9KP5hjv/dyE2FloIaus9WXSRmy3BsOrnOz34Y21Q3ThEHJzIUzPC9BzWKJqAiXhmZqFyQNpIPt
k/qfbsSvBqSTLaJSexAjyCb6KJ+cjdu04kb0KxNQHwNLCdnF8ejcSevf63EwGkmE+UzodGVDp+ZB
5rDYdmQGjq0EQCsB9QHiQJ9xNvYS9co+5Ki68Q==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ft/0b3HbGm8+/u8rq/UN1q9QtlQ7ydmhNvkUH1HFaaEw8IoZqW/LGV+djzXBf+a0L7Lslm4B8/ds
ZIPflSuox2viiVlo6Gu/oLKkTEg1tP9VJQ0SBlLuKdd+1Wtm5pN17pffr2TMr03eYDI2Wj8CqIF+
sz9vF9ralD5iy24MBrbk7D1MMaUjK1iYLEbGPul5XaMw+wCbhmYkQz1aq+m95hJ31EOKL5VFcBvw
0G1ICvealfGN8TBm1MOsgcXCDnEIfZlhrRoDLXx1+eTwJ9G46IioWqKUIgceTRCiJ0HPDdCrElbb
sSVKrR1ThH2yUQnQwI9fGdD6wpMKCSYrtlh7xw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34816)
`pragma protect data_block
ewowGykr0Xg9OiH+t3U9UlOPgMElQRW0LA6J5LYPrNqvTAoE3kHGawHvkNQ0FfMtlnF1aHHAvqI0
btSAr96Q338/FgmlJCdNWX2o3GKXZy0WqjyQoxgqiHbQIb1dDdpAsQCv4DdKAFXratcFwH5hqd9W
Mo3lss5esgQwQJdzY24+R8fxoqV18jOu2knlEp+bydblkknaGrvNUSgxsXcXyiTYNvUAxLXFWakM
3xD92PglAFS5VpOuI9Lyr4rRgirVhbKwmcYTkF/RAGjTd2xb4V0NvfA9ganzIQIH9Anfx8ddnVwd
R1IW2FBtSIGCBLxxw2XmdJwXnPcXtuZvMSimXB9Eamxa7R6kdRk2x/P6SBUpdvQxfJgdn5lJtANG
G3V222PF9AWqw3T9EU85AUiBk85kNbrHUbcv3D1562ojhZRPhSgNVENCOVtuSu7Onf6Gn8Uv5QcL
Ffb28WpThQaNDOYPEyF9++sJACjPnn8VGmJYLMG/sXof3oOXpJdeAyPq4bmIETtqZawkpzvCSefd
JRW3TWYvWbxCu2VZX35Fiv6oko2GnPi5PBWygbtDNDd1EiBevmYZS81Va/lqbix/RqwKgBgfLt8b
KnQa0yu7iO26D+JZVKfJMhWk3L0R34t0lHdyLGdpLG3XEaOCdAzTfjeTcaiRbLaThrzwFT9Hwk2b
PHGIu0VPW36aPSRup5TQI2U1zf1vONEjptU9Nt/ktqUoNTyCb4adlSo9k5ZnpGCMfuqVMkDIPK2g
+9mLCZ0frrFo5yPDC1A00DUGAU7UY+HM6hANt3z3GIP7PUkcUsTz2FCwiWm7Sp5quwQ0qipzuOW/
Fd2ew9UjetsJx9KbrIprkC1f6jG98PC3fqko1Mzv8Ux9QgUT0hLmhERa/9+a3Pe2qPK/4K0sbNt5
U9dKn9RyNBAwWsccAR+CYE2R/vDKIC31slkTm+Vb2VncXSxRpDZCOyskMytxlutgBEkGBmt2xtoW
GgdYmYEJHsaKybWfn6U2apRYJBitNEbkR0rys21fmNjQrqCll6Bt+nzdjcduVlApYLzQBWETm367
bWrabSvw7euCBxN3xIeAp8jd5bbVYpquBzA6bpay+epI22mG7MhizvEkC4u0bOY7NWr4y0poM4SJ
0vh8VvmbR6V5Ia1jGITSQG0d7jpbzC3wplbp8x58BiPVlNi/7pgL/5zaS032fEPepvZF8+Sxuo2Y
aukV9c5nVJbWmGyByR9YW92l98NbpN9lj4OlcdyJDEIlynlzBJaezYpeo/nfF7O9DEqZMfh11vaU
SVfqXDMvjcdV9TnxddrOnPPiM9NmbR3FKOK+VnPbpaPsRw5FvFUQO4IzjL56YO5wTJ+He0j+K9pX
Z2nwe9F8affQ6BRjFbE+YP61EaIFZ3A16ZQHonG2lX1zoA6kvh29qpzKrUdAzuH534AMTW0Pr0fD
RTVGwwoMDHYqGA51YGj1BhbAy6ELqO+cGU1ecoCoeuly4YzMfN2lQ7iNoC8FSN7fSmAIzX/AM2p4
F0n99Pz+KEXVQ7Hc0Eyccf2Yb4Z8KWxkuOsg9CWUvmZ61NSBW4EA1t40I2p7BX6i8Ckj+ZXQqbFU
ejfgPFedeuSPi0jhjdi+XZCWvmi4FBnJAIISm3V4UkbRewW/Is3qX9PiYvjN6M3lWGmBOZnekmum
k0YjIi1FiVeBA8A1tI6llIlXjm7oDw+NZqj98BrnEMwpSL4cKvHuIrAiuNXsks7crAupceHyi0Fo
7OGPtW1zCP+jZNlU9TNF1f+d1Ei69mS4K/1r55GJIP5dS7RtYdyEZlfJHSUF/YOXCh5QiqH1Oe8b
pwTR/b5tKR24N9IR0R0PrUJj+9SoRosbL3n4063x84mr8hcaSKjaCv4jave7FI2H7IT4hdR7cflQ
zTtHXbBkcC2DDMVMsqGtTeM4NZ3tNNU9/SYwfiKKcEt4pp35pBiKQhLfDyCZH62sOdnp6cdfdlCj
RtJL5Ug/WF8LNePp86sjwTfVqxPZQPjI4DSL34Nm6BacbZR6oHsx8ZorPBkFaNf11ugfSaltIbPw
zaFvs0Ibc0vuueQPZT1Bh5JtG3Hep1hs8nk7qiomoSVMh8+mNT30hSdYfjUWzANin+ACcNy9eeW6
8mU55Ygc9A7YgL+mIjZYlyT3WcT6uNYk9+T79L+PY/IgpqZ06+SWYH5nAVXQJr66l7dzvvpe+TNf
PU59SEmd607hqXHT3OT0aRXlaIPcb5RroizMw9H6na0Yi4y5Y1mIoDPwGBKcG67Jkha2wUDDCRlU
t5CV77UvG87+f2jl9S/wjYfzPOLacSoGq71Cf/Z+kYJmHol+WmFMMQqF+MWGEXe/pxmn7m9JFEMm
SE5VCJoEtA8bIN0vBI+E01nrcZ6MZGbjPI8Dvi6o5hy3K9e2acaGOfrgnLBPIYkMB73/l113nwUK
uQYmJAgP7wClr9weSdpYy6oBEW/58hyqcjvisdPchWaicBoZr5DAYoFqEWrLsUmnwnzimAnDUXrn
4P4GifBy16J9+E5b6H/4iFl+MpL7SUw0dDvo2zlkDYecz1p7FYpqVPeO4l/XM9OeXNghbv20cF8F
4eC1Vz73jnpBQgHgpmCXu32jv4HT2qqqcqLY5+rVP1pyy5e7Ezec2fi3PpRO8znRpPeZS/vv0gyw
NwHrKH3czZqgONoQq5EEntopsSz+/qgRgKZEKhm6ZiaV4H7qqByW1wnXnlut6UEBMJ/5zUYLG3sR
2AkoglyouAx/sabu3iyO41emt3lB2bZAf/mQ/cc1cbiJnt/KkSk1F/KGgpBQua4tn1PR9chCzQzG
ibCPFXvlL+GT/+vne0yNiwplUgxAXEARXvVIUvrx/ss4sdk56F2GTprmjZ1E5gNKTwuXDxS8GOAY
nDaqQFjiMtakDXg7aumTaTvgzTCWDxWRJsmdpcl1CR7okcXpeBStikI18Cpkprx9KPbf3JswF5L+
QLFEVdyZjDMRYMmInIXpWvyybThX8nc6y/yTpq66X8Lr7qVDxWQNnDMyZZwKcIdxJy2juqH/MMgX
8wIOtoN0m1JzTR8l0nhQHn4HmnB4Ftbwtl3AchfA7XsDS/SNY2VnYuAeqTpFV2w7gPYHyD47lPfZ
tVsz5ORLFgyMeFHfAs/47Svnh1pM4ZFLi4HPmmrZ1vea/6VYhfWs2zhPkKgMOHcKyHXUJZgqiLzg
Js/rTqx2JPdQ/WlKJmOZv6axm6cF5pfmWWL8596lNvGIBropDAErY6Nn+bbM8GahyC2Yxo3G31WU
c4cVoY2+uoV1wm3ne1MQpDL4zMKyIdyKDvA3Z8z/wPAqfxqaDFuuCOcCRjUYApeNDEBpSzU6Ihyj
f4eEldxya3gC0ViSKoPFornCeG5NfIculiW2Mu2aeqTiwC9XmTBT0UDmiiI68IEHwAi5v5WQSPMT
oAkukISqcXMCXjydEg9765rB8orUDuOCROR8lG5IoLkby7ZjB9picEZksqu0AQE0DPSuqlcAOUBa
0HCe7Q47jOKS5S5VBupNtVnbqw9d+EliSessjKsB/Jm4CryTabKHyJMk1b+fvA3guN44itS4rlCd
W3QUBgneF2IAc/TXYz5n/hm1Q/QfSt+xux2x7R2c4kIxB4VhIlgF4yZpTRMasJHlIGbjQCruSlOm
6xH23ujPT2SCEkMndcQVx1hDguN5Z/+5Ca/jPoYKwNkA8QdkfBy5o+ERIkX0XyiMDRfARwGEpbhj
TX2CwlgID9Ku8HQ3lOhpfyPp4bRgfSvPUpuS0NVVeqtuC/i6VLHNioBW96o0qLJA1oa2pYYxRAd9
qCaoDBgqndPOy46lsnPwwWhFFmpxbAHkaa9gaPZPQ6bD9D0BdbT/MKg9s+oH+WQctY7hSmw23jcR
DII1GYwyjrIO4gzWoSMb0a7p5OCAkENGHv3gvKYFPOsLdNz3LdOZWulB02UctcBd3EWzCjkIb87r
nAcvbpxy5nyE2P3BwFcliHsPyKsSpppL0cNH6ePg6mqqyelNSKxY0CHqjGMOFN6+0jxWREd/yP9v
06ijg4CfuGjYgebYG8QNEMZ31q7JnXRwqLsWHyF3v9gRhoZ7wxZJRSX0/qlOX3zZneCZ37nccbAG
2xnvm14XYYpqrqUuxduyr0YyYfpPiJiVE7rIzM/42A2+lpy1ZzqAtF7uU8NLg+2T7aAR2Vp+ILG3
m29BLzQKDBUcoiiW21Kc58uWVB2lzl2bmElR8rUaBwPBxlPJOKroyutK+l1D5fhPcNse7b/trOl+
qVuxXnodMO+YtoDdruk/rke04F0hvzae7vjQmW+TuqK287XQPZJE6oJ5iVcDPmIh9wdDpl4Iv4Bf
RYwniItuOilGr1OXevC6kzyWoUWU3QzLKBWPZijVYBtFcTpaBYm5mcbu8rHOE/abIcBKqy6PlxAF
JKs8J3ayLMQg4BeSDc9v/F8KPaMxL2vkFESgc8wexNwSmbsDvVKVAJUHWlV+hIhIm+SsFpqSD407
m8djmS4JfDuxYbzXpqPZGIvE1IWTqvKFF62FhY8808T/c94bV6HApNq7tmFS21lPCKcA4qoQeuCC
0/iCHZjXwMPji7LrotAgJtr8US8CmfcxX/wOnNz76VdBp/DksbBi80rQms3YhdawQGvLqkQCNuSa
rcP5NpvEZBZB1KDEWRag2I4RdHew8QseHhIbcNF8yvZY2WVmnpl/VdVvcvZBbrY4AmckcSaCG678
JpTmHyzge2AqejKo+nm7x1hd37dH7KPTDzzYJbbimf12E+SaheZF2JaC3hVonMT6mb4B577eCgBK
TXouFiM1x9hV6KOUAJCRG7gYjcq1HLuooNnHwOVd/Le3n4zXEQk+cpZh/L6Oj6QwmoKjEe8Icfzq
G3yU9a+bWNi1OCWKxfq0OU6RV6MGZ0PyEmQY/DugGioerVCuhTyLv9maHD33dtfxXVfUiSBcqXDb
B3SsLFMsk6oTTdYN8h0HkBhlgufTvfySbUDKJAWMP/O/q+iRyfkmKYAaWr0khtX9ZVu0DaYVVSY3
/AmtVVF4rBc8CWrTHGMq7awo/srDJjC6PoI6wTDLOL6f8ZlVQOAZ05Vw9YfufbWIldvMMkDm10F7
2A4j0X6HjTArksrAHCsVvM2FT4meSnRd01X4Jz/wURbnOlCcOO+PMSu8OpbVtm8Ph08KhL1201hi
E7B88y0SdzNOYDkab5SGmfU3D00/XmYSOvR+BSknA0zCBBjRDgyoJ36/ebrDRtfYcyhIgcuBs3Sw
zaV8hofzKO+B2i3lUmuE754ZyVCsADvmvqvX+BYuSCirWUENtlV8VZM9HJk5H2Q83y4YVbsijf1B
muJsas7+Pbp63q4pXwtfcCCrZywxgTTtZxFZ+BC2Ya9a7Rbj116bhLPidMzbgB3a+6gdG4I9cPQg
f9PBS3hP9s13ireW7axLEIAPfMX2nRhf4zChcOnMqunt0dPLNHjc+wMtx5KoUWlxn0ZDtXO/SQbA
LeAPHE8putPSr9GyMrPQYJQsELAfhbeMGAzJXyfsyx6FRdTUe/U2SM0YuG/8zzEhzxacftplVp3m
7JHsZS37XDgFZS9PhzjwqPSdjQzwLYbSWLaiaOXWLGR15+zpoo0dZNqG2AeYRVI5YAAHm2GQNDeF
xv26DWYkc1bNY0X3MaS7ipUoHohhMvAlxlF4Kr1e1fMWkQQQu9nwhT3PPzcz3qHFbaSIUxnOadrA
3liLYpfLRQ+AjiN+ABRy4IHCWO3T9O/jRSlMLCOuN5idd9vqVPltnzJlS2H+g+WAPFopNjhk7hnd
potKLgFcSgtR9w3pMvyT685RlnOz2T+KCCEXlQyR843KsoHmJaz+75S9tPJx9/HC7GQmWAm0l+wh
aJyD5XF8nDVRN/3/CAhVBbuY8m0VRss2dcofl1Qne9dBSCwwOVS+Wuh510eUn6D6GZooXR1bDOAq
U/UrV4RIHS4FBbi5AXRNScQ6U1nr/mWxY9s3cBQ2BWsmL0UKThDfwLsMPkKicu3/ESkEm/ugfEPD
o4NPy4d0UwbA6+Ib7AuhMAjXjMT6RTtXHUdcqr6NNrzC8Fnn/4ac2e0IhNLLBc78qE8wkshWSNIf
mEL8TlhaD+G0ng+DEr9X30eEhsQDP996MBiIvuDf3Fv1ICim1QZKpPzsb1bb7HagIDiDNmIP9Y2U
f/1GvyLH/8wTTd1GoIGXjHi2JVGHcDOk9CwuTA1y5Y8KB+3ltt4yY3vD1p0s2oxSYXv7PnI52xnv
7Go4kPa8CgoEFyCs3ECmyC/atpdM7KZeHsrheAb8vHOXEoFqeCmL5wdul0O3FfrLXwys4pR4s8Tc
oxcS2VkmnmVhMfMFwTL/nHgdcAbW4ajuGxDOD+8vte5IRKv1tipbXk6dziBoMds80ySwjRxnmmu4
y0oGh6adAU1+XWCvIYjS0jpysjqU0xAG+8TKyAWDYMwrJJnpdyli8IehgVqhWkB0iZs5si/tIBzE
hCFUNHEQJIls9R4xK/lPFEcJSPpXkDHrXWQeKcAlo08jEX64QYSEy5Ioe6f1Vl7QnfYfQc+QxZNl
IEcuyym0cc0I10B4JutBD/3onJhYxeitGnKynd9nFsPbnqbc9WO+5+vWKlc3yrgPwUdkUj2xhUnH
hSf5qPNyvonMggyPuJEpAEzn/1tYLZ7DAYgRIz1ImX/m0sGBsAfmoLYYnfC5bVZKX+IcF/xDIeU+
+VpxNGI19VeFPsgRH3iNdh3p9uiwYPhkGYyaIpXneod+hhzSlh3uatNtsEdpcwllX7XDmY3P9V5K
2ZkPnrfqo575/76eVrfWR3eb3Fj020sH6pTa5drMQHJYBNOCjXZD6j+Og53xUVjtCgp8XodV6K9Y
432tbtCBLFmvXK6A/M0xGakW+o/0H1AZ+SPk0GBeVRWhz89Yj/sVZnAf2sU+4L3hsmPtMOlNVJg0
JraoS+wI+BYKTxLBEubtb8JErqHpoVSuPOZ5MRYSFy79+f6+AptKn5I2DTborhmNUcN99ObIsyQ8
U8Gk8kGh6cPMKgh/pzb0ESWONFgvxMBFoUY3ksK9VAo3J9ACqYYHJ4BnQg9HPm/h4rvZGKrWIQjM
QRO62o3xkwVFQdtw1X7KAzxtxUad+toKR+v0u22EXds4dC4BBJpbC+vQSLhtPo6B5md185BONCoe
X89Q1N/94IsLG7lDAbvsKrvhFjuqaG3c5OUbyAkXRmaV+/d+xJ7GSaC04ByhCRKUsQDJzvqW1gaG
EMsozlQ4hx2PMsbq1vUiX2qoo6b8wpn2UmACmVB5mZIwFEFuR82SyWw0/5mfXaYETmFoPM9IbrnS
UcpgwmOZDsXBfkdsR71rOzK9aMoLn1alqDv53c/YiV795Uhq1Dqzq/LJxPv/SexLOmYK7dXCrr4o
z+GSCdUven9bEPH58So94NXli58xD7KhTXbm1JVpLwM6he592zL+d9BCjrt18oB5IzZok1qDemBm
4d166HhiTKIPycFoTvZ/VPsVcfHWv72ongSNgGjXzz7EuG7RUQeThpOF+N+ARsij215LOFl4EfmY
dX1JVX/5RuGOq4n9xBjLUsrNca4aP1cyub5dPk3OivuCc+/T1vgiSIrHlKMPiN2UEZC+OLK3JHln
P04/Eq8JE1Y42n3M9dO5rlnHC6TvIKlc01anjmLStptfqc4udY8onFDeNOaHB5pvetNKrUhla2+P
JJ4Iw8OXufW88UdcDcqDDpzGh3uIDxcF1GnphCVn+BOvOSKfVFzQ1AYhUGU+nRaJgF0BSlA+ZEey
Rb9WbylAmG2PzHFbfhN8xyoQ2SPg7ipyBCJ7buTmKlgedCW8k4M7xsPaY3auA3AlaVkf3QqwAUEa
jL1rjVAyQUfWedYm3fAWscHkHAyWX2E2PUJO7EPkPZKj6Whdvdpe/LrBeJ1FjmBktBdFxHzDRhxL
C7NCrV6RDDxjSqPgMzgPRLfjIfEX9bkWevX5olLWYCJzifqWNj4gT9l+L1Gft5ybHAC171OntYmV
sxUz4rrAtxTubzcz8GsFJV6qSXFdVQzB/W+5JZ1B6Q+tJsjMBrLojxEZRIdzRxRdygPwuWFjyX8A
2F+73UHcza2+87OQ24eP4mn1Ka1rbEy8XwJVeRLbAjdnZKH7B/B6qTL1XtGQYPMrV+uXxdqnw/j1
pV9Mni0ZFJobQmq8U/PmLRH6dXJib3m96v2oFY7/FZxf8hWkfNGF+/7OiEvDT9ijGRorFkY+7Is1
g0/nl0oy2GcvnX4QojYEVLAxaFv1CKxAy6Pqu37RLseKYB7iXlmv6Dd1mr66LVm+aFvGxunR4dld
nxTg3Uo4eZ1gjAeVFeHzNCHu8vyZMHDFc35h/R24xGrYdSohlMW505P0GYkXiZq3UI8sm1hkDrZr
Gs2+2uhRC4JTfwWQt4FYTo5b4enFWtc1sFc9Ou1UR4CoJYjg2k3SCYbS1sraTb7d24sNx7MXJLdb
H/D4BeEQv/WKdtPhIKz2+VWmRfb70QbzpXc2SP7h/WDQCTCxuCvOSESTsAmMwnb5/ef77r09MgVm
oW9eYtD805ToiM/EXIAHWlZ4xCYzORqMCca+MdbB2j4kH/Vi4HURzm2+yVOsdZsiJNMm6AVOlTmc
zqNmX/HAutRd0iCNO5B38ljpjksz2n5SO0/tkKV89oCHKgZxifvetmLxJx5IUDOrKlp/qqccTDcy
HWWGLX4nL/YXQKx+j4tbe4qufZfcT7tzmk8v5ZBz1vwuE5FSodJvOUSSzVqFi5/z1c0a1XCOdAG3
42N8PVL+0ww1/N50K2obK1/n1uZCJZtgrJQZUNeaExJBhXtryIeUkKSI7e/cObkvwLs7aN09A39l
ZtZU8dapO9n9S10BMwAk+9aOg9c7tK29MbKma/LY5zyT/RaKsN9doWvwjs2qpBMSz6ilOnc6n5aq
YTylz+zkrJVj4c3VGZi/PMeuaE5dqVGJ3X3q2ksKlcjsKEcWzaihdNM58xl4Lv5uSR6j/FsJXRUy
w+s5ZS17VGwh7J1EICmrtfNHH66qrt+S3xo4wmh4D4PhFIEv03lBEzfAAc1MmeJdFF4cH1ySERVx
6IN6eQ6KDxvnQaw28tMAZosqFRE7a4brw4TZPDAVWD78lhzZgSitkVvNivFLpQwpoGAB3sam3d6B
bgf1iZ5S7Ti24nKb4WLf7v8Af4mmX4/ho8R3zocX3OqHaBRlMGH+k9hdq3FKU9qpyct/uzBFfGcv
yu9nhaspBWI44V68JRV7lCiN+ID+OjHQXlMVVSH3zVyGS3W5j7Nd/VOG0bwnRGH7xk4iI9h+SdYX
Xs32ENScCkdFNNNJU/bTymUKV0j4kAkh0FJ3jctz/gxJ6ILET3u/Uit28jxDtk5/xaI91APhZpgE
5xoKMc/wUF6XKX0AAoY5oKTfuQP9tODh+WA+9rqNGYRAaQauWYam+YbTLcm6fzGvPrtEStMcfdft
/HYl3H6QZM4zW4Pc9iEHet/KXuHlbOUvUVwB5nZclV3+R2tjfgT0mDX7pN3W//LKQRQLrvtieXsL
fkfieZvr+ss/UR4D3rh3D1NColOB21jSRz5hPR0BBJPqChZltG2cQw2w03RqYYcgG8GSCA+lB9Eu
170W4yp59uy+1Rx0aKxHZ63N8jU1vayzjAFgVINKA0cZVOeC5VjOZOpi4NkkQP6T1yypOE7k1Ym2
EEjPgZZKHhkGTn/jTcn8v+IoqgV//FfMwOmeQHjF5JBch8ipsGRjZabTJIMazTSN+Ym+laUxqnog
JlzxPqLsQUPX2hUYWDinapwcie+X9wxz4ohHkwed75ud0e4fyXVV1D6RASDr5eP8lyY053FHq0IG
/TY/Cko4PWIL/8OwX8op41Ld4G3VJbd8Br3bEln377kgR8c5lakffV6bjJ8aycplN8R1VXrYUoXs
OZBq6G/WDIYr1Gu5nqP9ZuQRaZF6+WBsegk0vuQxJo39Feqyy6w79GJc215Eluuox7ugSf+gpGjw
zppHZtGqz1i9vuwPhxKNE0YMu07y3s8TwO3GVBWpfsP2MEt30QRDFAT/dMWcnIKCBv39i8g9oVuL
+pA2JtWymaV4ngV4EfKZVt4MGzjYGLEbaCL6VpB/bshQQYZferkSrdSv/l4Fq7Ts1WDT79kgneoB
bF7Bkw5e40r+pf7KT7R0oBjOCgfH5/3AxYvKl+kcIINgmpgshIwqshDsxWzNXxs6p14HoEVr90f/
QKF2OCuLceaD05YhwWP/1mx8To5vgoiIQeKLW1dLORksdcl5GlzhzcYNMkZuhbCzca1rKgxK0HTO
vBGy3XV7G7SYioaVXhmstGnHbxpJ5KdUR1DaeLY6zcaJpETF+jgU7TjZVfh8L8JSMSmk8AGQY2M9
l/9T87jhh+ifdB1OgeD9vs2eeGdt7z0b+09IpD0SSDBAhcsthkik2AnSYiMgPGmrDUVhjXo3Pl5/
15veYfBF2vhxMmPVgdOdf6ZKnhD3erBEd560FOefad6yFDKgupC6CJFCeNLEWePdlqkvtZy9eDsW
4uFiXBGhSfxcl15bCHKlWbVQJp04isJXGl4mtsN+Sz9GUPrwydTQwRsn2ZQ69veNlDbFa73ls1ao
dcpX/Jb1MS9oARBY5TY4aPxzg8T+C7rQldgAYouyVVgzw3R9UX7s6aPGI3Mkw22GUXZHB+ej5GUh
dxZG36kdC5XAkfijplLsUAu/5GaK208HC9cXV34IPFw78vO14ZnJYf/v+U6XHtk0j5EgdwONtPga
bTz1+fBFE5vST9X+DbxvT4KPn19Dg3YAANGYl27s10tfFQCr08nJ9+GU8iyZE9iUtqTMrS5OjxXf
Z4Nq8ox3RPOROMjmC/au/LL/Mo0ONgUMirJ1HWskwlW15S62ZzWUjUR3h49EjoKKbjzKq40d40oE
dMyf70gcHdLk7IG5uh/ODZnRXUCPhaMWrZcRFCl0cG4OPiTXdacd85zoDv6h9/wKZOS/rkwPxIzP
UC0PEZlZQntD7LEIDUynDEbfmPrlhkFJ2b0TIMIhEZnDVpy5GPJVNzdZsSJW3SykgNNPByIs7J/N
5X5I7gpeR4tW6eMtpy8303uF6poLLCgegBSL71V4LK8T+jCIOA0CgSs0xIS/9lEy2jEhWRs/Re81
lhJGxYgjM7ebo+k/04o3ZQs5WR9lHbZkIComO7cAzVsbZ/GTYPffRW1gnnrfA6YKtjR1b9GyxL2/
ZgrnpQjLfAdV2GIY5RntgoOoYD4Xl0aPjgr0u4AQOES5jrAD/pbASBSx06MkQPbXW9T+LhS8Ysji
94jPbcRsc5tVvmhOzPY63EJxJEaY6qOUbFJwmn9kxdwlvqkA0sboxlOwIcgt6xZdsxb6F0fcypXq
YQ2dFBbJ/gXVAM3AX4/qwN5ekC1NVos3olqldG9+cvQjj6OhbnAfoXqdKdivdwDjGIqkJ+eO4aQx
ZhdDWE4bhKNbLZpwmbA3Bre/j+wTpn290DaYn69YI9em+lKzfWnjzVXB0KZt2S4+wtJSGwKr58Eb
OXFl7Ua/SB4EnSmSIhALPXJ5bLm+tikM71pGZA0FLjclIAiRFztdEnsoHN/P+QuoTUZL+fpcClVv
quR+xNe0zGErRdNJkC+tdxubJe1OospyWllyWyslj6yfmDjGUzP9e1wuF9EDwmfb/cvVIYpvd58p
/5csbiJDR06wNwpv7+BmOGKlQu2JOUcgKYHvK3rDSaclqZNz90LILYjwzji5mAI6bEZo+QC15DIN
hUYM/du1RY52zoZwqkCtBx2fO5PM4IPcX7RuZLBaIfoFXES7CyN9LHbgbKY9hNF6wQLQ79upveVu
Gls5p5EJYd8XHtazsjp4wXE5G+DGhyzDdmsT0Iv3NGpRHLoTttvHdcX9fkY3fQrvgPTk/TjtNOWb
4zrbWdNnFsEXeZP6s3ttBGh8sLezGGTlT//jjHa25PYCPZoaWrcpBr+SFm5u341cMH6dy6Ny9OAk
dNxBEqpAlm1Z8NVUhqZapkRhRuqmD4kfuO6+1djvKsl+MAMxDN7KXQ+jTqnrVZ641623ZOJU+09O
HRjVL/ph1sil2Gy/ABR1PX+YLV6tOCoiVID4F/RhNT3AOrLC4Ajwx6Y3eBkQFDIbf2SZ8FD7LttF
IrsTHUYKhwkXKNqqSzvUjT0d2FVu7QlR5YZrSeMXDTj9qON9lhfQbRMcxgRPDBc7CcU+NCprWGI5
mxOIGff4P93ezO/tiHmQOtc6m+YQV7wGn1ehpqKKyQXdMKU/99QSu4SeWUUm2rQiYE3IAXb8itlZ
ZMb6Ga1EvX26DsCetFB9T6V+nRo7QIgQPAlnZ6HoLHiHwFFSXSgJRGyfQB6i64+AH6uPWnnsdgsb
CB2DxDh87MV3E9VCwpS2BVjnZRLGAnbMuRW+2/RDiqN1BcoihG47oHpTuo/q43DYi4FfNNmNcOEy
2Alg9exQXVyYcmtwjsyRw0CWuSyYskVAiWEsgNFw4G5rqMeYG5tcf9vaHC7LbuClXdRDNdrfqRGw
Apfo7MfZ1OU5nSS9Tx4sMYKhfqLkP3HebPal/B4ItXST86KYC3vxvYcctt6Xkcio+Y/bxX84ZlPf
AMtDT7YxkAnY7ISuqyXxH94g6iCmIgTPL4MeTxGjhEplChyi6N7aEJnOuzFqCh8BgM2sfdIh1ZMB
9yPyBp31KXhjmtXRmWyX2uoWUqHQQWSybRhJ8ARJGP3D2JJg+nkzACfD59hFWl/7xRBfXRdhRK0H
SL8cEasP3+Ny1U5o11xr/kWGTNPfXjZFdbGBvyEPVoAg6edFWr+4tP5kBlKYUulPxbIxopMThDu/
OYcZPwU644KylIcGhk1gHKTi9J1UYIYtJPd3daJaTBPAqQiPLTDmUdtT3RMQbuv9WyAP2QtPqL4q
rVR2uMHsJ+ruUJ6UaYy1u7P8Ib64ZOsPysHMbm3x2djO0CS1tJ6Wdr0kCM+87rctacIEMXBJvS6d
XxNZM7Ec8HEmpqBA76LTLZKMTu07G6gH+7RMLuGlMSko1VrJMZE9XDzmsc4UQx3JSb7HJyzyvtrT
O6qmw3TQcX3x8o+GmK3Tf2SXsvpP0fT78CkgQwObfFzeUj49hqQIx/lb4kKMtNWBWy15AC02mXzz
NXLS2E5BF15t0HpEpJ9VObn98HKNIfyOzXqHinvIVofJMAcBa3IK5S38+XTpJJQcnaHF575bYtjj
WjK1bJKfxp7EP/CpKW3gLQQ663x3OFrG0BVzUNzvp13DbmYtEE/wRApbBIDF8bvZ8S8rRza4PiGt
vMlkDz9K1TLSLCoDjcu/fka+oSWD/7myVhtvk/NZ+5QnRXsPGjOfxv/0jKaoZUYhAX8nbCphj7vl
Q7DoRJ7SCgQYT3h7+a0T/6n2PaWQVJ5aP/MJDEp0xem7uzZKdLgwKPQJdgK+IIgV0aqfTKdjM7sl
G6QtVZDUgQ6pCKUOasrb8st3dsrMVdWt8mKB/OnkdlVXCK+ZVWZbmIFNj4VcTFAEaOQ/2kU5cbb1
/7NmdjZ0F4leMKqt4gtMW4BSj24Eo/8wMF0TFQIFD84PTik720ELWc4vg7T6znhrfuLAGqYJrMHZ
nUNjdxu3ZvbAnnp3aE7s3DTlrPkPn/tpaJIeTO8tgioyWv0wAHKcsZ31w3HdprH8iBrYqSuO1Rft
xQTv1gQWhkTkp2Sv5pN+r5Mc3joR7NmsMe4xaSGl/90wPLwvG0VuvQY1yRKTkYME2I/dadjtWUQ8
LwPXR1kv2buSuhkYCjC7Im8C9t0xZP2tHNWXPIeB8kc217/S9HIkuf0fEy8v2XavOhBRiQ1J8vyX
Ly0fkORg1CKxBCR0uLAUpWTY0QSDmYzNbg0pqGXOPVEMoHTjVYOG5SK6VT4wnjzCZrMs666TG0V5
0slLks3ZvdtUn1KvhCXR4mT4ViLdbgHSY30f/IjEAs2qO/0TMAv+RpdIK5wIxWKENM3N8uelLELf
2JSFaCBO3pw4dXIFLlXToZGZCrQkZUD7s1UHgxrcel9w2l3t6veABvq0WXMTA2zZuD/F8GwthU0q
tolXUQfxxsHSma5maK63nmdsptCX2YYplRxnm9kR1zrcFBxY1eeETAc7ACK95a3wdokUVHbcITDA
4w18sN4DuDXYVEv5CqKeP1uKbtHduAYjR/jVNUlGFBVbTxeuNVM8jdYzsoFZQwK8Lir/lBZ6ytwC
pnAdtW8T5Lb74Dv5nHUAYgsWfD9Vg8UbQoBWAdrPo5HPrU0cc2I0w+6mOuK7p3EpQySqtlhOiLWk
yRtl4i/zRoa9tzzdVFQkjUTVabD7l7eGq7fJORMaH191FmIx4f2qQRY68qCuA6DUyp3wzCPnNUIB
0Xqg7Q1r/JJtti5EFqeZgZ0q45YDt4lpqPlW/KhotY+1QRS+7dTGFRaOjmDbfhvIgRhAypZ9TZOI
ioPhH0qofLG+GSa+Dir/icwJz1TELfUUvl85/B/iiKPUsiSj/m6pvmBDzrlRrU105KyiRbMaQToi
GCQD8GlKStmKr/ANiSuALLPeSTZnF/Hgv2pvs/lqqCFTcHmbFOY89oJuW7VjZixSyxbwbSAMipvt
ptafyUL2pTJUC+K1PtU2ummCKYHRWWpcLH1XlVIug26gPgNb96FSZWU9qW0js6/8xXvk93k2cYKH
XE0k7AfvS4vKJrTyNupfMBdQ0OCyCPWNom7bKYbjQRMmUf2VeuW3lZuOqaiGO0NLpoVbZxtgM1Vg
OY6Ff5H/F8A9130YI4JCdNZgDTGVhsqAVBABd5SbLoInId+q6Yw8RvvSfMyPJifEkQ2OsWJGW7du
Mw+yaGDCuBzUIJmcnnceog5tUxT2aZ1qfMslrRs29j6V0xlqaA+rIT4tC8bXbZIbTcHtprbkDEfI
bxeZ1ZJAKyXD4VenjQTK5n1lqH8qFPi84t8k8OI3bBcVUtAxzfe/GU3FnVOr1uT7ZH5V3q7ABiEv
8YMH2Z5nIB2J5h15FGKvMOoDI1DEsk9wCue1tNcAbyPOLOuZkXu+DzmQgAXVw4txPflEsyGc752q
cLQFAlgNB1306iECIti10VFdOpgEiY5bOebPpXE7ijuhN95VVKSdzmPEvRxvAxFh4YcoFyfXidFt
3Po4XNNyukVc6MOohBWIEA/Hx+Yok3LM2/JlGvP9bjz+NpU0zVsE3gkXtYvShGoJobl/R3SsWMVk
o0DLTABCEpJVK1BQqr1mu68UFP9m5rxtLJSpf84tkpIAX1sCwKyZZYZEfW/bVtC4NiHbNurLlYjf
/HRlrKFURHWhatk0vHENC9TFbgDN3dEKGP+LBM9D/t7NtyP1K7I/QzuKvk2BljfoOSkQMmyVDDCO
saAaMlmZXeVKqatUzHyQK32SHHWRpUvh7+2TIxVjRtpaAMFaLr3IUdYRp9EPgcml0PJlHSQakAIf
5hibPEhF4D7RO5pJ7MBwGavVag030j3smDGwrfBz1kh02/nLwSDRTEHVuFWIxELvCS6o/Jc2fdND
Ngcr/kQXHO4vgreQ8bq/kFfr2xVzmRtxYUPUeENXTDCq9kUop5jR0EpM4Fyti8j67IQERzOB+iDE
SiPD4b1Z+uivqaV15OIGScCW4lDodg9W2I5OK3jUuuZf6oNLzzDz7C6QCK9DWiAX42zTIj3Zjmpx
nOTIMGSDIoWM54p7pCoJpl55DcqWm+6/fhFpdOkuKTDxePr5WsNKhM4gr1A3hokGyEx3JLhngte7
t2Z4Hn5tDZ7/ZgSWwufOnpxLY4Z8wdIwnj8bmUZj9z0dtrjUC22krtYFfQUjsc99Oie2kP46pCGf
UPuI9tZ6gCgj910SjNBdKBcOzEVl/rd85YQznNPC7Ed5k5CiHd4xnY104J0sd1owvm2Ip58xKGAG
aaVkrxqw9bv/MXgZwe2X08WP4804hGGf90knR9PZLEGTePRppUy+2PF9bdoeXZkaKSe3y8TDR5lx
NkuOWa997Ny/7nQMNjgLOSIhmhV9li0wT+roqC00CMVnjjnT8ySg9jr2D9qNPNBhzWncx4QPAR/w
pqAVBO74cSCD2ZYys7IaBEID+UwNXHyaRvTTUEKTFf8wtUFz6Ij1EXQlrc3+8xiqBGQGK4iaFFgR
yEV0NFNXWFQxy/S3Ga5mY71vKrYOp0bODcdTgXhkZIlsvrXDx6MmwbDdThze9CT8myz0yHxG4hOW
p0xNtjxyWrPm15khUC9jlM22CEGX0GfSZ/rEJhfgqLJdRDA+c+hHuygElFh5KnIpN8OI+YgCi1ol
UUI4U6BvjfU5QnrdAe+5ATMEQRhSOqK7dDxxOl8A8wfixsMwwEwq1M+8m5a0HLDTmYth4rHQYhlA
xOZHeyMe+G8anwU9+4LTv9ROH1ziwTvP9E/QREgyiUyLqZsjH5UFCbj7GNoLfpgH+UrpIFr/jhGO
/BEg3FvclyD3b30hKvCVje/NWI02sh7o8L9sFirgg92ZVgH7/W/9c6kFtSEEAb/mqQ0ewrXnPjdP
cSdh2mgJ7yVjOf1vCcZDl83MjZMqd8x+ipVrQA6bhg9xPeS6Y6c7JdgAW8Quh0EElfnXHl+GV8Jn
Ajykcsv5YswmwbgbGNvufJGnjhA+5WkI6cFj192Hllb/FM6ClMpdhjOxy95/re+/3S7djeymOzD2
tokbo7AVfbUFur3bWpabstzM9bd61VvReozyEeKiM+GcT9cG5Ozdl5KqOuRXW4aCOv2Janu6VPrq
v3OaoLHsHAVZsh/ovpBdcc+zIJR+8o/Fk570+JQ8JeeHcaRKKeApNJEqaPMlQYORPyJd7/PgAZXa
pub1vdBVxR7Kkt20EYmi9ynLyfB0TvondXX9Y8/jInfTEE/woR3YurahiMDY7E9Yh33qHLkdODM/
j4KSeX9YJ0i/SFCRMrpUNmbHNgxpmo1JZB4m+P+i4fTLvtsoivFE0lPckQXG7+uRg8wdd3PF5AzS
5mW4w3AZJvLwK75G6sOtLflikWnimEG0Tvej6IC+bj2lil+zK5Z4IA2pB9P7ssO8xqF9/sV11O93
EXn63a1io2JMXDNl5my3rpy9ypJn330MIqfVqkuumCBwmkvOZ31BRDpFHWsHKATXr9595FzZMfi3
52bNW3Fq6d6B0EHCGE27i9fPkPh6doGNj1070h7/usGaznPzGcqc5qVOJAfaKvGHvL7+0Vh3+qel
+MlbKS/Aunlfm5Qn0AuuEh6/JOJc0jKdpw6uI//rnG9jPVZPag+H9rRBvgvUi52oVxNcCSbhEWHS
HpBuNe7JiIpDefFUxyGs3wKo2ovUcEkvsjwmixZuco9hdcR8J/yQOm847n7Ou5wM+NTtVgdHqHe8
E95r6cZxX0Vn4dM17/TbUqQ87gG9cN9M+HE/QDgDxe0wjJk3gGr+AjZo1ipVmv1DhikYeat9LyzI
i8lFBGwQuJMIlSFRH4acNSkvjcPcywNrn20e/JNWJIRrUccjU3W8YTLiIaXBYtmyjZA8he1Fvpqh
Ve1JXo5nLFy5eABj8BxJxZlxrJBtTSpxccpERfH6sb8csYLjdL5GB1uxDVg4jnSUVgi4QPIAB+d2
9gAhwjEDAq5xGQwb5r8Y6sijrsnl7i90OLPI8Bd9ogZDKFv12cr2HuMuMAHaPo7pZkXqfNQ3Ce7D
jmwEZllB3qLGlXem2lgx/14Rq8I+qNZs+aMX8t8p1B54v/QfxhOgRCCn6rtiOhP0mtWBvuBg+ZD7
k1RdTgsz0qjO27UcAKPFyLibeS5HfLslDRMW+/GW/NJSqAzCckZl/mKlhHw11DodBuJyew1pDatd
8suxeQgz+x8cak8y+Hx8TrkhFmFL/kgyn91L9tApdVTAUZCkSoNmdGClonZFI2dDLqa8UeNOBWbT
iNG+b7DRweqmmvCvku6fgzqg8OW+vukuDDhGS2vbQPNuRHl7nz/qydQ4fW1UzIcnQtT2RKlbo55U
xGXpTihP4svc1kz5QeNF42NFa4Uter/9Y1r6e0izHZeAFpl+TvwHzQJmcE024i5HkcJObJlcU+uI
HS+rBOLmhtoynsU+k4K/B1k9yKtbcBLlLtTu/0er5e8ZK+DoC6BPuEcpp0cZKjeWn9P6WE7ALCnG
4APB97YCMpLis+KBJtfTk5dzC7vOIrWB5ndseC5TI+ZTD77mQmGy8XRmpJm02CHuEyHbWiR7zban
ehdclWUs8gLvsIVjtvgmft4KDNcuGFl2X2GPqGKuF/xjO/fqi0hPTToJcDAFpnd6vCC8I4f/IcP2
DS3AQ/YA/iPzsLVkhwDzKLzEY5mCNS3Jruguc0pr1GGA2K3AzOJWP1p3Oo2zGUi8eGg776epXU6Y
SKd+bAXX6xXdacMc1Y4Bxhweol1h30Mxlv4+a3JOzknGYAlxulDxVQd2VkIElcOIfGwdVoya5mki
A6qj0/d+VR4h/VbZfx8/vmjhU8RN3lQhxBGorm791jUtHua3KYTI+Sr3IlemLNbheJygYDLe/LkV
FvOH9T2rLf41TmeTiiy4Idmz0xlN7KhVn/g9jnZXr+IdoYycoQLaKQG1vUxkkXoEXGpRkREW9u7f
m9TVjxOGs3P42cjcGbUQ26VzPhesgXrckzpKAkXLAbjc28abh0duRv3jQzRJfIhCMP+h40OfRVyc
NZzVqE/aXbcmymtybAbwMl5n6sFUmOWTHEdaP30YhxrRa1DFddxBLf2SWnv4TKDT1aFgchm7gkRG
0NscfYWFkZtZ5x/0h6JpFP2QcseeSk8lNMMbh//Yt0jsSE0gflXhzO9kxoSbhw1EIPZZWXdhRjKJ
k32nlYIL2HIU6Uj7eg9da7JK2hKW3sAQiKRj0MAQtD4lnPuZ97r/d/gaidU2mrLnMPyTZs7iRhSQ
YxZlNBJ3LyaA+ORLmNVFOZG7uH1Cjcz23hm+QuQsiVSK48QETqHOQ5wC+goSORMLikwtNEp66t3r
r5MMmGKVcnHBJYS6RdvSnyJ6yC50+c+nDXoYgwnHgFSpQuJsffm+6kGd0erqG2dQqNpzTDolHvrl
yKFlbmhp54Ie2w9jvsFk8AOFi0fhMU1dJtMNQTlWnEyu/AOPznWLmkVLxYfZa3Yc0FK0Mj65U2yR
pO+iZsmx2q3Hi6pLqaRfv2fvOk5Tx9dZIYiWZmNi4VfL9UGo4OUJRCnV7eCb3pV3CXSyrGKn3elX
5pM8W1/sEt29hjNP25uWniyFWnfc40RQb0TKcAlgnWmYRSKamal67xTwFdtfcFhJCb491X91lzdV
lNebzwebsQD0jxK8DJhzWFTDq9zmhutA6rb1dswG29jAk8PAV7Fp/+/82Efc01jxHQHLDgkKhXXA
VSAq3xEVogFE8ksBUwosuC6diI3WWDOAuumzj12l8eMtGKYVv7sziCO7ld+sRi8a+nFxs4AZJm+R
aW8IZ4Z18J36RA4AqovDmlLy8jHVOjy8nJEV7QuSvPaDZix9kKJPjgIdHqbFaxdmDvZmuQD/5llZ
U/TTHvYUcTzbERvCaYmExRKfPtVw0qBT1XZLl7IhfETYoiTNx3mIYnm0mxM9AGoS5R9pizbfnJKj
Nogja0g+/XDcY9Iy9lTPBINAvOaClKw11UNkv6CA9SrYnOu+qcL3RkHJpaAAGERP9RXwYQFx33iq
YNDBn91EgvyySzwJoQnt2Kk58TOlwA76mJk6x7ULD2BvhrlOyhQt92PxbR9TZ5Uz4M9iOIM8cztI
DenetDdbfpGSpVLu3QZtES8cZ0e25Y9ovrUR9//t1CwX6ZK5wJn7lPG/gn/gRs5E6giKRGc5+eHk
Zs/livvM+1bAmSGzj1hxy0ZaR30eIE4O/fXceX+ZoHUkgZiTV/pPeoI2ImcR2mLrquaowZ4UAQzL
hJdNGSU/TFa/BmS7DWYmLi1inzhZrCT4++2a9GvC1JDT762Nf6VcHindoKc5E+XFYVDuMMvf/TeI
WuQMmNj8ux45IhyP/OJxjzi6otvwoslYk2A8UWM0IA2Y85iD+tJ4CY3MyMzgGBGrvrGtr43odsiX
9ab4IDOM3jWqTsE4WxC8+wUuAgBTiNjIJHJWrCbWJFLmLu59UxeynPnS6UN4aPBUrpHq8kJscoNp
8BkLVwOnqakvN7FDwBfIvOeavH6hrBu/Pzj1Nn9ZULkeKtEHZCKaP8jXOivT+eag+Uj9bjztK70e
xNXiwS2fGcb1z3r8eFDYN34z/a6YCqTBHynzL2UL8TYBnWoIgL+bnb1X0Lxes20K6l8PBcXp8oGZ
TnXlNhZ3L+MvrAquG99zaFOihU+XXvV/o7X5NQ5+OpbtZZuze5ZtvaGTXVyiN2ylpcAfreP/V3X5
Gfa/n1NsIVLEDJSH79BGOXJfZweVg95cSNkHQoFB3EbZ6N4ndxG2NkR89jnQeZ8mijRnBfOp84La
+E5HZGD93rStxZ6h1jG2LsOQswzK9xKn2PRUiJ/R7S2ejsXoR0wqXSFtLBKUE37bL31HI4LsDBw3
1LiZf4Bpp9/xRjC4z5HJ75/cHDT/KGt06W/7C0TTLMIXeisel7VahJ+book8+yx1WX/WTJv+fxqL
utUCyE/6uTC80ltAdRQ5CvGUmGxgR7ru3sPIgrliDaAd41lmTvavFTxXqzsKpPz7taDhH19ekOEd
V2NjQZQo0g17ODri4UPxO6onG2UZuwRE0N3qBTz3ip19hEjXYrawjkerTj/nkukQPHaqbJ+COzNS
mHxztaWp0+kYNpmL3FaRuSOf9YqzOOvLg9h0gruD8GclT1quRE3MguJKiVUIZHpex2Z1atcWeLyX
g0qxbBjV0WmuJ0HkHFedBmWURqzcM5EoX+1JlThGoiaE6Nz4v7of1TbPS5HCfC8l1lFCiMVjNet6
WpWvL5k2hamCd4Zb3BggeovyPXoHkygcAQbXwIBWGwqbX+EESXcPYSRxyfxhUd56FFvXD7vLSTtB
hvWOwt5pC4brTAO4vCPer/UZVBARIcHL92IjeQ4d+NByipnmmUMWcXTUD5k5xU/rHs8N6iVtA8pT
SGzdd4m5eeFSsnxVVzGRGxWuy4m+vlHcV88gKL5xBdV/f8vq3ZweZ0hIs/4RyYMpZFqGNmbX1ilO
WnvMaa0j3uofqzhnDrJvzubixPgWbc+KuiqLBMxrmovSIGTQRLvknw6f6Kb7SNk2lLWque/PbeLE
jeFb/gLn2uiwriFPu1GI1yiULG1bfUIwpUuRa3Au7yp/fvttwCvzoHXNcm2UwygLu+hAMPDrWOqr
fQGVvJxTV6TJKKSrQAN6B/AQhgjVMZYuk2VRufH2XtZASO5o88fHh2odEnwfoXNYNPaHx/j/pZ6q
oxpLXEgVDL3NtLdKfQV0P2bx3rYYCqrXmxirbSJoHIsg1PDxnVfZuQZIAFh+pINv7XcJInX+uQ99
WZK1h3QetOAamFGqgT3eNsHrsHN79sUGLiNMoAJg5KOq/V7nMv7sibitoP87S452LmIRNzh0tVfT
GQdOFHqjeMaPxy7VvqV04/zsHygCSeIdj/bp/aAauXcyM+3w6Gab8tw9rCiGhYtb+Jr19jUCCQA0
mlEuROP2Zs8NpcrjWnaPbDhxSCcWYT+RRaF7KYYQeLId3zfW1Zno7yXUpk4cNI2GnMHZSgIQWCQx
CNJ/3A0oSSQxyIljoJJlA4pEKte37ZUy7fbg6CQXy7PpGWS6W6ZC86t2aS+kpY1N2y61bHIAe65B
9vi+vqYX5zkXvubQrXgOEdB0h0hfzvGIl+BO5PbfarVbHmB6oCjFNPZjx5zYsMnIRpjR6s2+qVmP
0sWVGZNaKE5Y9Wm4XtzM6ZuJSYYGadBDsj06IFQy9S3k1+bbGn7hWQSA6yNFs4dBaZd6qp8Y+jVu
WD+5msd5poukr74/vO/BfCDFDVlYJrtHIQsWp0woRFuqQnrwOBaNlohrMYLaQFcNffwZF4bkbaE/
hCCMDtlPJWaH+gYE7cRhAqoazrv7tE1d5dRq+0wbNZtsqMloYOj5a0SsWEfuTsxDT7s7Yos3dOYP
4MsWG/WOXV6lK8iEROvk5OzMosQkGG3y95CyFj2f1OU9N/qhGfPCfn4QAoGGitEMH9i2r0kZOU2S
HSos0U0xa4FkoqWJIYU/M9y5Ks7Ql2d9qizhEpfIKKLDspspe5L70ewrHBrgQUyAzy38Ie7i77fC
hUn47Lf8cdAsIzJGMTSASsEar530pNsnaHaDpdu0Kca2kyNO3Ekw/7ZYWTJF80QQyBXeKNv13I/s
JwXYzSsDxWmqlWBzL9RzMKB2QuYjCVQxLiKT4m2sFiZT2pkuvTOvsRpFQiNltsfTgKNtlPeOV80Y
ETa0DMgSwWPR39nc4tXWZMc9xlKBRhiPgkJ6l0xK41nCuy6J9MiHaECnpd2uyF+6pOGiQ0+f6Yu8
SN0NhsnxA1UMjgTbyU8nUVv7+cZtOuA0t41gdNNhjKrWznHrQd0PcS8aJ20TB5mJWXAxF1ydDPvQ
wqvF886QxH6xTgSRKcBsMPImF8bOoWRFOUzTR3hLnM9dGhS3XP62sAqCTtxkTPgPGAcJ8dtbIu/1
KvK/HiUAM1zwR9uCTLkmMNvUWcfpTMuCDjxwTBs6wiEznZMbkq9h6FnWgDp2/XVO1WJMZZ34lOrt
9nrwdwTLZrTNc06vcpSh7EAwYVOoR2veGNb8vn8R7Zr8fzZKTtAAInW6Mlf7Vz50il6m8X9g3KwI
r5esgKXYRFEtQafJw9RnsLdaj0Y3iC5NL0yWcL7MnznlkSSc/unuGSh9L9Po5oA3Gu9qqNbpQCqw
T1S2sAtyzDuL2DEDCwno9gqmVdMOqu8LP0wWgeYX5vn5icAnvl7rrDEThpNBA+/mHS9Gvr6Zb7IL
qJbczQwxuteQf85QoddweB2azNJ/Cw3zWZEZQMaDJ3XrdEelbyY7L7l1o6ch3bTnv2nNBh/ZZ763
WMv3xyveRqCgxiOmuqopX35khXH6E93+qcAClnmEbK1/xVNhRi/r0TqbwDR1LgHqurKwQpWYWxpI
r7iQyGDciLZNLQKhNAeJANzqbrt5mk7U2mfPOVdly0gpbb6d2xRhTrU5SYiJtEJyQETHHOLsKQtv
6YuQR8nsvZ5fsqU3srGKMdSHy3QPaP0b+s+xr0mlQlbzpS863rfQ8QPtjeqNynynWUBouabcvHhH
Bo7BI9sA/n1DPtxWXCPpjKHq++9zwZVlscUcUivcV+hdS+UnQ5SYgAwpgXU3xU7UG5eEO+l0LCGm
wxqfzSDpBJcPd6ZU0L4FDR9ppXMfa05SPP2PPVDxmgsrS51boCNXvL7VXHhVNKHA7eHzI5QtNyHI
MdoU/UrLnOJKGivoWb9NUGBJE95ZlF/qSb6fU8zuwdkwYZ5dttJqXQQkxylBQkVNiLjEXAocv+DS
sc+Jss9ZuSZXHi7koIroa1cXlFpt+TCA/yKWlma+j32ii8J5q7PfMWW8UOfWUNmbRJJu/bDdRylC
r0rYRr1zonLQQOGPEUvQy9KSEyHl+0OsMjifhN2Cz8DBcPo6/NbWQdavLszsLQo7Okw99wJU+p9o
+9I6ETNnCpGYMAEIRBrGyLLtvdXZ6VaYAWwOfj5Dk2UWrrJ5mcNtuT3BGmSG5bFn/mzkWE5IV2iQ
YjMTLhUfRkl0/8yUT440ga1lvDbhvsKM57ViI33zAJomJ13DzpnOmtR+L4EAo7XeXdmZF6BGXLpN
fhglNpsReJHE+huEqScEyOT0xJ/hfco538g9cMnyz0vWjKHY1LMnTamM/rCtxBsMQBiGW5ncXfxh
zI4ya+C7cEHw0srn6pINmWAcLNEWohM10hiuE+qU2+gbW74RL9eAQjuuQkY8ipJkoez6lIVFHeJC
z3b/xGjS1Nk7fS4T4X8vjN6bnmK1apsOtZZryUDw6qPVHRwUwTvvdPPrzt3dysznvsOr/3kMHqBq
YlGkTOmKumCAptZcCa1sb9UtTQRocK7GI3tslOt4tkYsOoeN154DzjGdQSqrDh0RHh4EYPfdFrBF
xaNQscuQjhLFslKzSyvm/bQCFY6f0ieKsXbpAfwvucldIMUHK+NiuTcQ9NhyfjZ6JzNyjOXX9k7I
v6CgcI/WPId17RnaGan8MUoUcx3WGIegE7olRp0gCF3DuP16FzWgY3+Ni2GMf70PU5B+Z0Bqc0S8
tkyc2QdqvI+yiowNVGDWaCZlP0UTdFACxWGSd6IJfeE926akrJEb5PgNcmfmr5GFz7xA8/yZRQya
KxxQI7UzgM/DAxdN+fZigpVK9hy6DC5WhiFDhLeehfqSBOodBo3ULzwTL/xBgbPVCjH2YknR2vTK
mcT7eLIJfsnd9nArlPdze6hVm6DO0/2ol5+KXp0lLP80Z+YO+VozqJQ+AFnJzoaq7S6fFDCbIYVq
NVX1B25uELdbInke0pQGMulHZmB54QCiMwYnCguBLCMvG1dmIP+pKgyCVwcJda3N/nptLiEjw2IQ
klzbzfh75kOLn2oCjIDPnqHp9KLE7KVhYy6l6WABPYAis6wbPyATfAoDyY4aLCD8Nhud93Uh5Q4r
MI7bhmkOx7QbJEljqCwcSf71mXGblHtL4dSyXWjwQ7gbkBcFuFv7Dg4U3hDiftcgYjgDo/W3UHJn
Eeekkz9/B1EFtJMlTV2EHm3eBIOuj6+JCjNIz1pFiLPcrv2XIjIXObtqKdUzoOcMsE5YrdfdLgK2
bvorZ3t7/g+R2+/zRiRlSmvquh1V3VwVcTgabfbdfNcf5Nlhs5dTo8qyoZu6mGLc7lhkmdQ2YyV8
MG/a9WIPyDcowif/qpszO1nxIMEz3iXM7scOY+lQJZHpBLm7hzVwoyoLXylyufzpSnRGN+l/4pWe
ecIhH9P6gCEN4JwRlf7i0QBX0mDRRuK01FRVkCZxJuAeWgl+PA87J+XgiXkQZeK6gh/W0Xdtk4Hp
WhZkAwiwaU7Kl9EtWFlejsWBQTkp70t/ZnXexSzTMch99IVg279ca/ZtBNuASA5l2FTds34pJ0Ni
ipLMTH7JoP2FEDa5/JpGsYQI4g7xATqvmqkRPWysRLQBQoCgyu5A3isIaMNN9l7xACoAMIAxBkh2
CpqjS9IRgN/Z6/KnzFfOEbjBPuAUuerw/BAS7erKckwMh2BV7GjlYZwCICLKprvcG6mBfXwur/Yu
7xGiwwUYHx5SkLWK5QzQRYg1JbGcXyGPuv2zBxCflUtkeMMoofTAbn/pzJbJ05ZCKqBj8B8l9xXa
hUlGgDkirLpkPN/+r9U2zX7zxfaCIiDpaKapTbdBNHebCkNZy9DIWSVZzePXJKBu7L0nJJDjjavc
z6KUsPW9gQqj82FVPLPGVs9INI5SjvYpra6rSTUzeyXTCS4p+yE7d3FiCBNJ9CGZjvbJHaXPFKfH
9Kechowy383pzf/gHyjMH1+hVsffHoNTTmUGs1Oyb9FCfyqgzim+URo4QMxNnN+1Uoym+6ron5uR
FyulXl0NqgFTOMgDjS3KgW/X2E2ktqD/siiPMSiBpBbTJkO+0jQwmxW7YrcDMmf+c383y/g13rJl
+3b1zMQsuBNUYODQmmk5YpFMsFfzCYADkQwV7KbrX739vkgMCQWXaBim/zNyZuHagZxh7gKLtpMz
N6xThQP8j2u/5vWB9xz/HFhrHyuOZ2JCDhsj9F8NJiFB9z0/5a28lms+m6w/Tj/V85PcP01p+rdR
8n/1uZG0avTjWtMN4Q3d8CajtJY8dAYnEDNBCiINFmohFDVfr5dJBhJ600DLhqI3HDLudBtwNAsW
a9H/iA8i0EMMeoG2iJuAnY0QM2GEMjdtBwDBc4iDAWFhPl/XwCuUxMiKR0QK0q5H1Xnr3SMwJGSH
ySbfIa46UVkYNzf80ydC+vEQmOL6SpEgCUubO29hghq4+v9bj/t3lcPP+cmq4Moc3/0LhchslNVC
ohUUPowj8Pymajmay075UaJHFIq94odaXH5w/6NOOPGYw8wZP480hWEIh+yzIpx/7lb1SistDULK
NayGeXZAJsWseky4xjDluVyzsSGQmqMGZb/eo1vpMRb+mr/k1PbUd6GMaOzhhjuSaqx9uhkifSFl
yGNYHkr2G8kexhV1CVoBgyY/PFuxCS4+bN2wQ/SyI+kFo0jhIEdXBga1/yvZpcIQm6wdpaFuWDt4
Wj5a028txjko1QOc71MBi9ew44iDnl/A87qSzpLNEtclaKfUIJieIABUb2dYALO17BCuoEjKosam
Ns841km3sLRXpo3el4F9TQReG2IJcEgkGTL+fJgSFci4N3f/JthxBKUJzeLnZ1OqsVIWta1s1D5C
h9yL72kH25C0oD1UUn4gi5rBE+xCpZfvT62p29h/eQZELE29BFpJ/0Z8cPQiKdvtRKuxigWf9EeK
naYhAoepBYkZkO2BZpUfgoiwZwsdhzWeD+Dfwn9zDbnV4dKSdJuBqDDmPbBcJd38QGQNUgKkW8EP
vlOZGCWvP/s+0VXcFunMHmeI3yrdBzorBIhCw+LtgPuBLCtknNHBsVh3HPUShHafD8OqHTae4ikf
meAAjixVHxRhl0R+Row5glPjhqvLQPSBrJgqvH/Hhl4MYf0Vidh3jbWI0Ph8bBsUrytTXPIufyoc
tAyrKzItR8PDu5CV93R/NV1co3EGAr4MHRazp1WB1ESOD7ES1LiVVW9K5Ly04uo5AgOJ2zECN2WF
hdrv/1iuEcXELvzS/sHKT5S+taw8fKTTjCSQZTMSD6CjkxwLtuPMx/L6iY/SbC+jngfyKAiMxYOQ
OpeIY2vhiB1lTi0AaqZSpRi5lSCow80VHDva9AZiGWcX4/YnG1R6s5n4QGz8z9Ax80+PFC91GxtX
ZXfsyh6LdtdkWRKX2xbiHTw4WCPoq6w3pEByLpSBy8ojgGBqWEhEwFSmZ21toTHPQJCE54DrK/UV
coJO3mCYbioKhvSlQwcasTECh3NIe3tUH/bjtg+/kezMTAjuRAtjsrc2lowu9+F/y7qE5LfEeF23
spc7Pr48558SmgEtulWjxSUrMB83bOmCdCMUz9t8yCRkZ8OqOOYcEkikwoyM+VbRaf3jt+nIDwJe
OYKLk/+zNxP6VXNv/8iCxoChRKYJ+FRhs4TnATD+Wpz/n24JV89bDKGoYrnXOkiu096PE2OUpPHK
+d3ZqzhLoPaAfa8Vy+a82A/ga2SGlStbRYjpHbhq4FbZZO1h5M0sAxB+KmcwnptoyGsS9JyMBvqA
5S6EcKDR3YstybTy8MY6suHlpEyQLEoLcBd/G1UBnFP3xOAalrMZTQOw8MG6PXRRh+NDjH+xX9Tr
W1tFkriax+cB8moYNB1SFUm3K2MySTirYtc6/A8I2wpxhu8QAmQL6oFfQKmIk6/TSDIimO1wabj9
Jw9VzLelx/T+DvyBj59Nn25UC+lQ0z0i6EoQdQwFH9ZaNqPk7vt0Krt8CPIpFj0GlYAlVA0AtpVk
9u3OoSpfScgSJVcC7UeznE/nujcKrbV8S9Xrl0Qp3kwwHb123I+DT/V5FRI4Yw9YyX4OTKI7/zq5
ZPgsPcc2Fzc8SaR8kDjOQcr/ZvExxrgdjHTU09rlJN5yNf679IERdofqLclCUuokq+uOSEDjJNeY
0vqdvoJdgxzRuIyDD4mtN+CQvQDifQmxknCETd/HAEpsWwwrgDgaMKIIhoncM0cMsj1uT4A1jfSh
u8HKBPepjXLlXHXk55HFzD09Gi9izcZud7MRwuwlWsDprCpN6ETJUWfA4+47vygiFULO+vKRSVCU
eHyHCSMLYA1z2DWkkUAJmvLlR5tnPBLcSDHNrU17U5gGIrDX/ebXSJUtyo/hmfioXDB+y749v0Vm
86Y6x8lJ74Uovo+eDsj8Bu8W6egz7jcTGxASV530ESGlJ9cuAwftUnpoMA3R1d2a+fn2U67k/v2D
qBcRZjwAPw8JkTGnNV2QPngxF7u/bSFvHxgcPtb5Zzjab/IEc/n4rRWoUf1c660O1oOtwuDmh2Wk
OtKpvIaTvGxFOZNqWVe1N20cH4rLkswjgk4+afc/GvCEbQSE0JuDZKRpbR5TlpyE30unwH4zCNEw
tO2OgZbv6f8Ziw5qThgucbfGIqmBEmfzr7JcE8g2+QUGdXR/6QGgyv+dS7IQLtoYCvwh/8zhp7ma
hpEOrzAMaQ8DYGI6hPopc7m0mNysvqwNaLP1oFpXED8iq6JI4SX93DTNBoowJ3/KkwLcOsotl/mH
cBsTzPIYDOq7hygX+c6KfsMtAMD//xZMUcj+/DYJT+9VmBU5ie0+5TQPUXjzLH4cMehREq4fph91
cJeu4en3ekjIaiVpqxJEGJyFndrXg4if2XyXzdb3wZBtDvu+cpTTUkUoTfX9nGQ86x1xfGKtyXym
EO3eIBSfiKIyFkjJ50gUXdXM2ckOzZn5wpnRrBp+Dg/C9rm/1+MRBnaCN4cAtvTO/HuuXkFaADgr
ptn2WwZ5RtAOpWlv2Lqtde13YItY2GqdWnrgjSXTQbikXu/72xI/PBcE++SMGAH8P2aRxo0ca3t6
V1I7lH3ZDT9k/zt9kWGBjUiAvDvp0jOMUhRVWhBYu4cq/1jp3WlTu1rfEIpYJjwHgmCf/m7BCP3C
CpSUSHwLjqQUHpLjddUAXsfXmtF1CaJL5LVtihhcDun+z45EVMy8JtGybFP3zy/gYieiVM+tWVgQ
NZJ91e/BSmct3dc6wV8qEZCuoFM01t1iAnNbcnrSC2ygToOAO5prTMgMBD6Vi7+Nfr+fbUKczSvV
s4KXtc9rBBjrrOKPDa1rR3oKWAoNxx1zb0IP4GeP2S+CucvdGWeghtNpPPgbVH8d0FBEL4PJh3P1
8UCTGCPCst5TgBtsfcPJh0bPm/KtwZTH/h3slm89OwUdqAMEBT7tOVYaonqavfLtRgr86CKCYT92
kbZfhSN/m6aYeXEWAhPjMkR4Iz9aXfgT3mncQnSyWWNJgBYHqLElTFFaUjiFSVJp2Ouro0KCp/j+
ksihjDWnS7VEYCxvQT7SuW7Rv17cYUAz2RPVVay2innstZ0UNITZS0kxABFIG0yFqpW5qSdSmu0L
HzwegMjzKf9XdR+wV7PXTQN2UIDgyv6wrIEIS0Hm6Uovt9vDpMNaZcX3rnjUkMVuU7a1i7bekwRb
aEZKeFcAYzpI6WaAeLpUCRskl1G1R4ap/47mQijL67JP5DtZRkfX5gQfVLVtun27LUrv1dkArAFt
54Ac3Oc0Q/H3FnQMJBs/3uygA2iAbPYyBxrdnoYKMurnlTtIiDMPv9etDi3N1CA504BCD+N+nXJf
Qa9pQp8BIj3aKga+r+vUIXOid+55W3gXnbfByeXbQRbGsxLiqRuYl9xBV5V9C9Nuw70k4trXTBF4
YLpOdgw3O8nJaA5ioUDVd/Epz4Jy36A4EillekbH8WMre+r8yVFMq28OOAwHzyIV4hZd4olJgzpo
InH0kjvAEq67ZHypYwKebLK5RQx6BoooqRaEFlWNE6VyZonmSLs8paqkQn/ce8Jrrr8kiIsEClxg
8PCKZpuyOr8AlwyNKBafBX9Jdb/B3HRAzLzp3ql8a3bAiwIf892u+JmJpt5xqonMCJiip+IWAbmz
PSpq09/sSnWQqD1Jl+fJ9dKsBpqbnKC9+V+C8llnHAF466vfciHGcz9Afta5RIlGXc0L2vcMhVxY
oPlVpqjyZ3JGBR9lAvhG5o8W5sL/rnCzg8nG/nd/feI1ObL9kchHj/vRIHpkJi3/etgJuFWQu9jP
JmIvrXXz5yOQ/seXOMsa+aUC/gAyCRkNkjePc0J0cHhPn8IKI3cYZwxUD7Ts/Kvobr3t7oadYudX
rhmEzgISDk2qq541U5kjTkwN7gdsdDrSEDaQQ8Zr5DE8PqpN3F1eGDb0TDYE6hlyNP8ir4sI5twW
+dVD3eac45JD8K+Kae+lRl0UZpeKYX9r4ObFK0Yerpn8ccyVYnD1ae5r1926Npo9qx2KFeJklby2
05y/CSlo22t2sxLyO+EbtjCg9ji444U9FgEqQfNEM6w3reUXJ40H7CZQubt96j9o8HjG4J2C3e69
Y2zhNB0ZQykVEIqIoDergGC+rnV7HBAWg8G3KJhzRyKwK+mlgUbASwC6TIdkaXbi9X5qRpimwdL2
hAL1sfb2RkOKXQZWTFCQjRLqIsyMhklgMdNuacgE8El9Rh1HgLU0vo49hPme12zDxSabLkzCiUBi
l0geqpG6/Y3r35s1pBnWHrWegbeaknVGyh78MECcTD95NITboPrLThefoDNYXSiVbU8zfx55CGEt
3VysGcupbzCKxzKB5RUBLVDE+i/WJHr0VhY8+Gm5iHahh/yNd1aJN7jlQM9vaQ833DF/KFN+vmG9
y3jIycalrHxDsucIUVBAv0QWKByaCd/Hi+Htcf5U6rXL/A51M+31i3S2lQUEOskYAIeJTWe+B/J2
5wlRtkHepCqfUDyC0wUzOGG+YwtMqXnJ3XAExjKXdd35o8VXSJy5Aa1LdlWjPwgWg1HHWXF4Jr73
MtClQTBF4I0NEhm7Eowtm1ejAORUptzCalrR8Ar4MiMi/PJsWfq3szBqc7kZN+DYwwYhKRWTNs+q
9iysGpbtav4y5Vu7QL7u83MMDqxq5TsRd/mYCSrYidTlQykBwAsICQTW8CklelsHOwugfyRFzilg
ZYgVlhO99pWF8lSigUujl2hyuZJqjbCOMUHBZEeX2J7ExgOxQJYQZ/Ogcsxl2+vxupbC30rH4ysB
4gGCi0uDhcyzx1LnmfUPe+BDKC9gFg7np+lDAEaVnh+zgtNAaixqSpNNMlfGnE2rWjZI7gs9U/5u
wrnaxVorRMFQwhOwfbVOm07Xx5kh2NJjv66ZgjMcmCOMPwq4xRDWdPPsgFRl56e+KJmujsVYJysp
Oq+JQGDUQr//DGTDohuj/QKRUr91BSVDFrNIS7W8AaFCEXuTF+fEe9xCGwpjErf5hnV/9Y0fjgVk
UyLztdNNav7d5am9vVDSrxZ/MUMudj8tNxLEq+v63VAChGiOyF2vGIwbcMg+iONt3pnxIdxKW2gJ
jU3MjpUNL8CNok/hxeDW2Pych94d82haBK1x/U85WqUYF5bQL29qv8FHs0VXh1hnyixGSxo++tBm
uIoI1hi1CQ8AvDTVCxG4xPKW+KJgVpmtGAgd3aBCzMhgDCXQc6SMpvv5V3vAoiXP3k5C4tMlGwhN
SjB5Sm3G6gNbtDGXuukZFQyfTfyw0wwDpp8hLYHBTKbgQF1hLdOy+KCy1e25ecykpnb2Uo6GG0bJ
yNWM20aPowvP3dDILHOmgxMb7lka+EaxMLF2ELxfMJfYbmqS6BHcr0g0k6PqZlNmmP20p1IKu6Ej
8B807VuX+j08vGrx2x4t2oQ4h7fzwgyz8e5m6kChuh8Su0hwK9+MviKEMnc6CcNH2YWexau5auWQ
FGOEJi/np7cRYsrtC2zN+2z+6qX8Be9jQnTi/RgzwI8+Pwj2FosfL5uBXohXjue47UK4Lk1uo3xL
diE+aPsQI0ZJmQ41mk22CqCDMabA//pBvPtEFi7qj3cZ1DP81Ehb0DdR4dOOB0AaNv8q/l1KtFYp
U4GH+06nghz0Br1QNVwsD76E5DHW5uqWLLPkQc+GxEADM7EiDaa053D5O/5SdKDhsBWNbhOCSNGr
2hfH5ZA6QdJbWpwnEKykgW/Phzo8WceTSJP3Y714Rc0JoE7RYORQlMNJVi3SeOVbLIrnutTET41y
e4T8E8Ln/1JwcMiirqN/9dNv0MYIp91ZNT+TOfzW5ZoPtMO8xt911Xdn9su/qMv9BGr4EDU0DWpV
3BXBG3MQahGPFe60XWYqHRu53TVwGpmvQfyAbCcnxO0C+kAe3e1+oA7pzB8Sioq4CBKL+aH8DY34
TWmt6uVHUidD/yh17tn44ShQxs7cHbfCiJXWsdZPaDdo/3ENJ8hr7aDLO0oRquGz2i908wPjPUj0
aU61GjlEDdgip9/1V2Sh7iPTLeXpq44saGJ7pyRNWEz7y+3PoBUyvpfbVEP0O2XqiYdfKhlfrOHW
CEIZ3EBPLf66SWRbBVriUtL20uJ7wfnKO7TVVgaisSHTHZvtkx1ycLCkuFiKOTOkWJR4gCWLIUkZ
+Y19hDjZy3E2AGA1d8YqTM5Xb6rE0CGndEsLdIzFCLEUncLWq2UEabj2DqfqslI8I75HK869ucuJ
qAMZoDq87lmH4cWlDBMTiSK7aQDSsLz2CPenCxQo2864edSHc6d75m+/AD83FhHxJ46Z4wySvEHV
Ywhbxxl006PgKPRyY9/C8Rf1tq2U7U0vJJLCKcGfZy/Dfztq0IfegCqFlIoLwPYTb6D4PSka6ugx
nVFxsG5GSDXUziJH/mtoEwzsF/OJjaKZ6/ckCHOdbotb1FLT6mAjZz1WYeeudhibtTDRLvwMb790
GISvwWxCIg+UnRskehJe7vyphkB7PE1F2FPhctf6SMRSg1ikZItWuHoKYWMHkALcIQEFrsCFoHhN
dJ6pJsM5kdRy+YYSdPnr5ItXkiRGvTAxVytULJPoIb8z0+NRAA51l04SVtd6tzMh2WEiWIppGRD4
rih5LoE39YtzhMNsEXhZz3AzDpSmwr2NJfaM/VgXVSv/UBI7qLxPtXsxiOXY5FgQs6Ityvo4rVZw
0Zkqn5l2JysNfKYlKELh0Ka+uqb54qNjMPCytyyTAQJnh9CeW+kNYDrt1xK3u6BpRIU4Hxr2CXtl
F502wCMUCGtGiJTP6rGbU3oRcDRMBVZXdS3nBKn8icK7TcXavw8G9ZYMEU5bVnsFRYCDlB942FTl
syYg5+GF0vqke8+swfZTKlmYtRxtBSB73nHDivRsDpKKHeDCnAFMc9DG8MuCejWvPJD4wYgY/TCb
YNJXkoTgbUkF/Spp+svBRHd9QpeGqIqBg5Tu0se4SkZn7MG2TldGmJh1Hkh/O1U/rJA6wPVsYjtm
qUayBknCO1ClRSu5NpYV/CBGy2dTFmBdmNid6ba4r6V1UhFZxsNbos2/KiLyRUF3XI9u5m2eYVnY
lcocWjO3N+7ARVcSGf0TGkSgdjkiARY1O0WccYPfILKpY4OQcbtbPywHI3MdSrw4OZVeAoW+nbvr
JcxAoetpTJtlZVn5nTQCYV0gJaW3nTrbuR82OZsL/G/KtzltOKUU1JPITWeJVPQHeEJwFbM/SFHh
K4aTfA4A/sEJoGYjNQ5wInu8Qnojvg8a/ugaMDO2/svThfvsG6dM1QtangRUZswSCXDcFvE/Y3Jv
6gr00R1x/b2kFDbBEQyXgug7tcIqL2khqnF4ZKz/dhhE2UIDWwqQ8xIY5rA3nfNlQoetg9yWtVxv
qa2Zo1BARIZ3GADZuUqiPpg3TjrG8mbBRAOOSLvJpgnEVorJA0UTEqev/jIBVw+LMgA5r5d6n4Lu
eznU5d9yYzjcy2LdX7wQbgZiAwlIvIF17KgbqYDCabHAoZOL3RndPMVtDpPsn8OvKdylQqLPxJSt
fTAL7MYWy7l0GLdViqpNNhclg2Rynj6XFgEd5XVgl3q41tYM9MN0adWtQfXi77HuoGhCqtxlheFt
WZgh6XWxO9tGTWAM9xjzdZ1C921/85mreH11eLdUN8bwj5ieXUuqwNnvyjZcjan3rXIgZB9nHVB5
G/fyynEJ4ZarGn+nzkoyi6F/N/0hEerCHlUK+QQ3M3Erb3x7hSXES66ipQAm4FPgCb45T8FO8SKG
l9mRx4MdilRbU0FoSi5f6Sd/TJ1j57bqCIvlAQu2u9t1ta5mUmrfhNo2pBojQhygK0hS6Gsma5dG
Jk9gg4znyY6NX3niINQ9k4UPXmxeuL8Ntr+AaY4HSN14g0+KA0km7CkDPXvCIGbRr3s470LkjNp1
qHbw0h/bC3cBJwC4C1YyM1oc9aK98+nY3sfx0c3Fm87JJw8ENr5+qFF4El2GeLIPStjaXYVglvGV
xepgjrR2tZfg803qXglYMUVT70wFZr0fGWTaOSMU6K5inM34hXv3KNKsLEmLpuQhNeUotISg+OFb
jaHBe0jxFjaQqYJD9U99o/nUutNOCJ5FLhvNkccsnT3/ZRgrhOiMD6VKeIKy2KdslkTFfPpYnl6B
gDeaw/dc1fk72VV/RV0vpqjNpMmI3r8JxImdrW+bso6xQyUI6S0i7/rRPi3ainG6ew5cBkDf4LEy
8omdc0iRw7rm1ZnAf1REXJkai6afGrvYuL9lYehjnjEIUSff7bryZpDDtZhW0NxdagwxZ1tjDjCe
L7kDa93C+pgFtNNa3qg1zWOhsmiiQdFzCntHn0k3i5hxyGhWnJwhrFy+WwJw7gw0V2UypbMI66Qq
AvcoKOseLVLQX8ZpidWVpBTlRVsQ0iERKdlMThyTEnrFA1L8UNjh6qEPS0jgUMhFB6opzbyfzZa4
hINwmctr/MmWvNdOce5VQHgZnmuv2TDGOKlNwcnsXXaqVDjXz2ZePWI2Y5Xb9Jz3I/WSYGEC4nGP
cKt9w9s5dir9YGBAwrDoyD5Gir/xFt2ySXlBCc4c3vVW+m0kYCWhDLZe+P5K9fhuh9u+WZkYHQfC
TiA8G5SVi178HEcL0xk7kVh1n7rhw8+EqHna6+7mqNNoUqNoIoQZ6LjkO1JI8of7gNFe+k9sDafk
uZXVwLC5GUrdDFWRi6HVcMv3gq5o1SMys9gktNiE7icmQxS4JcMbe4nTXUeobpB4PJPHHn4nEV4y
qymQwHEHoHGovIiadx9HIATXohT0P7CvpA6Ts6D2W/p00244bJQIV/YeBYEBLfHGrSIFFRHOz+PE
54BrW4Rib2bbtYSVnUU6UszJmwwOKKCGMwY+4jxXpD0zeUkZ0kyAtCDQVYAbXDU3E5NHV/7BNXv3
R5q29u7e6SWxQe+ejIZfN0HL6TYj/vptBM8cu2Na5ZQStyZDEJNGXWB9cerVLgtxQnXHC8zfVTz5
mwzxI3jvqCHqzguMgaxkTcjmG4TVL18Vg4YZ8qTSzcj/yjONyhHGAnhhZRqlnphy56DgkPw8IAfB
ak/p+u47RvfxgU4K3lpN+9lBGPn60iFKc2374v/+P288RMnKTWoZ/dqM5h0fO6wWb+nEKyVWKw1n
TRvnOeBr5PwjzKzES4D9VKZbD6yayBBndniDs6BQj0wqyU38F16p9qY8/kRDyoFnOFrffFHk9ctg
emMU2P55lCxg7Isxv5y4F7xo0Qou3E6hOf1mmO+WbNq4c025eyCNtmeRQoJy8mFN9P0Oq9nubPFj
9aUnM2TEnc2JB7kVOhPvQz6e/fGK7Enq5zVGASky4NTdIzCYJDtsgQNAMa8VosJ4CLyleGIuhCt3
ctW7ka7HwvzGi9XsRhh10CwtDhis944IUXgpvbWn7LjOt27PWC3T1NO8Yt37+Fqp9Dl001QVJaZV
IRAJk7BRnA8ZGU/dTPJT8/RSdr6lyXvz4F4UhLEGbNAflu0TmX6LvulNZPpunkkzBUqgbrKFtsry
dskO+ykzrkKTCzimpLGJLL/+XiPJ0Qd8TtHtUzFoNMZfR2xCa/SQKRsse6NcXzVuiXvAdxrn17uy
+igYucOOntbQd7aAE4gQJAi6wMC7Gb7AXGURgUBQnX37D1CrENAykH1oy0sbpMpLJa5zhWyOoIjo
AKGXmbHe7rWWLILpXnB9nOzWZLk7ykq7indGE1rtroSNZnshI1pwd3P4mxy0ZXSOoMbeuO0Hc7tt
iYnzz1DxOuzg+gw90nuxgFIA86Fuua6ec9Ssf3r9YY0sXGgEiPJOBI9tdRRiinEZGXBiC+fhd7c0
scTsWcs0f23Z/ALQKBGYYuu+FzI09LPBsFe72YVfBNDhMaADESyTqGkS0va04xfMwIVz2o3di67/
WoKa2E3v5+qrlDFgbPIwBZARCdPld1JSSDNXMBymc/RgO3TQ/oOJ2TyakDnN6ZocS16cuzXvJYe0
VyX3D+7a5HjCVg7Z0bezRWjoCoX92QYbveSdyiXXL301eEDXi3dGSLMNpZ36vB0VzKU7evGRZ4Vc
NSUw8u56kyzxrRdRMbbhdSUNeoSmbsmdZETeZdyuOtzjMujvbNQOoW+SfPt6272Ri9Fl1nO4KIbc
WZe9PuT2dU6f1fwJ8N57vrxU87eXIQojW1p7yaJW7M+K76pm6ftxX4tcrlv3kGlqEa+Y5ZuqoyUS
ZH0ZcgwsOinBmOVdp8GH3y1cZYc4LS4sPuCx7hUsAGPIf9ra2Q4XfR4MFwggorexMltGeKwwldmM
fGqnW1b/4cB2cMNbh/uopl2V3/7/fiPJNPEyEiMe9Pd0rFiYnEPMMTnjH0k4k4I7FcWtNmApDZoq
Iw8jtVikGkdnmvYVlqgLFzNPUW05dNPXlGT6Abord4LTvmzKSiM1/xLlQAb4k6UMZjNaZiGFy6oA
jTaBb9MElNWDJwOAI2cBraPWwRDG7Z4mnhgj3SN88ajVx1RK6pMEorbtfk8Fx+BssjCdLKVDQ+Rv
3eUSdX4O+y2B444R+znTw8mdwjFhhWS0xA/69labJFHT+aiXLaO9S3HYrWGXOxLRBctq3L66CJmv
pfBZkKqw0GEXvia8OJ+Ypa+QXRA6pmwxcml4mVV0r69Glm9ASOYz/IJIw5Ap659HePbRHU+36rZE
HwdhZwocOl81lOI5tvODYnuXKTx6YVawOpf8Qh79zafmtl62k45NqnaabF4oM1ZTmJlx+0+kNaTs
be23pOqYRbIiaycViK63BlCzN86v7Pj/VzwH8tlKxyYvsngImkaVxSyXO/CWAjDGE7NhyepBgquq
iufSmqs/trCUUjzSC5pz2g77Qw7t3HVyE+4dK8442HLHgEaK2qmGEwIy5rczDSpOq0S9QRK/hYz8
5JNdFUe9qemV8WIV3LHeGX8sxN7jVEH0fkj8iSFwkiL4nCebPxcc5FZ+FOyH+fnOWkVSu3V6EXEg
Fvb4jYak3U/8Pz4jdyDb8izSPHJcxmHYftHUWNi+8uzlLwcuApJCcScHJJ1Jk9lRL1JVCVEclsvR
RLGcUr2LZy1T4+iH+wvj1BscHuZ7N4deEi4nUdVUQFZ9zSAJ5LIwILJQa+lLqneSf46f7MJgKg5D
jQbNArUz7O+IXVXTNI9tpLMf4B/h2WiTUcl6zsomOmLfyfe35pkV3NJJl8AUrXkoFgXYi8sWFfGe
LCL6HSPaHZz3Nl6zUWAvzzu+4EAcOc1hEhwXVqtZkH6ZEfzXvU6GpLVbVO1ICzRxNpzXinEdwybY
fzaFZh9G+9CxK02sqOZ+luppdu/POOc+32iT2+IwQJuXjPVJ3fhBs4zQ3xl3DDilhZXojScvzZcc
wjBQ5Ugm0/jirvWXpWbK0n7pfzhDeAXIcgYTXzKHGhKhsMKgqdWOMWsi+7FYqEUIITPoVpD6sIHj
iIa5eKUCOtYfB0WA3EekATwe+VG8Kki7ZnGjN4e8UGqFg2y/N4f0yopfTtiTXcrDa6XprYsQxYAS
dtvWY5Sebpanswb7xttnE8laeIHvEmjHI1vFzmj9zs/IW1r9xDZHesx0L0fyEOJhXKsZ5xmOkawt
6z8NFLGJuGBFM/RykB3V3+uvEdEemomJO2TNYYq3m8j7ZhrPzX8FTJPRJJNvS8mC216NExbEJnXx
ufUWA56PS2mPlojLotxHrpTi45Cle6JiVRVb/EUXGJBzaLNFxuH0+jQtbgIlvVhcWCS2s7eRToP+
ykJFaUVKYCeRrcgpGe0zp2PkaE87kv4KIzbBfTcCeYaFQ/SjZHIf6z1EhZynKIhuTHv8oLZLS8ez
Ag7xIYZQx1BYu7aI8dUnWITjxFcgU0rAjZFRvEpOi8DVMCMTOCICaHj0H6cyKD8x3XEDy3JftTT2
i3iDC84j3deuND24Sasq+rAQxKlJT2rEk9JIQmezoHNU0uBMOzDoSnqZxC279RzOOEx7Me2qJkB+
r64+zxne+ddcROYwiXLrsq8j/XlwUWfj6+gyGPubuJjcypEoZENwHZr/ozJneNI8cYuRpBhlbjgP
QQR+rw1Qewdph3jHdT7UPbs1GcolEme0b4vtmgvsokAyuRPaPCIu8Sp//9h+MmkvVhjgNEpAxLke
yDOzX28lcZZGQrQzF6yUz5su4yXl96gUv+LyPFscnWOcPcc5RYAZKKSoEFBzeN2xGFfQR6ftrate
GGONsytTe0iPrLoBSslC3HKlm28xnFv+Og9to7H5YylhCaT1UpKbnHBGI1cQFeeAHraFDEDk8uV9
kSjjZlmNEkIaccH8kxoTbnmy08luOnYmn6JKnGzQ+X17ywDZ4kWkcuVZPVrxL4CSwCTgMgWVbqvQ
9R7GOZfDYCND7xGG80HMC8YwhKBYoHGeHwmZGcBNzyMYz68goEHGB/hqfq3lhVdg0bRkuOIWsXUI
2gIkqiOwEeuWqXmVtpEYfbH5NZ82FvPOcCNmYhD55Uv9JIJ8Rrmi/nHIrpALHFTOC5R7oBZSGGpX
3n1l0Jbl6YzQwjmPfs14GNy3dejZkYIPPcsGqz2NkjY34gsE0USTKAjJJKAiv8BVn520vb5nbMPr
8Ddtrkfm6yxbPBISfI2z5lZz55EaahcyQRcX+fJNR8EorptowlXif+Mn4YtediP2LGUQaFA+S5To
GuVcVdkzJW2Wber4EdgPev7I4HeLU/xKm3KLrS3ENWui9PlC3PCQaqnGONtBRXnfgVpBFXshQ/Sq
Q8OmZT1P9VCb2KWY9pSw4GEjrMSA1TjSBZVVVzHYkY2KoOW92XKcIBPMBhlznO8p0X7aRChKP8Ry
Xz8bhJHPo4Mgn1zdEZWpkR3Y7qTJ/OH5Ph9+b8kLyeAS5OTvfHdUQG7dNTQEOdlvGfhEcxvdqJLc
83pI912JnVyA0eLAcxk7FeSWp52oxZZOvWPmg9P8IPbVosXnnTS+AtIItf0i6wbcwQmhzftDErY4
uMa0zpHBZFIH/79SM29+A07BIcLf2Jhg7Wa9yuybnjeMxa81dDe8ZwibbQ0B/CVw7TL5kYW9H0K8
aELGaSQrvbnO26QOQAphO5ojJU5DIjUG0832XccNaorItXRNipmRAIOwjjx4ZxZl8i/d2/PmDsGQ
Dptlcg4LlgPyyDKJdrrim5PNfCCnogLxHkZsTfFPVGTjB3mXaKOX6jFA7zgdhYisT/1hs0h27CJH
mRX1Q1h14wZiDq8+Z5fSjlznmS4ereGuN/a9BiuMhMwtn+46Pv2lX8dWbCW+z0ZlIZnMS2I6cDdt
CDwB9V3eecEvIKDfCLIrMwzr9zYC95SeQc/C82GH+RqPvwWmi32/5T0ZAH0bEGcOKMIauLRzC11K
7g0Ljnxe89tRO17dh2/w8Mtm3luTdlUQnNJ1OFjcK1IW9i9UzSfqQF9NcUOKyLSbSekcw9lVjutN
YwfXLkcv3dzVwkyxjZvrgsHtvhV1EWp7WiigdI2LHdbQRO8GoUeb7o4npRKlf4iXKmG0shLnhf1m
JU5NsLDFU/vmJD4/MoKt2MX43BMX3/IekTZ7ckdJQzm50pHcuZ95jhi+gnVe5P/yusnjTcX8m33K
u5R67mLmQocXOZNm6lF526DJ1RWLzELqAiOdLw5oqFOuFKdAifzA8oVTB3cOCfu4Cx0X+/bEIqng
Xahst0jKapCFgK1FdlieO6x+aAI6VT+qzdedB1Scq6ynJmth/gGfLYck+KRrWR3DjIQVieFgJ4e7
rzVl/nUh+sZoqeoY9n0IpFFGBSt/oSXLmMLuHkhywxH5R4kxKhmDJGanpdLJt0nowlvTfV62DTYF
nGpo21vX1jg0gq/b1kJTtXjDRha+nJAgJJZ2yYc3PP2Ouf45xb9k/kL+0iOmD5HHGG7UksgQXGhy
ArnE66iyX55pFnE7XvKfMzSSU+eJL+dwyPl14IFWNK24JnDZUJunDqXzFNtDl74AAvGJEuS2ikvh
hX8I/s9hnHS3GQQBwDsd7ce/xFUWas8AAFTyOvbJPprky2OE6jbFrNXX8Mgm3MKj3f23I1HG0Ync
81zfA0aMu3yCiydW1LpO5AfomwYE785lXmBVdyq2/b7VBZXRg/rhZ3OFCFan1UdbjdFA7e59h19X
jKJRUBM6ij3wp0fPH6qMNSX/jGSQz8jOCGC4mVG597jnOaPycG0Jh54yAYuf6hkZhmOdBmQ8nkc0
eXIjINR3h+CZHCRkVPwPeTveogweGcJQIQrwshT9doJp7fvEFW1T1j+XD6i7tuKSLApsMkDffdD3
cVUYEoPADmNYnDjOwn4Vw5+evqXE636eigfJnat9tpuVyXKYGN7BT9QmTqpJbIjv/iq2alLR5bKv
BBVZ65df3KqS4kaCQIGj93cBxH1L+dVZAQuMbtJblwB0SiN50mDc3aWx7Txyf1XZlKiGSkjFT63C
vHxSP/B6fDIptAuFBt0+uNwbPDLVhWtm0POuwgJLVMsiHrFnWCHpwYoeuC9coJa8wgV6XJASachp
+cX/i34NEd5TUJAoR6F0E0uJnTs7Bo8EpasXQX1SnAu7kwmckI47Jl6DUgY+lKB9oErLEOVAL8rq
pJNGDceUxd1qIxfyBwIBB3UADzL6lVWsORuY8FBAq4r3zIb9ZhFRpYGcIFCRIj+h35uyhd9KotFR
im2qCMEVlYt67JHokaoyPfYL9HWjHa2fmbKNrKf5PhINjmsa40uukTCZsIChtO41uAz4j1itPyhk
MaAFLUq8tPKP1sPhv6K1Ie616qz5AHwFZ71eR0YI09h6HojhJM2nhOJ5YssRR+rOfoYP9+Y5tq5d
uLMsmzytsFXYznHLs21+YSsZOWo2uDV3KP4FGueZ4f2hN6rIsnkPrJ4hF1hys54CbtALtMpgd8Su
XMqcbxGcI8DxOj+xHQ0DkzqchmONySdBl4zF6qQokq3qDPHjwnsQPtKfkU8a2EWkmKgjci7Fryk+
zZ8fTkTwLcKySlMSf5Buhch+Dhcq/l95yMYXS5Tpk7N0PgfG96mCDdkwO/iWAMCLGp8a+jwqW9RH
rIFQmiKk1jJ/KY17keXl/e8RO9szKZTo0jBFXow61pu/TvPRzODDTDnB3bERLtsBe5s8cyzLGl44
/AsiXkUUZS3A1WQtw1ZV7D0KSG3Aaw4BKlKeTy4R2Y7SW7LGKg9jMeox57dXQqoLNO4b/fyzoWMD
Tx9iSJuSBEAsDOAJYUMOlstbFFLm3bjOP7mDgWOVmMdDcwDDTPcXKB5z4g3vvIyfNhIUZVj9TiZN
oUhAzTS+34ITO7IOmHF+KwxpGS/7gvnvndz7lQYYaLo1aGyBDIKRQR0G9NOxNc2UAcHLhKtY6CkJ
r3AIiYigzKEB59mbwMgMr38DPcLCVdaP2nN8ahrWAeGgxbkyVCAfFdCKQh8sKbMiTiihGVhEHmeL
G7l535BneJV2ef4M0fbakfJD31piuiO5ZBY+kRHi5eDGUCjuRGIQ3NflteUg8WWinIl83c0bH8L9
mGyIZX4q+njwNHIrES7bCOm6MBTR74fPS5RF3y54mSlnu2Cd60x9o/I6Zo0bHZnX/dON4NcKWYNP
cCPz6KrRVK+N8KfZpHLYd/X/b2o6sKePRj+VInJ9iscUgyfKcRrC4wcIoVZesSlvwkJJ5QGEdLrI
+tgo1m8eHpyZGKze0sBv9p9B/76GdcB55ooK1OLxXxk5bmcHDGTQ25h7df0Npmi/lne/hi/rFNE3
+dQtvxE1KHc/1R+NzW8C5Q8d/P8CsS8vhtCSV9MZso0xMR1sRg2ZZqRLGTrIutqCl3Uf49Uq+jMe
Q3PwGcD46U/uYPK6w2GsTh0QglgypqtJTPM8uKLzhYvUxGssu+XLwBFm0qFDJVx5M3UnnP8pATH7
LB9KAIUgpep37b3YdXtU1WcCPnGVj50NeSoX2mph4FysujeyKlhM1IiOTAm0eiUXVHtxn4DS+kiF
WJGbYgP5Ztv4YGGpJKE0wkz5/pG4GmgHqXFJ0h3wJG53r0zLcl543329BpSgmM5pwIBMZ88q6Go3
lUbDcBEU4zLymMHLUPt6fP7UMEgoxQT2HiGZK7c3DNWZym69SdovPN5fdJXA+EJSrNpP45TIshmm
SMwJRgdhk7l/rhDPwfmx2njM/OWTo9tLPPyp4BGWa6Qbcv4CmMKPWGFThxkVoWwcv1gx6xHZnAOE
9TZsokKps3dVeU2dWFzfhKOdeEa892JwU2lHoVyulicQbF+SYfytj+xKV+y+9qFXRGHlXpLTmbw0
BMGXWGJso/Xp0Ixt66LgFsAOjhIS6OOq30Lz6A3mSsDWHKgMV1r04YCW9iLT8w6F6RRueULIN95K
pdYI4BjA9eHoBl6EdRrCCJF7pQ5S5JvGdUgBqBYKBlIKgbvxlVdGqrwxoiKBf6Af7jb6HDn9zeNz
EuL/Fy7LudAZYWELvxnpGYhYDBruJsdFbK2PxY0s/lHb47VtTtKofAd3C32V2ZWuzGr87B7owfPd
uiPN8wRnppD/mJTSPBWuem0jF4OtW6t93l97mMPKd3QtVOcsaWdqXE25ZAOgOZDIPtXl5wFZGcbu
TTZlWSdqOXErrJ3p+gFfzTYmAUrNM0h897CcinZjxFIJ2caraHjHKk6OHUoOhz32iCD042kmk8mm
HVnrWE4c9Q6mw09r8V96FWbdNy0h9bpV/Q6QC6RIJTeH3huzIyVKfe6Pav2Xzt3ioV+mMlnWikDk
Kv7IJCZ0/4t2OMVrUWNyGlqlvKSbggKNWOSI4vq+tHAh2pFta58sgvUKyRC8IkqSGW+1HaAgkxMY
ob7gYj7LhQRjA/bF9IEeZmtchQZBCSiRI4o5JrD+TJ+XXM0v2OSG7reLE6q7at3C6ppZ/XN0Gtvf
9kkqew2AtAhoAwLFnqwdsvOYHraZwo3POc04sAzi1dHXPywgjeYtBeh2+ZAYe6qEbb6agor7FKfd
P+93zm0WR0gaFh1RUHNDyVsS51tHvIQe74mgUIQA3LD3hupP6XGlx7GBMbe2jvLuAGuoKBpO+D5b
Re3XMrVU0iy8kQEAdj2zYw3CKyHBpuGbH4i6uVtrBUH3/NBCfB+rizYkjCneXMwwwzbN6uEsfIPc
h5h6udZl46uu37AJscz5zbVJVuFQ72hXmbM85ogy+QhRX7Onc4MeRY5cINiHsm4okvMR4e9MhIlr
h8RYYjC33lz2dCZ74l7/XoBcPgEetH03bUYyDb2LXamTdABOO04znejb/AQ5fOwgFNq/ZmIlJphW
3aZe+H0SoHpE0EEJM+2zm2uhQ3Xg0Ee5gSXeTuGaWyDrAhbkV9cIvK8SrL5OmJ+j5YjDMIlyHBBd
dpO9LZw35DZbOK/Uo6DWX1HTnz/Yk+uZMZQWcZS1m+qanoj0GRpD+w0Dr1P7uygCJGo6N5SsZLuL
QSBnBK9FYqLYs42XFsNHifM4Atc6IH2wHp3PcVlab/o30jvn9Lg8Wfef6XRV/H4yltfaoarrUOyQ
EoN8gpThEXzhP9Wm2za5bkbGJKZVtPx8KBqu6yNGA5sziEyI25Ei9Kg4HJ1siXRc+n0QJveaN0xn
qw9JrWKyip6dOsAu5cGUciu/l5qgu6Gp3HRWbhqXd0CJPtXxsETLBk/UUHbXH6AxJSOIMsCZEwYC
MWsvSE6gmWfRvnTueM41Ns3XksJVmPYahI6/zUUbXQyowxtdVCz9Fww6ygOLEtCXqNN0XZAAUXMa
8U4zO6+H15PRhxRYAzkzE9xVnWuZjgZSQd4DohFpf6jCB5CwcEoUdAyOr458h4I9YRukbUQF8YvG
Ludr4j10e+g5j8gUSJDmvT7Pbp5QEfsB+8BzbB3dndAyONtzn7sVlwim+1cahtqVyj7uMIPtiNdf
pWR5AFQ3S/n7L7lPNGCWiejIOyUAx+G8FdHIWmK6eEd0UORR7jLu2pG7OG3HKFZSkqfzxV3w0EHr
BomP6Nkf2lHGCAsVpS6+D7j+Rwl8Mmtc2hTtjSBe+FX6sumisoCfmEzX3yLTqTpXDI6PYVuMUY1c
/1m97Z4R1Tt4xvdtTsCeAWAhu0AraD+jKLUmtrmMBGZ93anUNkK+f6HH2CBtLY5qvES7fsyOIBdg
JifbPOYTq9KNejQOynM1JbpwH3HeABHkogCsJEgOSM8e/CL55p3HkCWdvf4S7OMoza3dTr6qes7f
LNNFAE2Q+3+lSZSVMbk3O1YVe5xPruKLCg5G8lRiQ4cwy/IEeZqOg3wDjI1exydJ1Jymokdo1XAn
k5avKSXwxFv7wX9x5+tx9iGWC0AB7UcqAoeFvZCIie+lMVnnJIkoedovKeIhcCJ9JL3ODzHkfDRE
W93jpZJ7epTTr9U37qfxT897JFrXKxDS59za50wF0MO2aVadZhm8G7B4KqGhkiVU/+asx0Q4dVv0
EqdMgxK/kQPgQYUxyuHMK3fu9fOKMZvPVJhxxqVVDy/qUnajMkRbsmcyKugOV2kuUkdybZuFZKrz
3S3cxkkQo2uceTJQHDcOz188LZEmXM6Lox+Bua/7d3vpDOymNnGffFoeInPdM3/YX+yvF3poUeUz
N3DuYG8+jopIbP2nKNhlNdWGcx3xqb37+LNGRg83tJiRjt8Xp//L4OamU0Ai/Eq5vsp2FddcvR6P
Lfxyu+PdTBr3Z1ZveLQ4d3N8jq1t6MZQ8jXxi7nS7+2Gzc4P3LKYyOS57u5wz0TlEm3c0gN3+il7
NhkLU0V/yvVEj9R5J7CdTHI6iQ/j1E4i38+kogAV1vee20ZoP3+v2wY34LPxmjhkSWFxzF9L3+Yw
S4h7zpNNQVV/C2wTpjbsLrp9rZBgcBfxU3NOcLTemd3E+ie/GX6jNBGnjPRdJ4cHdQZww2JhZt7Z
H27wGqlZDbio1fAQyfykpPT68nUHd+bOfQ+9DDviMwfV+U380Qhvl6DnXVn75b3oX+17Ei06YEE7
oonWA6x5sk5lukV8eq1UvsSStmY3Ro+/QwetHnggBez5I0ywHpzglHj6eSMbmvZqruMoGB0YoEBl
yqiWxaz0l4psjOtERACsdqlPzjP2GBPMjB4TbNSNibsckOlybCLr8wjO6c97fCqCbmoA3TzB7u4r
7btS5vz7zTe04zD8YYizIsGdAIeyK10lF4L/e3eoaDTAVbT3NWGmtyoNQEnRONkgb/o6wqTamN+X
Kk9L5GQhm9i1cOkXIWNcZ5YU4nAevVYGUaGn99XgnXqZLfdgfkW7eTkUGhP+t46xT2QzltYtUvtM
UgJ48PwUmfW6Do0k46pycDt/c9HR+AZ8qSTCDuA7SMbvSWGt1MV5SYP4qD2tgztejfrO88cili6H
UWEnMf62fMTblULLm5g2IwVjYVUHvypVGAnM5OmSA7Mu77miNCUwFA/H0bDlNIQ+cipS7mI67Ccv
jlD8/ScW/fqOESVunlWMCyrpVlbD2pRCz6dPvX2nKR/faauJPYyKil3avEH9NGyhBHz/iYxy3RBf
KATGprFYIsFW5/cLUIXXBHFXUfbxmWZ5wKrY9MEUwJ0Sz/MJmNzm6zZM4Vp4TPAeOYBvZE/mFhkD
gBrOqJzTnrNig3QICOLGbt1C4fpHmdWHFp3SYdffDkR2E7CBev1OmNUE9C5xUnru8SGrZ7KXGpKB
HwDoo0AwuFMQXdD7z85iDj7CN47QSR2XMaDcDcU/BHrvn8n+H90L4prVWbsyrrwAphFJik+hk510
o4HZqkBh0VZ6GyEtR9Rx4s2aS/VzXEm9fzuWWpdPJg7kAXfzwUV3jHRFGx2gx9qakHE6R/d8KBfG
9bbBUZJPseLPrUtaauDtI7V9yDq7NTaTaSYPUeYC0keunaZRwGAfJ4v2FZuNwsP9UU2/UkM7RTUL
yamK6HtZT2PAkz3nwJnaDqxmQ/+Tv8x/QBzXKcAu4t+sQlWKkwaKLzi2MZjmOqmjx34dEazVAkn+
iYMg86oraKDLZ4p1XFWQJ4Ssx/x0lpDk5BCUNIixr/pMPRW85jF9pCrU2R4Px/oefPhmPZ9Jpn1z
7gsiWuOHerzdEGEaqI3qojoVl3Vk7iDPDPigwZoJqk03+slk8/z1faLVF4FXWXSCcZga/B4dEaXm
Dj0OYAzeQ1rbslJPNnN3KcfKwva7+K4oW0iP28JjxpyCBrcHk0vEYYrWr59ZNscTpR6NXFqfDkO3
8y4+5k+fp8Ubxn6hA6Ux1o6lPIbH8Z/bSinWpW+U3r/dr3ilG6UAvpiBuXOvrRqCB2lMtmcoG+FT
CV0DYmC45w375IBW2VrkremEbofwHrOIC59k66Blk42juU7B/7N9BfffFrn25z8ogS0aIFdA0Oss
idU3KN1L8mmW8Jovz92Auxl0HnfOtSXmNJ0ZJgF3QVze5eoAmzJ2Qxp7pgm+xby6/bvWPojTpkR0
YFYiIW66b2OCOqTL4M8QZ4R+4jwX1D0p1yy0gyxSsY88cPrAeIE3Hk03jpIZkruOFHaK11BA2K3g
2Og8mc3IIVjH56vdBsVwKew00UqQWIfwQQjFF8b73pJg8d1xnmPN7VeaYZEJNs6Yy/7fVW+RTBmE
m96yEgubNpKCGJ9OfXyL+Kib7eHfMPLHnmMnx8VkBWLk28gGXW5AsDLL+w3MH5ww4/9QIRVgVd/y
GqhWHtjKB5WNvugZmVHB1XZHYUs/8Rxfd0fVJMg9f45kGbaMzkh6GxeGfVpgIL/RPP1rhU9u3NnJ
0xNSVWE32o2f4xVdBekGBnWYZnc5zPmuez5UQRRw/SjeR4Mc0ND14GlxLWcmoA==
`pragma protect end_protected
