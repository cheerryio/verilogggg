`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94032)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCbd/xufmegFFN7ofJ3JnOOHp4xf4+yzvoy2wwiilC1g6jDAa4d8V83PJ
Zsq8kDORpRx9Tpabv6inbu2SzuFa7msufT16+UmPonZT3aB16U/GOkTXY4KWDHnQIKEX9cPAIPr8
omu8oPWgSjIRoIXfI9eQnhGHoaY5gNtXeuAFsPOd8L0SbVSkh/lazRjcl9FFZDVbLdMOXmo6aEC8
SbHDFjBwdnGDjVmvbLFNZHlYo2+qfAmzQxjCDtHeRKYgacof9Q3r2t8vlgJ8CDDAL9kqnxOZ6fMF
27Rq7edba913wfO5arcQ22jareL5lpb5YaqGHRYjxgBGmTd3YhSQRVGOCSHKgU5UtY2NjtS8QEsG
zfTb0I3nUeHgiWeeBSSPabNqRu++QoMdO2L/1jpKm9ZI60cC3lSNhxlc/1RyvdYJF/bLj3FTjs3M
lNdj/Y7dX2S/XSYo60WnCQITThMSzqmsdT0BQvL8iA2dzbVIP/jB5j/AelhgtT4qd16dX9MesN9S
HxQft4sj57fiNGO1j/YbQYAYVIHy6puo6rn6W6oMYlZYBwwZ7Ab1s7tY0npwknWuqydDS+PHL+l/
H9wBP8FVHek7qh+7lpiW5hWFBRsgOTZ9GDuUhWMoNt130Ktk7n9hKagF6o875pVPD/svMvdzNmyx
x9TtcxRq+eKGDbFoRIpvlhCbfdDvD//vqq6Xviz7GDPWT/T4ZViTbuzXVNsdOtClTxA/lSfyqkbI
mdRaSZjobPjeOXHx4PRMcRapqHCKKKVAH8LKYi5V7Sa3cSgKRYdQxtzw4j+zROyAQ9MBm4f3xtr/
ntoVdt+tkK4TYGPxyHW/1jPQVgZflZlnzpzEwjyW58LHSPAZaNuEJUirWFWGFp632MXx6V0fV4EZ
DbGbkuL9643sRqyUwRgJkDM4gc+KCmYPKQak9lswwMJPJau/rE5JGIPm0qC/7t/yMgFwvHsEsNyG
EhZfC+lHNnJyNUUBlf3UPhC1UwJcsXUwSwogvFqEIncBr+bI1U1RvMB57/3HwbuFHW2KgLOvKys1
x8Igww5YASC204ujA2i5MPLqR0qcOwOAiCkU96QcWVgSyDEAjjsz0OwAGQy+vy04kowS27qIPDht
rUO4IgysrahjbxgpI4PoWZY1PCukOsRD6eHpx+yhSt5/gocPt8HNJKm2R0DmyNDBgmp6uphnqCBs
quJiocm1L+imcQdPdPdGy26wxw5o9kG7AlnrYTwWI099wG4aNC5L7ly/cth7/TPMqfKmE6TuxwqU
U4qbvL0I2FsEgyE3iqDYxCL9wv43dXdQX/QJMKbIVE5O6p19zSCvMknKMTJHTkV06AYVMs2sVTYM
kRYePmLe7VK8HwuxD5qX8V+zX5kXzaTeSF1mgReplmM66ucZOIFEX9g/5V+mw3jrVbH/Xyy00er5
c4v3zTv9Uvsrw5sTh9zbcNeeV9S69Vg2lp1Owa2R8XmR+FkhiZFMk2PX60vNCpx7EgFhr1r4mkNn
gLgfg9mRFgbvUgEEfxhrAtFUT4fKvPRl4fK9xl+ZPwSB2TWt0bpkxwWrTWg8Mis7qho4685BdsUM
iKSo8pnkTITI/c3LUWVozl96gPl3huPR0qvLDDbXqFguUOKxcSD354wGSHj67w2THc9BDGxK2o8u
WZdcS5c+lcjiHl+emJ4VzIFwMRL0m/U7tUs32ySyPGhDpM+yoFU1WTr6AWQTpX2g1/J1wRAHKXjM
nQy/5h/uHc1QszyU4LJFjX1CAK8UWgq0hGq7x+eP/ghjet8ZlAF17RNM05uAQcToaRERt3INmTDZ
xSzYHlKrmLiYbcVN2AvCH/2q4tT07vdQZPx/ofUIDohhRMM7diXKnVLaZ3RqJ6FaSZle8Fw8q5NI
oD6CYC8qj1cpH82s9zZQYzIJIjpXjxmEndLTTJ8otrO1GZIU9+NEZcjrwhFSNsp/tSPs17xFFhRE
6xxKs9YFC4sa10S7A8SIy67zWD++LhoU5DnyMrIv2zwGaygC25Ixc6PWa5DYDJXrL3EKWQcfHfZe
HmYmTW6TT5boluMOQWGhZ3xzKVnObspQfAB/Wp27DO7OVgPj37duZyPKbzc9nich8+YcN0eQOvcT
LMZVUfrAlHa3qYpzAz1DTaDPGAO2UgRop/E927MJGqn058krxUG7rrpiWrKY6OHKHhqjdq04vP+R
FIEoIZq9pMD6ZwKIJPbKKIx1bW8IR740WjTB5ZxlnBi4EyY6zvS+KAhMy1aR6dLrjqWgfk2LABFo
FQaI3wAlF/Vt6D336kbpzK57OjeXoVYJv9mhDETgchDOYKwiaK0McFKZ5hCNhMsL0xQ1rwEsspps
e2iL6e7FQ6VZ5owOY/E4CZD7TaqSxkT9VczVCFcmefkIjWr3rW3v01/cQHWI/a9PeNO1VXqsAZud
Jr6/bf7kbKhsnM8jj3ruxb6c6ewW6+vXng0BAzvoS/QPX+62olLFmBAHS3zHhCoNKiWud21x1Plh
pbN7vUbn3bMKxGFZQYSy0nnbWyEOu7SHXSchqTY6lERnSvOPjVBUhmrIQ8q+4oaHMG6fKwJacuvl
t7Mb/X4/NGP0Jp6y974h2GhoB3bp43QFg9OMdwTUMThoEHjBqzMrZR+QJwV+0Sdqqoz+W7wg3vws
NasTUBZ8gv6TIYuNqhsUElB4EAYNuljS8IHmUd8DpI6Fh7PoZXkBgM/t1gVyppNSBfNF8LRxm1uy
uCCayq7SPkns3teSrUBWKXf5gADXRWDafgnwTlAsAR1OgkpPmlcNm3cwYZAknnPKVy3RlX7Z4c48
eTLJp9KyQiR1YzfMIEQNhfPT8/Ss+40VStrmAEwCPstCaZaTbU8ZaHKlD3fpq+3OGvQRzFZAaQjo
o0SFvJThHOlV74RFWX0DcB1CcHTWUIMhyP7XpuxJuBeqAt6F6vKsPxPbgnlB6Fn9C7+Y13przGK2
BKnzgldEtgCxDLbfBnubCYnyP9tQrLgFg9oZ8D2vNPclN+8MjMlv7hCRi8L2Y5jWDp9kCjHENRxk
gIpkRErGweahSQ0Xbsv/9veEEGqPohFqk1+69b2t8sGfs7l62eVy9ztaphHshdMEBX8V55GzmKPE
cr/UBKEFJBJrcb7jbu9erSTcf8NCQ4iG2m/Z1fPzJ11ku3jBnblH6Tmgg98BtOZbgbvApxqTlA87
jgzIizNS5N554/vR2UFkN1GjAMHNU5UFNrQzaMDG79UWfynTm74OxmEou4W9pBDNvvrznk3Wgv2/
pDRpZa37cQkJXODkqrk3vx0ptSOjAlmy/KeU4u2USMe0OCwgrNfeWiwZOAGZaNjvPvr7Omucp2T3
eKa5Wx/5r02GlclmPpBk1+M3PQnmxkl/6jup6U1o2ZcI1avROO1WBPI5oqx71Xbugtzm8K4dmRjG
mIeXHBl5nPFyNhYXkqJiHOLzUYf7xX+N4rorXMjTfLpnh/j7BL1meJCPz2cNLcjQDWxRfUFrsQQ6
VsUlpiwX8TUo1D6ciQ0JoKhYOCd0uRPQPsTVedPU4dkTu9GXww8RzhEQOBxxodpdV0pP5jQ7uU1Z
5CNdJL972tPBb4N1N0SHVFDz9+ZS6vcFRzRm5b8S6DxA5YGPchANlOANes9Cvc1nXW56c84apND1
iylZG3fTwlq/yfCUOSlA2+MKNmW8UUON3/z3MH0F66my5Cb4Yf9yhLgby+rjSmDeAjH2R0rl6Ytn
AURgf4OkcdeMI8CV3SJ0eDIog8eIpKqpLgWN/mBveA7kAG6EfFjvc5IAgrc2JaNNwAjxzFT/fM2V
+4EmP+bCzOJZbPPMwgvgoUsvqXvvEcC4fQHjEy8VN9wb9SGegX+/L8isBDqvF12lR2dZjj6KtWau
LMvYCc/WTE+TfQxFb6ZODo8tlEXdb7sFkFqAwWSGGDlwtI/g9MY5Rzh0rbCfwferb9uEN4Vhn0eI
N65pjJQF/yChalRpcfzsqEltv/sXcT5iuB97tPTvS3C68KWz/i+wsG7ofhPqMweikeOU44+1A9Uo
Gji/k39miPW2mjOZ6f6uWirkz9dQL7QDA/Vp0ZxOw8a1UwhY5n1v4zKLuAtsD5zgpPf6FbLzg0pa
uI6OBOq7RGwQj91rMUImlgw4CNAx9vlMFAoJo6Faejb9k71VeO7Lul6gV4UdYKH6AB79Zq4WvseH
07GUDbybLmWSxiKIgeAr1BUvaVVtEuyVJbgiiFhiIBj5ExG83HO3dIoAlBTBycvSRC2y4SBnVLwb
bhgPeeZhbZC1uW3lJu74rzWpviahW2RjKKpLxUAdvkMks5dgHrkblhnrHpQWEZb7TOfUD7XVr7Dq
Jk5AHAPnm8Z1ckQTWM2MiRfE58D3/5XXv0Y36zvAazl6CpYMxGHCDz+Ypye6SSMsW2HzY1V3zKIk
Acm4LnmzM6M/ebsh80DFSzUqOlOsUOVOb2Q/qOrQu8CiK78L2ZlREsH/1omIcmwfhgS/4Yr5zgSf
9z/iQrUR7NejkN+oDkk3NMNCfg5nFDrkrO7nh9QIr9KOCtgKNw1J9wcR/8Ga2gt0pcl42ITJ0sFO
5u1fq9XWULx+q1s5zmF4j7BQsd4IvccWgx3BJ4x3jiJTUyLp+ixsFPwh4INc7b5wd/OrAZ/02VnR
nt7gwLhDO5eU8S4qjD1Vkkh//PpdAVcgxlFqdx5tfkVpBY7HDMjPLhb4229qW3OA90DtUlp712UR
tLvccq74hkYopDDkXmKl63S9XFnMzaLWVgxqvkj5JxTcpOurwPzGaIYU5v/gDy5+PCeXkSOywWbK
pICK6beXdRGyGd8di2N/cGNoxsCMOP4DMXgC6Q85txtHDyyhuUhCb3Wsy0gT3wT2nBaULA+LbazQ
2ayNeknKkNBmHWog7CpIulZJu4QgGxQO4GdfZWnCzP6zlXUgmfqcl4ytyMwot2fFu0avrq7ctBUS
BSGHzedugd7QTJWECYMAqQZr5hMmBKFMFxJWwaDHi5gvhVQnxX3uGPisGzs/rYYeOXRykcr9anPH
gJBVfipOs0/Qqa+B3yVjUnlND7S2VIvMHpdovTQr054TJsRZgsrQZRPQjCC6eo+D6hEhjYV5A1lX
81ei+nBk7NWEyymYqdqj6fExGhtmtOaNnokyxWO93Ywi79Ghdlg5EsJX32d5oTdF8sKYn5XbSWZi
N36PnqpfavTNfONuwqic5lR59cXWu7eBUS3GzFwGNsuAYqOcSFQoINZMcV+kSh7Ns8tvmeKj9Zd8
jy6vlIVfOEZQ6nepBBUNIC9qYuN9jQubUTJPG2GzTw03GKC1az+G+C9H3yyVkeqtpjKAcIZkUkqP
9NXdSjwlcQzF8tKRNhTCKZvRnKKLWux+Zm+R2FGeM2+n9xK20I1YrsEE0fNPCSxhOoq3tC9uqQJs
5IqX+LnK9dT4zol1r0e/kglWypgFYLoahIUKwsm45oS+yK3A3O5RMGE2tGn6du24hu5UnrGbxjwH
MtMurd6mt4V3LEgEAUn1OO6nWPfYWDo/VUeL8u3WcE+WHAY0CRlZRLk67KHXDpSxb8uFy1WKJMOQ
9/lyWQIuA485RptNMv5lgMVuvq/w24KeQiUVfSooUVek/ToWrHH+JP/WQULdY0YtDDBYsRa9HfZS
44BhQ3AYJhGEEYgD+hwylcNdsJb954cq6fDwvkZRM+ncsQZIK8+rmmYCIwYRQI4gKoYdb2TV2lAm
cfoQyfXG0Bbz63YhwlGOX95Gq9Y70hnVvBSGd7J6qIGGE0RiDQk/WHryZGGd+YI9bevC9xSX3kEf
ceKNWLXjxWZ7pDXq2K2sHPXIbkiHZsPgI/StZ+HDEHUkM69ivpTOUYOTSRLuDsZnz7z3wRwVb5Eu
EXr0WxlGo23VW4Wrs0efKjRtd8L3J7xUkd/tptL0v5zAxx72MwJQeeDG/xUXYFfjaWKx3hsIEc+S
HzOsM7cGN4Ib+9XEKmxb6CSSIgayW0lYF1l7pIZimGCXZnNWuj32zToXjYbo2v1WoWacK7xvaV+W
r/deQNvr0TrSjcJ7jwPPmKOKngQDeOG8eTBBrHKWu2dvcxDLHlYsD8wwLlbJsmubXjS8dWfTaYvD
JPH/X2qhtrrv+8FvyJtXPCFTHU/4c7yfnW57hMiQRxxG14nRjYK9yUlVwbqtg/54yvIWe+vEVobX
w2ajuwsvIFwE3I4QyqPICHFDpo9M+DDSwe/rQi252aJ69TKzskIViHI6QKzYnYD71PN9QMomN2Hy
N+UYvVYiUL6tvg9MknX0yQkd98WC5Re59PRjlU2UkVDQtmBj4jOGqsETRlfbN5w0G05gV0a/p6Bh
3Aeo9ryMu/FQRslSdnKof+NSqFpVCFAlKyGMe12SLb7QNGB8gwB0IegcxBaLoiwmzjgVEiq7fyML
xMQUbgIc+lF/qxn2wTCzfd+bK/UEYIorazAoLW9AYAT7uQKJsCKcBQk7pjBTaVMS1T0fhuyLPdUP
t5Xh03LX4CZ5MMaZiVRIJv8r9OXRablPwVgF4g9pBKqowIH25Nwf+pzvYkMsFf4Y9wri0NEVPLRl
Kit3lachWslq0JdFG2BS7Aelzo58mvFpmWuDnQwc7fC8wMszbHv4lfQmX98cn+4FiDwmP9m4Dt31
G6436MnI93bzN2PjedaYg0xinsZrBdTBMrCv1tCCtHJ2Sb1Hrsgw10c614JdYqxqjTxRXRen82fb
OY+c//jwrbpll5sHNgcCWpWENCxhrqo/rXyxFquX0UKgLVWLXwn97ZZa9/Gs2SxjMBDDV4+oydil
IIUueE8nLcoK7dDGF7mcSRkpi9a8VHKmkd90V5IwZRcD5DwNlNXcTeH7vlcJv/PTZG7bUgS5sb+B
Z+3yeqE1cp8VyGUYEyn8b4Et5Z5m1t01rd92QQuonrdDOHhDRDdRyuV67eqRZ4Rdsswcm6MCos2k
f/qwaz3w1QV8Jg8eebcn/+sWqum3V3pEQ5TNc77Y1SWYs8BXQtQRsC7zENVX2aop4FeMHW7yZEgT
UlGmE0RMYoU2iZwGRiwpy3dLvAekFXrrzFdaztFRjTKLcqrjryOPH9HnwAjyuhl3zOaz3uFGZUFY
aPqFBTH6pTwvEK+T4DKdcoQrLTybVdBmI4zLkKQV3nVeq2PpRr3eBpgb+ad2bF1FKE1X5VzLLnek
fX1TmKDRbyHT6vXrR/uVW6dmWlLHPJgRdeEgwfn3Bj6/Xy1GhEbxOjlmID27/wboTe9qqAEoh/+d
SKbzg/f4yg73bqWPgAl93Cg5RwfLZ9ZVALa/v9GbK14B5f+xhgYA6MwgdDSZIO6aIjTrxSZhXTvi
dxjICGN3xW+m8VaH2nUU8D95tj4mCDshTBA885/8DyEyJYQpqs/0VaEnmDrE+/F3bOsgfJE66fvu
aNiagZiIC7RL9/T4EwwqAL6CGMgTB1o2B1EwpVs4ljfUZcnJyM+pNkZSDqp8pSiJ8iDvdNhr0lMB
R1mEoYct6s24FlQGb7Z6SXmpwWzwZbmds8jvdXXQPX7J6n0eCVoZv+BgGL8zL5kd5z9WjCAQJwcb
XL+WZa9JfM0KUd+yb5/lpP2dla+yuUTBSBy6Vx3d1W5JXztDWJ6tX64M4X40FEREZG1AOVr68H1c
Yz9zDBmKjE6AcCMPi86ZNAAGRDSvd8owMnKzG6CKE6YlQlM0aSKKqzGggn5/8hJbKhDLbgeWumGT
WWFOhTirddP5zE2TNZQSUg2EmPxNILhFHtjqUJah+L7JiXMvXib50UhFXSw3a0G2Y9Gy0arK6IJF
exqKTH2+/92u9z8nNtXIlPLP26pUPzq0emYgOeY0FegEhr7J+srZ9QZXnXGMDfEJhVdV0CFyvHSB
vL9ZPzApRS7oxbliRe7q3K0k74uDUzZLmwN5h2RuXi5fzNNmITJ+13sGlTcdR70ByF+4MPGGuBHJ
PJ31hntN2y77QuaZ5cq/9ClLSHIztYtQCwYNtHIP44baaomC2lJ0agdFbS7W8KRfEVIRwJVFGeOh
HbjGRhgSWQ+MkjVssOEuxL36NS+NyUqOJSu6rdU5KdGlMSmr7jrkdA70qfXGyBjoCY7cWfZb9svx
A3UMBD/EHX3WH45xFg4dgWGwA73NcH8/f263ds0X0stLYi56hZqVW+s5qWr9XqlYYCAQjKmcyyZS
mE6NVuG3fQo2QKcUCNFbbp6H6iAotbRVyOml2vJb54l1yiNhshh9/DnSLN/FFBFhVPCACagRXAft
h8TeuNrF2nLXbo4W/k+U699VgN6XLUPZt5bv5zPDkzAzm5da2+LA6544QW36CazktZTM5O9GEiKI
/cOSogx6ga0Ze9woR2ABnT1rfODbZxY/YFXye6/Kk7uhxVWDRBRJbJS3Ya8UNtYs4a6pSqz0cRt+
2BrWB2s19tGq72sGLrfByNIQVOftiLE7GuQamGYeetcRLEkUf9MFZXfcdxU6LS+WNZvPogHixycE
C8wbN3TCqt2VVHejBehkJwMtFZsYJ5BMTG3igSukAK4uoIN2xqzzQYni7Ck9CKgMS4FXs1uS7pQJ
qHBCPFYKfk27eCciifROuXtZJNrwaSLBlNK7WCzG9ArHyHLlQrlxpqMIhktGzoKjTZ9xaEBryBkf
4ZtdRljboW0EdxsRtYurbiDaBbFCr65KkKPLjQp7+HWyaqjvKep2tcMACKncV0fltwNAXn/qG3PC
4xjuXJbzXw8cTgSVXxhY7rN0vg6+z8DE7bDGBU91mm2zwkqSYbscr7O/Au9QpC8Lsz69eeph6z9Z
tVo+64GftywvUNdgjIycziO5WdGBmrrxcna0nQgMaEyxThFvkuRVpLXlDyZciibWeNVkqMrukz+V
v+HknsQpwj1TIV6Q/R/6RG8+BfWwRV2eDed+lNk8gUm4umCXrPMYjstSw5PTv9evJ9AKTJx19Xf9
KYBYU3C5nsXIvoT2RFyOVSFpnzZ74TcYHp5/QGbBgcULr//MfOyMxnJJnAWv49d3vnoDWN3WnZr6
W75IesejDuMe37aOW3EidzezVbMqUco+yI9rioE0FWFyq5HM+k+IAPKYn7/PFcQPM7PQRXdqf0bc
nNhmYCgD5WriUQa39wRV/hqserOz4hgfUn2nTiAKjUZ9r39mubD31z3DczY82RGPYnDhS2gw0TAG
VGNmttiIQ0oKuRxDQRr4pjTMoLuglStcIG78w12FBgv3nugEPkVtV8Zx5Rpg69sZow5HgLOZRH4O
BXZKwtdHmOKwt6FgaddU1NpT8xXBDSb8Yjs+sYLUwXdbVVtJJaPIXX1ZnRSth9cOsh6rgCu2Lipj
yRo4acs5Lu6YY+6N4FQUdBBiW2nBmQ9zEyvpwCcrVPuzXS8OeeN7UERzb6Gql//xrJI7hl3FHMcy
cePw0STbMR3OTiuzk7lkTPwwwGVtlQIByc2dEjv2WcTo2hylEq4qZ+l3hH71iq7ZJU6aqjwgh4pG
BYeCEraX63GTNkjw5NG4x/yVieMjYKYuYeuL63VuR2H5FLAq7MgDJTtNDlqFVTuxlk9bIHFySvft
3A3mGV4yA0V+32LDazBGa9o1iaNqUfFb2pYkU/euppF3VjdUinqP23HBwc7HKSp2Azju8cdOezYU
Gctxh4ie9Lxe+sGCFW/mFU8BprbX0tXhVZsRH5BVYSWG/+GJFzQI2W6ls9Pq/T0xEWwMSZxfhOis
QLnkV6XUMoYzL/ezPxaQw8WOaxCcZkQJBTD1Z7phfOHTDdzccHDyHw5VoeNFS2Ybw0V3QMsl9mWb
VBLXCsVBQC2ThPA7JU4fwQFPHotlBNhSPlbLxNqAxsY/TVzfr6nEfwusTbuH8G7zU4Mk2muHjn6z
rtVb2DVyiubsPsnZ8W2RV4mppL0TpGC8wJjqDLm6pRmTBmDAVFun20xQV1UXwlrGeWOTzMECaOxD
A9lIArW3q/f5QXFgeqYPmDA2BJTofKxjFOGAaebnrN9M2AWDTRkxEpDuce8zohYbCTfTSBxI4CDN
D7kJuC0hsKcJYKME+QlPMWvS1iXOxZIPRVEpR1CVVFBSF9Ux9dJonmn2izX1Lf/fv7oE0LRV1PGy
YkPsaGgKJlhI7pZZSQh9od4GRYxbWuBuRYQfDXuud+wYXhWIfpfkYB4JWphsEErUYIT5orjnKlsN
3p3uWXeTilwWAKbFv4ZSY+KENwi0zbttepmRd+ZtsMr/50zGEeLADbnsmhrt//cIjeF4T/YHxbHK
ECKPpTd1qpqmpj9qzqVcd3QLEyIQcRSWMs9LHN5Y1poO4do4sGMQKeEr6Oa/PObqL4KfqyUKZhwf
Ww5P54iyVKaXEcWCdzHoe7Euz38k2UGgyNuvTn7kUzwPSNGWGDITEjNYdmQeVBgFbaakqIFrWFyY
qPRmdVg6M4jdTL8TgL+M3/8EgfytqHsRFCwkMUe2wuN7PuX+gt/n5IUP2XMv7vCe9KVOvXyvyhLK
JmJ59w4+e4wv0bYi26CHeUj/t3RSdQsfyHjViI0TH1sSOj0Mb4E1CvUlQwL3PrMDzE1eESBdj5vp
qBznFLRtUMgRODtM6sBfbb4+ZPabj2xtUCORSsL+bfN76WYsHaP2Rqugyi1LPvuj8tFwhm7CsYzN
bZyENEttK6UDj38rPT869crTqDMYCpjK5oMVTXsNed3Dgz+No7jmF/Tz2sytSPw8N5E9rwuGvKu5
0A+wS4Id9O1L4pp78SiLKq+7lD4ZEDbN1gREvLENCayt6jV0eOOSpkBVlC6k5uEXbsQ2szI5Gv9M
Ie8QFiZBRODovmh9FZoS1lPXO1juYkfGzTdtIOpqYTKqrU7BDOYjxm02humtD/DY9DVSa5fu/9WA
StZoIMI3aOnEXWARRcGHEuIIn4er2u6nZpBzhjBzwEoLkA/oN/T3JK/O2KfTYUpak53CCDDinWP7
dfiqi6Jvqm06MG61ZT6XAp1dMRqF2TWm/z9TmBIVyh0bQ7wI8cpVNNOE0kXzNc6vJuHS1xbFMOLP
8vXRFxqZON0OI6SfXPzL4LrKIAcYTVOgFhWzb2VeSkvxsD6d/ytRebVIMCOVl2ZkSP94c1fQpN1R
WWicL1zUYuncHQeRLHF/n55WXmHHWxOFaXaXF4ZiTF1nNZLtu+9tJvRIFY38s2F2ZZVp+kGgYoxi
Qlx7e19tXL+d7EsQNkNd5ivbSvh6Fsxy8aYvS+wPVZrizqJRgTJGGkuaaybdVnKdH24Xlp4TDOKP
txZlWjq5uvbnPMdpxHrVygD2Uhx/K5OB0ZAP7gDFQx8Vb7ZqSfHkmpi0J0nTfWFnUxHX2HBUHylk
YjbROhd8i2a8RZZ41GpB22hhBKrwnzQwW0oLHtF+2OLkiIg2fJYgd+gVfP2YwjT037ftl3W3+byT
EeoNKzUTx3KjGWQpljB3xTVPZh4Ldb/y3QQFfdOtubeoFZviqJdpsyIXQmqV9QrJaAkbYPTGMpg+
NHs9kVZ84g4VARl3z6fLxi49AHjV7TWNc7otuEAQ/Bear+UdlOOtgXpne//Ijh/8Ovo9s1VOhakn
Zl6eEhhRjoW92Um3K3I+q9rHn5Oc101x7wyfgBR6NcuJLFzJDrs6Awixa7oWhHeTcCN2StfxeEsc
giNZxSOlmKTYrCgOKhSvwp97jq1IUkPlU/byY6+FdcktJH49F7I5UHiw7uO6iUKWrcDKQ0ePf72M
RDeOEOVe/XxIJjclZI/bxTsnhucKQ1zPDD1DT7/+/kFr8mjF34l/cWGQ0SeWSLEiFDxRw6ggBndA
mcW2wl5LLBM5pjfs4xUjzxXYEIoV82iuXOWpNBmkZAFr0prrK4RSWzmsnG2AezaCgstimFmMmvIe
7PEDOBRC1+3HuyKLb3umaIsPD8XHnWEVtN3AQObsRX+i5QaPKO9yJYat1l3xPiMGHeWEEXpaIAXI
aun+thtFm7R1VuWG+lTjQl9U2NwjTaH4didE5IPmTCNQzPs52hOnC6rscWlUlZeizrUGFNeEaSgN
dPJBaSuYqp4VYAYDwgPaWJEWMEdStmVwnn07ZXxE2WrtAYw6+6Ys/Qu1NvVK0rJRDV03iXlpcfWr
CQZErxR4snpB8bZ0hhipxWEA2DVy1KqJbR1/JBFP1P8lQjEkjM7M4XzrC0DTkU/g7rGab+9vSMoe
r3bSpmfEyPRw6dRvfH+FTZUAy/CFQDo9Sv7OQUNqFGZ4cYVMbbAByqYBF9thPu2N/Je6KJ5H6g9O
Der3WBh3YTLdG4fmeMrQwm2/UM+4prTWhFutC5KZnksCD8UyLIiGZ2/K8evYO8+frLrU+JHtdCi3
iQQ4WtdglgjN3BDMUhQedE1500UoG9lAU3+3gCT/zK6HDlZoms1Nr6YzwXlFKnI4y8sVDpd9DX1B
E+dUtfsjz+hKzmkJ7zIi4q9I9Vs+jyly0Jz6nJ/n7wLjL4KRi3VTgWtk8uYqmSsyTrmUs5iAu/KN
IUnhxHzNSqg9mbgBxTk7OiF4KN/7G+97EeEfCn9/1/zScKKPNbJNsZog8QWp3Ek7zPed+ILLasoS
lKcE7QVy8PDAKchpbRzUMjSeb0d+fhM9JzcVKDvixZggP1nlk/noR3XHysHsfh8CyXbFToaLdFbS
c/Z3e23BUuGzcL6r1UBTfdOuSBTSr5QMCpm1FtW/+i5MyWodCmFuohmsC2ufqAf2Pr9yQD+dR5/N
Zbn5pSRGHgA+P9i/zd+I+M3EjJmBgmcC0fRReiv9gTyhQ/EIk0ZSmw3z90y7ACRQD+xgQTf6EIuH
m6kDRyQGu7+ci3XTeVk3zarOL+Td+0y9rgHre9HhbNcVND53pOMBrSEJJvi5bAlo0m431bID4k92
ly7S88s49ZeFcXVmU0OGBHm/gVzrSKeFh4I7w0xjh4a1eQWCZYyemzx2U9CK9w465vwgAhhVJAeJ
SfffMXY8u1ef64MIda9g4qcykLPVZ48wgE/Eh07qT+2Whi1KPSwetaBQzghzsLPcT+L/kAsDeha9
gExEDbbNEY0Jm17k4VS3nN/8/kZpVc1rw1tH49yfxfu4lIn4u0vS8hCixmY6CcpVo/y+rbLjoxuL
05159FYH0zGek/0CeDmA3T7UwljVJLtp0OvP5m/kK+++KXZ4sOppzg4AkN5GjuwbZu/K7TP73gpt
SaGDI1Eti0S3rpZcPrt3H71McZkMpeDvIhiUtRImNkMZjLw7bkgP7wqVGDspxoWgo8/EPs60r4C2
HhVDKRLvjlkrAFkDB7D2pwGdmcF8QmM8kkDnKxLT+bScV45t/C7QoiiI5YcKp+3O/dUIS6Im2uGF
zmfIJG34kLN/H2f7fLNE8EBEowafA0mXL3/apgIqV4zGx01v4/V6GJ+0Nc5hLhOesBMqc+SfH5jG
BcGCfEOXoYTej1a0WfyNZu9lGOXu+tVVPnxmGE64lPxVL5zgA+rpAjicxOemmxwe6lp1191k77hY
++xfI1fit56dxe29wJWpzsHaQ9sKzwMd69q0TZfwjH0mg4TmWU5RhdxuhUKj42IPyO04kZ9h+IkE
o+aAZ5CMWvtFTczPRu6j/XF/RIlEyuIyfluX+DRM00McJ+BszL4opTkDHVooUntt1oCGiTeFAeoA
0pgHyPuW6qlYoEIPt02U032HMZ9Lp6yRK0B+7diVTIn/b28FCfRtlzuIH+py+SQVepgzQb1bvpQO
bnZ2EQU4WZqaBiVNi1SpIvOBkj1WY5Awa56oqMPdD3i4oJcKrkzYRwVK8nRfRlBSTThtP7CEonLF
s/eaYrOaFPtQK48yXY3WbsE5tpVHivzqIPdaQbrNYqBPPZMgbbfmNUdlz1KkDusDSSc9ZcwNecCT
KwURH3N+odWjTGuJdqwxPwoyJ6CVYZc/A/Ff/TmVv9EO7exrm92eTECTqAcEiiJEkWTO8rZOxiHj
W71zsmImsCnoMu271h/aFRfNd4ngBkbj770rHoc+NsvrPPKi6a4K0vxDN/AiZne2kmvWGJgn4wiZ
kn3vNfHKUHQN4h8inX+MmGT3J/NnCukNtctTeXuf+3aaF8tIc8zJxpEbCCBPIw9jzfExEXq/J4HD
Jn1EbvDB4dCuzLsY6Yq4secGQCQeK8LkgEbDcX9/kajEVVMJ/0UoOsm+QBNCwcOcknAiGomiNi0y
I68JvjKEMRxI6ydS1jnQJWUG2zxyX2hVzZ2sKxShzT8YWH1laruZtoOzYp1DuIEX13byXBMLMldx
pZFGVkcHZ8V9j/RN6I3v57aA10Imy1ylX/BAS6PKD2tZ7CINzjMkI88rTO4gOsnWcAIEsn0cVbWO
lnfUlEKApTuPAt6dyMQEqzksGzKKPn2zfI4cpGub2b//RZWCyypes9wJ/lCMwpzrH3I682q4Qg4E
hdzGBgklXMF+/fz1tBrfD1Lq5OBXjNR8BxLY5k3tCykzn9muLyunjrd+KcWhf36euji0FYjZsivX
BaX49UhaQzl9itUXDXl1xmNepPtKcBZKbw9QVNaNpmcuyPMhiB/hFM0frjqywYIa7OcCSKlf0407
CWme38TBJXVe2Jg13SVwL3wf2lrWRS9E4c4klzZ+raenWWSmDseDrQ2o+Ko8Ro87GFNRyB9xPxa6
Bs3IR0jQaCQu6bwlfiPByGX1JdNUebBy55W1n3b08p3ZFBeko3GgiCVa3Dj/BLiADrOppmkTHh1g
5rgU34T1+L/QXpRDM6N6Rfw4NBUO2LwBeHNi7H4InE9sAOKF0EhGFn+6UoXddHMAWoikDHxq6dsn
4YQs5uOE4BnvJfA3V92hFRr43UJdiFkVihiBJYQT7J5bNxBbwiAMFwFFZPJKoacubEcy2hTAottr
6zWIJGTyIPJqAUdsKCOc41/7RSZttaYwNz8sdy0tgnU2M0lfvriJU3HjFfvP9XnFIrlfKGUwaIAv
5cdAkn32iUv678AuoQZB9L//UqDHpyrgRVkdFwVRmHYBqmDIzcg6JJx15ksZyl/bTcwj1RYzXEij
r+ssrnLQoog7UKs0xyhNhSlLSW7qpXa3w12GJ0YFj7ICemmf6n98xdDWf0pJtOt6oY06v6x43rro
90MxeEfFfIKW/DJF9BgCwy/B7vpDgPsnpgT04MU4GG0X8ULoAA4WsFCOXscsQd9Un0amOqCU/TjR
8y08tAsDW47Prv6u3fo5YFADBMP1YxcP8pNLbEzttqhu4/UOUrb0IQQ4Rwl2t4Gj1qD0Ufpjde71
OWzgG2ZLvruI/M2eMvIPAxmnjlV0chiEIi0cBbQVnTH6ijF+n+IcHMjdsvp+VkusX/Y1rEHhyyge
0KgStjnf4H7ZfPLcURGrUD9hVU95KfLAVfv3RlSUvOBNRWTgmVN7N9wO7t9d6qRI/E4GDaG08A1F
dw1hyi6H7SBU08HKyJK8ETbSHr8hLTCAQqIUY627a5ciTQFPPW9A6IZJOX9b4splqv+CpgnL3z1I
a3WvPa80ZecANAhUl64Gu+0TIvdJrCfW6nrDbRyx52QQqba4AHLR6TmM2rNfVaC14+cFH3fXin6e
4DUnkgBfUvXqgWFL0RMq8xVlwO+K9FPEheejcwsokpY0oNrCxe8RLiYAEN8EOzSRN7uHfPDARtuq
GIw+69aBHflQh/c1xmSaFHQ275cUJw25/Kd8cIruaD5VpWj3XtZzI8VpYZrJQNZXvoWfWA2Ho7Of
Kwmlwn+vCFaYgONqumqdNNKHfC2Whn02LFeVAPp5svl+7fmhK5zuTmlpyN72zwW+IACSv1HjBi2x
PvlT9kqAQ3obkxwqDgDf8da2dPfgggSvT0b8YAEKMdm+/tJ9TmDCMcpieILikTk7VY5V5y1Amdzr
gZxF3BKfuLoycbPv6cPoMTWrtWYuowSPjIrh72WJQScWCzNnUnIOBwxejoujvJsZO29iHdOkVrR0
IhDIHyVI6BeSIJkyEbC/9A4ZZKTeNZwnWNq/ccs+0GDI6Abg4ZX5TTAJPDsTgRPtCkR9zzXqK7Fw
bA27RRiHtBknJDa2ieij4e7oNOqlewDYCzQUanEYLKs9PWTExD7TOmp0y5posd91OjQuGt/+odx2
zJ0BZLvrLvtt1q6+VN6JgAIm2X9rgq2PXLEujoigztSvwGaMp+EwbbZkTsS+f9lgUJyN7mmd9FvV
pv2Mz8D666bp0FyBichtVAlVeBfeU1CTXEW7Cv4wsOz0FoRqJLQmxAIg5lEoyf3SWzgfsOrEl5a6
kfvD7aZM3aCRQO4Ih6fohwvPi2A/2HBfFMn8zBhYUUS2tCcBnCmMPLQ1Id3yfQMUFqkABxyYrm3z
Eo+QXKJE6iYQxbBq4k88fRQAFrp8FVbajYoFydadJALdb/CUlHRHKRlUZae25UozP8/rXd6EP8Mi
WonzFSG+ic5RKNZ05wstG/aQ0qRUKTaThwU7AK7wd+4X0+sbuUY7BqavEYw2k+GE+r1MQx1m3/8Q
8ewbFXjdDOAY/k8i1x1MU9geutHyaWK1H66lDJ7T8Fm4rOCZKWJCNUb6QYeC6gD65WTqYzw0eL02
VFLcuuM17f0tMvfBzrM0BchDJ7UM6gLAugONdSfVf3F1dfLKUBJBTU/HQfbFIsvQgv4v/KgvqocV
kWT+3KrjZ2CVKrRiR02i6j7KZy9wWZpIRPOhfeMfWG/Yp/qVs9wXmRvqTRK4/z1/6knxAWSfI+sO
wDt0AbnIOA2Z2Nf8xCbA/TviW5H05IhVwrKGX827iWlG+gU9OixI8+dAzOsTa+7nWFzPFXWt7+4Q
K6lPJLGjpPavszZ2xhZnm6EBiI/xfSqBTQ1auwZEvuzHKO9o2YzyYfGFOlRdZ5mp8hhYx+ycRXIV
cYnA1/qz0iGa2bmMrLNdAfCRzpYXVg96QjdApeglqiYLajRYDPZbI2GqFBNUq7qT0j5YTAXEbfBm
bGPUUSKeFbPdc3AzkQU+NFKGCRvXMllIVqQPizPTVEFb2T/fcY1YYbimH7HrjdlfSnYsEULbBNZw
RUflbbORjWXSACgboPktNE3wb9HPCGU26qkMMdQHe99003bRxGECMVjoh5l8fhTZJNWinnixx/AG
MXQv2qQV8QvowfdBfVDbW6nB8RD6BIGomHVoU/I7DbDR/L5T45lFObhmeXM8IWHAOP5cdNI/ksTL
OqWHPyOjcg1tiSTlL1/tKco0hCTTZOGoynCu6gmMLefYY1q+2FvoeDct8Wy4Uqm7uGN043mhwAxe
EPTFEa9reEG4SZs3SStUYPgylKJHwa9lJS1O/jozDOrI7sFBboGs/5hVdObnsaDjRS9gQJZv5jVl
1C/wsVFrFNVBd6JA/8izgDZzG6nMcOjc+bgy02llNzQkT19HgYRZ7aDhnmd3yQJu+V36Mh5hGQrg
aKhpaT9qznlFOIilAwEbcD/to0UQ7p8s7s6gFrLKAYBimswos+E6Dc5TAkLKmLJHOfdOfjEYa7Kb
wwfv6PgZ/qVqKeg1F7+aZ92nYcPxzkzAaxRWZUV9EIlr/jW9Uzc3/ly+IRhWg1tndugfeiKjdv8y
UIW6wA0Ah8EeeIbLfvt+mQ3YcgI01jceSwJD0FGTr48puHdmEvK/gtIj718PRR/+c3mBX9UXFhRd
7oJ0VCvveLKdH3N20TD1DF11c1trHPN2PldQQb2hcbS9yCB3ywX4Ci5DvXGoowJkESaxqv7sAjPj
sgetEVOQA5feDJzdmN9Cvk2PSTNZy71orfD4LwLnQn5Nf3q0cthnbRvER2iy1x4AvNFQ1kJZS1rL
uaVzm8ifFWpH1OsIzZRQcWldR0LEnrdxT6F/Wp50a0/5d3xRKXJivbjIXPKGwjzxAnLDhxFGTDNh
JOzz1r/+bk801/0tK56NkiAPrnDBadCN6wJDHW03IMTL9sJLZGmtbsOxd0XtENmw64juVK9LDV7u
HK5U56W1XOf0JQWd7wopESn5cHmuMrXfLAoC5mvV/rEEIy9tMMDihpLB0dr+mAQWJeuQTBha3NGy
wkE77AqHRAYmAKTTKMDHim0bBV2OmhZqb2U61TOxrx5I7wf3VUtenAAJ7uWiATE9tO90jWHjpLa5
WODay3NmoIvjgGcbPN7qPt0i62C88WpUUWctinlQOkhER7TfAJhKzwvWcffZsQq+vckcCHbpJ/wO
HWsx0/4kqyKksKoBRMqWyMPcbFqg8Gtjv0sPYeBU5UAujxNUv/dlB4q1qkI5LK8+l3mzhT/gH8Mi
zSsK1mebTQ/AMtM/LZKamT9ZRNgxB4ZZ95L1rU863Sf8KsR3fTcuZpQwhwM+FdtFYAyth64+Tf/G
WSvc+AuIKanIO6TI8K2z6O5DclbKeNzOAWip2tudcwS5LkFaLGkcVcHb+D5I6oGfMT6xYxrgi3jj
bVebsALInb4H4JcctLBTydzMwFwyFpblHejywEDlJT2FawBoW5RvMOtHMUaepYz0AdciLjn9ZwVi
75o5Fs9JVBOYxhwk3480D5fzLBafYEn2HUPuT8+f27DoQAdexbWRZSfXs5cYGql9YJhv6k9uo+aq
JfaWzY1GBP8R5IUdAEkX0GBtk6POuLoLS1hgWTkIyArTV5aw48v2s8sSSpePLJnnn812ZjDvGTwi
39082Sq63FczeX+AGaz8kN8OdRUFqRzyqe9RgD/wk3DXvFCS35XU697J6xCN5VsfRf6FwEczSGn4
PorHodWJkPsDlq1pwvur3lQrMSWRVdWsDkrJEYbj7Mw5YyMBnRsD46cc8rTNXfszcQyQPtgtW0ly
CW64ozMU0+GGCDYyHjGd3a1NBg8O3YgOn3Uv3PezL6iT20up3e+jvWcUGa4ZjT18u+kF5GDNt1Ah
R4aVQK8PqCITZHayv902QhASdIWrILNcpY2Pln8M3DZZyIqiTeMCXTyLt5m9aLaxzv9OV8uuP9wF
wIZUxULuWzJx0lT4IJYie5IQWah7FkaJibBXk3UjYcS39GAbkRiJALt+ib2pPzqPMTdUCNmbyfJI
yuVsQZ13YcwVyKhcks8tVIvptH1GCiZsTDeUZ69LQS2+1uFzhQkOMNLwUuKX9Z7xvwDBibjoMsWF
26KG7t4qWwcWR1+hJL8ohxWfOS2VVgiL59+SX58lpfEmVoYNwdG8+LtKF0RpmaG68WAEloWEHFAx
79QDlLLPKSg8xFXPP5U4WbenxkWf1rjfxSsDGpi2KOlIJFuIsV+UYymKPmq1u7pOuot3QfIhILBk
Se+wxl4eI/fEMVvzohhaCIXdRXHux8fhXol+5/GGD70Uwukizd5VlU0SLdkwHkMje3vs+GOPxDpB
pVYBJcV5dvkN3Y4upoUSM+AKiScN97O5529tEdmLe8seT/gTlNVTaw+azmJHtS5E6xnF16shKadV
+/4B0wOafERGKhi3/mwS9B7Tq0Kd+/e9te34/fycNOZDkYHydhXdSkWD4a/9gj+lURdoXoGIAwnq
rSf8uxMO4OnRG2vYArG61NlHC9u4uAsF0DTOI44Zun50m5Fsf4EQDjEqlcTsX1lkwgQXG0hplNJS
hd0YKQnByeerxrqG0ccPvHME1vvJi34mGTXMpdmetGCSMVBlcTjMGrDNUlIMqYiixNwA2cnUntaj
K6WoBUF4YGbvFaCioC12OEL0AtLea7B0xsLMgLZCIuVGRSVzkWVT/i7GYaR2rUAicYfGzAJY5Zaw
1LvZB5Q5jgs3d0A6p01olfqBVeja3YLwkZQ7FjEPGsYsCbjPvUzVJPcnkubBSfrkz6eKZbrwAEkv
8ahkMhLGKuh3vj4Ky6odIeYEMA52iXDUUFZI2oZXgy+rsFShgT1IS7JzzKGN4jNDi3J3zCaGpMyE
oepySYpc/SLfm4NfcXh7FrFP2UviSf13gTHjLQGArBnSVtJkbNUmFprKgYFI3J+UxNbxn7D+9OXS
4m+aMIoMwtt4KU4iyL3O6PegFacciXyUZqXSwO+Ue9tX6WC2MkOe3PHktNievqg7n21lEwG8QFSq
1CZE4RBuXNM/eknCHiPLeg0WPMtqCDkHdLdmILCuPZUlV1VUoSlh5MHtH+Coo4N7ZeMrbG71bvmU
CPwZ4zLls8bfIOqBz1DVOFRZSTFylANrwYB5qzDGzIiPwXdr2XchR5ye9HK0Igf3U8hRULsNNRE3
KS1v41bZvnWrSlE9D5xRfBay390DWvUNIzaYV/FXLYmDEWxsokcypSsGcoGn7aTpNbYj57vtSlRy
/Eq77wmDCqF0nAV8+7MOATX1yXpLLE3RKj2hggGXn8+2h7rRQQudXtG/q6uoYLLFPAjCIGlU1AsQ
1/vS++DEyK1TvSvl74ylzBczkkTBS5Y3M9jMb7PSNBY7d/m/bBAo/4OnnoGd6de2TkCURtRUrYP1
VE+AIWT/EtkWV9cGmNjwsFmlbepggjwl6Ynmj5/EL/e7TWdvHH+QXC8mxzefg4g93t72un/lZ9+Y
Mf/tOStEdKCULcbj+ewS/g8pt2sAF5esk/GPyTuOSaUuFrfCBJqVGYu7/ICcrpMYSX/YukJWi6S6
HcdAuKakUNN9Lsra/skYfEwFywVX01nZeZSvWk1BaE6+l+VY8dbJbmV+/YcgukUCJNstFu8XZeXQ
V2K6/Kq6PpultfYObsJd3clQzibaK1aYeitV+KqnsD7qL7Fu+OQu5EaJIIbiEDRkyBkglWZWz+ge
KSxVjeo6ja06TFBj+F/jTIVxp6a5LoGQZhRLAbuKUrF3Mt87lIerA9zS0cP00A9u3QxfBmsPU/YM
fyawO9hp54PjIWnCsgLmXL+khUd/1lpuxt7FkB06/dpIt2CzVpKCWy13K1h9CW3j4gd+tMi6ouey
d3HNBATnBunHMd4MIMmdPyzE+YE/N68hQA4x+8NN7R3SFS3RlVeO6AlBArF2M6MBhHMT80OItpHK
YmOyVkIq6bayBi5vw/fHB8JYN37KuOzNDbpMR6nt4Q3iTpk3h5cyEAKsIjxLAcPUgQt/XcT39y5q
TcDp3xUNWtGCUzNE0rCR3BBdIbF1b6DJOvQRFdjiTNbH+69LvXrFi8YHavIYKStCBAl7KsYc+fiA
FXYwsiNETUiZo4xCtR/yJeKV4/n2wIOM4PnZ2GN3Y8jy/C1kaVWysXfME9391AiAWe3bzIUeCKjl
jJ+JseP2RQKYeJmJm1IukGhPA9E00BWNU9uvTunDWB8ipcA5b+BDU6nt6andG2wLwugcRgUpD7kF
CUgxPlFmSkV43nDlwzpIhitJJQBgscCE5oOxd4INdpFmVht+izOkRdZKANa3ruyKXaWr4wfR37KI
yQBlp1qR0OiP7cQmYCHi9I1ZZ4bsp1O1yDuxLlnB8R/Gh5oOjNvwDpVxmQW0vKJ6eHrK5zQFAjSb
qbXLTATts83NXPOy5XIaaD9+dcpVwilSK8A/uKxqUvIIM8GO2llaiv8ReFvDNB4BNW/XJgGr7cD8
zlA1LK2LDOt4uXt+Ajeh5YHuBS6YvqKGcMejIQHjx0aAvnLqTlJtzwfc9u0bwREoH4eZBP4XA1qB
GCV189uXq6rda+wsA6L2hr8+WwBy3kprT5DJ1VjJhBKdVCXEOYpWyD+FAA7vTPeOg8fKeqMh+0uf
nfwd35jayiY5RXYR+p8PwBpV/3n2PdHdbILQAJK6/H+kZL1bUe25ABLMFAIzcjJcgvag8llPP25X
nJFfKA0xjpToHjl8V/2268KqzBLghuz+hR6qtUwlJZPk/tICxt87+cTHhH18wHhdF6StaUfCzNgO
kiHrxkoe+rLwjxnVviNN2dbW9EJVxf8+jmDbvydMGjzjo0d6AtHnY9qLDPlXFuExmauT6UWw7Y0k
QzChzEwFlwuZDuEPAibgkK13eJbYQC/Zsg6+0bUdXp8L5ACaTK4tTkjKY3HRHSgiOQmQfEDJmEzR
EQ5kia6wkY/ldfi0GpcFWM2F7Bn9HT247PFDksMKMZLVbjUO1FfM8BJvxxvi/aIqeupX6NnY/5J2
S9P1oMfOGaULiDwLoIqUgJTPkp40v/XJtnbpeRfKeh4ScSD32x3piqn5/wy9LgLiOmR9ejtoanTD
TH5S662X0ekABE4hePY7siamXMKR0mMhkUG9zMbaMkjP1JLkqg+tVbl0h2O8PHK1SuJtiQ4u3kgt
iEjx8Z3jCQMfqFuF5vDQqxNF8sLQkZ1giPQ+6lCgmZogmznd9dAHzIQ9QuH171SNeddnQ38QSfLk
VDquzKAk9l82b3tQ7K0Zx+8fVtpSxkJ0gAkmV/ewK7wZiZR2N52Gpq9jDdyP7qxL60JuGmmq3WLN
HNw1FXmUU/k1uhAXxFYpS3551ioQwSxh7Mv3ReK//gTahiIL+FHnTFnlWLiA7Ud8l1wua4FtumNq
MQ2ZMn/dnQzVbQTX4xX6gSJSjOLm//W1ZJ4d8kHhll9cCebXamTJwR53NdNYVEycfTWAIUUfS1Qw
jbv3zBuZeiqeMCG47IAkA87lRKU/B3wtPBVzuqlbgNzmhyaewEwAp/Lx8sFxiqtOn7clc92ijIvJ
1rD/wiuB189VAhda9VWARlJwIC8RXrK5aXIMumzg/3dXPozwHtHaGA69OOrM4WZVBGBMAGJk1ygq
tjoUTTIffy2RvHRPcO+bhFChkyssbkiUWYJTwCx+UYWJ5SQ+qfcmVVpKB0T5YtqPS7k+tXPUi6IH
+K8h7y3IReRyBABt/x0epZidt/F84nuOwUD0tRHrC296aF6lukK0rCKCwHNgg37dKQWnpErbBRXk
kyflV5pNnWHilL5ViCW2jmEW7hjtX3COMN+lJ/4040x18SKawtshFufZTCCndJQ8Oui9poX5OqQ0
LMYlLlY6xqBtuEc6Jf/CiCoXdqPsBhc+wTZt5/Y40l+1lxrHpRvjKAKtwDTenF+8FCyqrTJQjzD5
hWRJ5hzI7tkpruvYrSlaTmlHWLKvEeJTHDzVAxdk2jiNGtGoP1IUmmroOZ5x2EcobSX9bujkpxOP
xr9cKFLtnHU7xLBjnzx6aD4q/7Z6fidPmJjjnVCKHjQWmrOfPFAlEk5Al3jlzmhnl5LDDs/MwCjw
8QL7E7Dcn9SLSnrF9vQEVSuxqGz2cc4769RxfcewUYiQyifE5TFBu+e6esl5nXddL2Ak2/nHM+wn
DieOWV5AlmbdCzm655t5XE64iSk7MhvMHLRnfUB8NrgqunaKYlsj6vg412GmwYzMuuSU12vdRbBP
xBvBVQ1oEl5E1bEW8rnKSYxOpUZqwemcGoHR+Z2UzZxGQulfdw2nxR+7GpQFQuFHImXt45pNoQA8
2N06IQM5lL+Ml52H1JMPEakqRZFI0k7lzoIki7fyyw6kU8bIjdFFYy+a04f0WSenf2gE4l6JVcig
twAFm3qTYkdIhgrvjRXBknKdQ6+NmF4FDHaYu92hv0d28AFTXmaVNZcpfa1uzBMQ9UMlkUEW4D+5
eco5ST2/p9XIqOnKKJi7IC5vmY09L2BAkTE+JMxGIeoGrKCYHj9oKptwJ5oaq0f89/R8GER7nns5
yio4r0NhqF0jd8zf+oJv8HtV7jlCDfouO7xkG/W/Qjbrc3rKmIFRvX54+zFgoaPnHz2/fCa2tecJ
8AFIebEZgS3RSq1YCS/axpcFZk8B4pJ/SFV5N6ZWre80UnQEZzdHU3YNqkQSU7NsfVvrTnuOdaZT
VKVclKEDiLoN/1nuvUfXfKsg6oY3dI3Iu+SgO5XQ1mJIMkhd+BDIQEtT7/ljwR+o13Ui2RFpL3wI
MgdJuUV8DjmfDCPOGmETF737l+fsKg4l+7z83pbJFHmmQ/IYPXpFd4EMyCNvf2tO+KBzOehTgqY9
JtUWQ20nU7bqaDZE+ky2z6QbT+Nzl8nznQyjCGulcXWs6XO4N+xRMWMNvO8TIOfryLMZDlvLjtRs
VIN19j6MblgPVmPgdzJu1DwuADIxlXPFjUneuBcgbuRD7L9qZ8dCZbkvt5IyciI4JEUQI3FBHoAr
7iMlqt9z5Eiw3fR1Xu6m/9ZHcFp4YLhKejr/6CXj4wOO4smHRbrURcs5W1Qt8AT2NvaCqhdDIH24
IyVSYTN0vB0fpVio9Bao9Zfq4MQuyoiqQLDH2Ppb89KvGnyGw7OsQNhICngxV/J951qmkS30GrTm
uXle1jLYMWN8VQL1qGX8SwVQWVVH+1RvJvHuoJ82VvjE4vHyAyUlQ3zMmy/oX+TtkJtrcJjXspxo
0tODi71ijbdIFKfkwBXcdHBHNx2MMfkuS/imTFSobULMPa+kushMH6T0iuaZQzo7CozjcYt4uWAf
jo6Tqcz9Yu4NrRBxjG7HFAcKP7T3J52QjhoVbWUfHX43wbv1dQ0iloFaADoVyBydozN2w0u91z+N
LPibSRBqNACBg2voYfUsT4f0CgKDsj4mKIeYpwnvFZ8mmzqVhcmHPFdxgUJpzSgNJbNJrHCW75AQ
qj4RhIXuEQyxt2aZHGaGB0mkqVc6TvR8P1i5/hVVdTjW9aNLxlbXaq9Y54WJ9nlk4aA8VEXNbYny
9mDyVAW2aXnNOaAKRJw3PMIzQNKAUyFJKtqqySXfuhle+HwwIQxPaMg+W6LnWMlLWLIHvSlNM1Vl
6owi5MInO1M8YiUAFxry7XoF5p/+z8a5Q/oWzoqu9ouastTpQ+EYmLPrp6qtlJRtWl7yWG3j8Ozh
a7hEiqCCrIjVhYusnDNN5LZgtuTmMj3SzjJfA8L+kkVBTR35wntTzKNNUW4nF3ILwsHmVpaQmpbx
Fn6iapEW16pKMyU8eP3I092OQK/+EZKGYpAFgiKNupWZQC2t4J0iqLN2ht+VFclhV79O2OwxdTtH
3lNtVmvJdyfbTtmymf2GwCEDk2RbZREIT5zINoGBsWM4WUEAVTkPlHStjzMvwKia5l7fcO91r+UN
wfBxqymSTR+7tqyvyfsm7Y9gHzP4sIvtr0MleRaMCthIqRwmuFM3h8tUn2GL7YOlHYPriOzC9gn9
OIN6JRxMhISUYRLGnAvPLGE6sDHghozY0JDEWN1w8I1Jo8ehQYWRyX4fSGEZRM65NPYLyqD2iGJx
8nAeDv/VzuSIENVIrRJzuzq9gpwiSus5EecYjmpYgsazGqFHaLfZ9ncZXdETgrU5S/rRg1O6dLJr
ktfNNBbuL+VjgxrU7ZDFW8t5UASymMTLQOBdvp+89ojWaLsxRptC9+PbKRZ21yUZw5wTCiX1qKzd
fPI5OO73Gf94F0dmGKXqNMj8oKM16KM87tjlMcyg4jryJOoWOAYUnyLjVqS5n22r/E9M6OjWCtaJ
cWbedP8mCuHWVEbk5DcPgP+It9AybQYRZXtg+Vo13d36haq1O/XaHCuuPI21vn2L59cSBUWoT3wn
eqvA95OCCGOszieoCGEreTIwunIsh5X4s66MrOGs2GXja5vkbJfzwgaWp/JkczXvnprtY2+t1l70
R5FgGwnglWQXXpWNzpi06knTOnSSDRIDAYT9hxwr3qeOHpC+2UQ+t06EnzozSF27v+1Y6Op2gsMT
iNpJoeeCWobVxROd6IHkGYgl7VC+BLFfzZ6P1sRdp3soQM5k2rgnnPLtl9rMs0C/h/vHsW/puCJn
bPoUw1F737hAvMF1+lddIkj/HUJ44Bf632Oesd0fI5FCfGxOP1Si3R4G0n717dIf2xiE8fwM9HkO
3eFFF6PZseA8m4d66PdIYZ8mL9kN0ouNepsH9V8ELwX+jFKUCX+2RP1DGa2GEFRlpoV8VgINc2gs
Ls5a1DqxGuXHSQUaqxE4rlXR8t6oQLwEWFqGuvPJ3EXb++HawKho1ObihBJaYrvNQGUkOqsiDZ0e
4/utyir9KuzHYnlYA67t/MetFr1hnzAZ5f0ufZroNlTHd3bEF50D/tLnkER4Kj5v0y9SyxZfdqAN
jLZs6mHX8AeM21/66dzExvSkBDnfMOIU9Ge7KmWEsW0wlOKJL9rr6FjwSjV/koHQHvKapjjgGDWb
CoVvnjFlzqyjs7CbXoOdn1s3+nWtHx2bbqqUdQ3sZjOPnfrPBwYTpmWWFrt3zti89AyI/e6EsgHk
lArwKFDq4Pp5pIevqBAyHBZXBt3B3Ijvf6vmofRekw3DYrNp+iEEUoqO/3E73DfdrwZ7iAe6+9mQ
3GdArVPub1sOPYq31McPmqJg81w+YsQ6mCovm5PFoFQ7qVovn8ujCQw7XSVnzEngutzuiswyXPnH
e3/dfhzXImJidtNgrjgC4o9Ej20tk2HH31t2f7ndGLQKC1rw1WoAgDT1fDEFTLs+fP4DN95MYblM
Qc25kui+MDrBJkElnnyKh5s68Wfmvt5bEbYWvMjhKxoAr2ES/R8sggX25FNREezHFaR1n+k0gzjX
O94zHTb44zrDQ09eROm4RpbblqKQ2HN8naUKCzVvz+iPJn4A3bQsDtup4RSv2QepytRIvPpEMEdC
iOfgSur5eVVXHSRlESvORpa1htcBbq2r/Ee7+iHhYVPMgzdD4xHddqpLIlvnfmK92XEAt4X0WLwo
SH7kjAgKDej4S9bBJE/TEz9NXc7xiVt8IW1aOxescqa79L54fpAkNBKnni9BD9i6IYGo+LG40Ela
Ou/EsYik6QqZA+NjNd62PUoro15fwsyNCQRvTKsa7rgip+aVbSxq6veOgiRsV94Qi1hV8ruG7s+3
QbZ04BmlyUAq0vwX8qjUV8A4Kd+uKEFRFqL6E38SeZbT49gS10SowtKws+6rvY3UARGA0B69bpS5
nFMHanj1O+HBYjzbDzKzWqK/pRX2yRQU7WSljPnGLrp7nPMhlXajYf7r1FYkOwA4YOoMIGEww/mi
RxSB1Kz3SnweaPJih3Ems5qOeQqboJEoOz4YKg8UKKcMq5n9Oqm8fFDPTgn9pZNTpQx5fVkSPTbr
zykXgYCjAMVJwfoYwXfGjx6ctvZPcQwmeDazHEkEBw9SdhPNQ04KR4pX+UmbuFMLQ1aum/1zY4n5
2/RpG4YRjElQxowYaD+27cW3cCbmiBEwA964S1Z1xF8cnUhzKafq14nqDL3JFhygT3wGIxd/Ncag
/f3rB4R5h5mwnxqfuWfGoL7B7NTyn0t84e9DpKzIk/zQ0ks8nNBOgGMRUN/sA2JqG405EN98ZnP6
wu2D7Dd8B6aljPaCjbYp+t4gT5XMcchFSE8BBuVF2/SdQDsur/UqGeHLGvf0lgByDem9xm4kkQZf
nT2aLpEyABTgcSQXDHDUZe9AtYHmI1CCIlo+Y9lj8MR13tydzUhjc+DaZhtOjphLgry165aCVmcn
vPNUTGfCqxP3nc+AORwi6LPuvWGHokz31dP/Dwl1/Pc/PhFPWepEoGXFVKHmXot00EECa7de5cXB
aavN3g97w4snRpSifnY8UeK36BNkQcvzAXpwBHM37uc8u2WONS+fr69JBDE6Uzk2ApEkNLdY2f+V
TOSoEZ9cYGGz+XYYZDQ4+FCRNtH06wfTBnU7zXUK/1Z+2bt/NNmhsPvTp+nPRXTD86UTmgYZj0vb
ugNz2lQCJqP6zCSWpwH5hJkqnPwBqXzrHpwIg+JvMXgkMzSEVwSjJ+LoCkBkAq7H3w8MOHI9yd4N
mJQ3uAH7sFbq0r9QBUG7+VGDGTn1R/5aAzsr5LoW2RXh5bmFe1LqjjezXHNapydGGdi1xMGZhWbx
Vm2YsuaRvpOdTN/nxNAXZb19su6buqV5KHeqFRcgRjTX1IeVrT/H/fQKRQfDT6kItGnkxsjnjWhm
UesxcEYCxUZ9ENyAN8VPck1VJ0FJSeDR+u4WBGIT5fLLgt7gqhoaM1fDGDCFTO5qKFzdmdYsUX06
Gq+tWUDZCt4sULFinunAzUlRHhBGTkC05Q4wl+T1pKbMY1sPwSEhO3JOTSZJGXqZnVpXibjWI/m1
oPY6yIy5DiqPxvn0nHWvkDAx2o7ioMPnrLBw7FVAmCtlshVx8ZubYNiHaQ+fJ5RrVm/0IDp4tC9j
oSMnUfZKzLThoH7pyEJUNyRSg2VGrmZknccbZXJaf/6z3dEITzHjPoKMTTHsLL4RAWvpwNkXtaAu
iIHPf9+GQTz8Vmyx/XiGFyXNUOta2YrNbyGtvCiVRm/udksRRYVJHil0boaVG+YNJlkStSwtY6b4
9+SoQu0eSi4asMNC1fgUAPpY8tAMNfl9VYeUqftxBeo3p9zCEvXW37CM/v2KaqJ6pZG1Ai3X3QQg
HvrhjtCPvDCYm/IqblaFBqOzkRaBWT8C/X6g9AbdCp+sDzyEvIqcOZj13baLWiKN/SABU0wahWh1
dMU3NzZe536zlywh7D9AM2HlwzU1k47f2mKH/qYgHuaDoiZ5pn3/JduUzg39Z98uQhAXbBbxrGO+
LothveH/oK9HrJhckDQdCPNa9lg0aLOrpYPtqTYq18/OoSglYclAwTKj5/5gdmCrlsxhjSKiI2nR
OAtgNo7e8AojHHU6OgPBH4Ewu72Ryt39vX9FyB7ETZaUnACoZHf68p4axC/9GMIfJDDArO3IVJbi
W8CnUjLhSt4Bezpcdms+p1E6HaH22Z3yMHSKVzcZAyP+vhAKMDdxW5OuIp449XMjeCCrL3E/wrLf
68cFI5ZJgkszHQCxKjp68VsNvMUEM4HuP/BAZzT6Z4+nG02yriLRb5OvYxgEtEeK4ASgtlEoineO
baNkWB/gEY4sWz+DXgug2nUJF+i8738md+fg0mlrrpxz006zOdxdfThZCrxqgWOOXNECd0aUPmI7
2lDVA/QnXBTsIJWLCzhpYx0oRREb/9h1qPQ9jwxWHT18BWfCgleckgVsFLe94fLemg03TIpMQbCg
bANex0G1Q+f+k9ecN9UsY3cx8XAUJBgU+JWJItoOWo/zRvSR5ZXDG/mV7JtGW8bcRTUsxkeigcpy
N+Yk8+3WMSEbRCjMr8QjnEIZ0VhbKLqP1XYoSkOgwPsf7DFPFlIEbQq15S3XZG+RzHW3L5ZFHXAk
Y5+fGTvYEQNCpHFGitoaXoUFFn7WkMcB9l612nGgh6O5cGPDRl22Z4PZs7Pv/Juycd4GfmzLigYk
s/Sk6xrbtqzdBr6cXjVd8fRQGT1PruUBw9YiM7w/C68+Sxzx+8MR0h7luXHjy+s2xAODxdrT2L+p
IZKtQ70XiiVXTv8G6EgFXCIAe3ppiHE4iEo1os90HYYN1jtFPNOMYq6rBGEHZ6suG+e/ejpFevDT
or6CxnnSCY3P2g+xf/yZbclE/MZ3te0VHrgN/pruIH1yJ1uGUp7YAi7Trdc0KiLnMUzFCrmimLUR
SCjJKgrKhrNuMWPr0ufXK8wBveqvi6LZ29LINP4yMdYENjmt74aLrFaVOYqCjaxGQDQ/486Zftp0
ZA1DtehmTbAemv959cyg2ZxwnlLSdP0vXHfkqYLjvf89jwTQ8v4oxjNqNPMMoRkavUteMFxl6cCz
DCzTyfScJ3My176h+aIOLIUnuAwNsWMq/eRNwozC+Tt8UfldHmS/W/lnwOkUO/pl4EeLIh2yaM0u
fOkps1omwWQvuDz2H8zmWFEL/Bqs/xRhYrq4G2mzJrl4IU22jiSI2ZOD/6dFD21WVk1XUK6jlhOv
ruuURBoZJcZ5StWdmG8y2U0x06PnDjaHcnq/q1hnaA9RkMHcu6W5qBbTsw1E1WZdUYLA+R+hBZ/M
tRPs13zjFmiFKIHf/x90e4IfGbgdJtdUrk79bXpYCNLGP/y0Kktw7tFdlAG3m8QqQ2fPoPXe+hrv
x6sB6aOUkoUzxM2bmLBVWFU+3ymwDM4VHiBHaTlplZ3svDSsqMaO9/LrHKmN8iXEN3imhQb8St4Z
t3PwUToZacTvPI7yOLhHDqDZcbCuS1M2iwACK68QK2kX5cWzxQiaNtJhwXHyq/aui41KaBhzRsMq
/Tp2NpV/nW/neP2kDxI+F6dZd16e6QTwkob8CnjQYI3mMp3qu8QcUq6xPmjsQx5LonronBhdQNsG
V3Id3YmgoBJoGZ8uSF9wM6JI7al6uI2IiULXyuTY4RI+kaFltSlXD9uTTluDSypv5vdSgHAOAHOF
sAwgm9FDsmlB2NuX26HAyjJYRvKtRr0YzK8yw7cQ6WpGVWBRe9CTfMKHQN7tAGdjKDu+f2u5b4oW
Q/KgH3fHD0dGzdPwEylbUnLQXZ9Sqr9/el3NzHCzJ/WiKFiu6iNqiPbj7n/5M3KA3eivFDVAKrUo
29xurcOsSCFedEOXuLZdZ/fSW7ZZ2EYLAam2J2PpQi+nzI8e21ng4P3pboG7XwHKyvFdJQTwcoJq
vUrkxv8SLp5jX/ZjDWiOZki/xyaaU61E7GREOtKJ1J1M3cW14Ls+FB8Tt60QxGXw0XqA74Jq8PUX
rz6/ojphHa0DKwFw7gguKreTaEZ1hjL/Yb84Ggs1efjSfNaJ3/J4TMx4UVVBD8aNca08L3BxRnjs
/UTMmiiyR6PeDfTLl475kMtHJ0O3/9N1qZ96PWZGeU/ccejViauxeoDQ04HA43tvfqkBOrGy9Tzr
JIbtAZ+2aw3B9D6nQNrZ255UKSrqPMkOnzPYWFy5beFT35RqO2wVlkS0kNV99j3rqEH+zNpuPJ3x
z7xHI8CiHhf8A843fLLSyXGoPzL4ZKqudGFz/61IqA4nf7JsyyHdnrwBxd/E1N5v+v6N0sI/Zdrh
5H2YAhjRBvCKWdZa76Q7akOmpo+ijfOEHAvCB7lyYKT0Uf6Bcyo7OA1JJL9SBfxdcnzCjpmCxIXv
D9fs2GBPla+QOfyXKM9AkEgjDQqiktsqmfkp39bIRmqJS8pZnAIVBFraG9K6etzZHN9AezZHrneZ
gIL/Tbij5i1kP87h5rT6KutI8bN+SBhIGXFmLh96W3p20sMLjpL0Q64MTMGZ7ZeFHgDp5InEnfOR
2/Yg3IABIV3aFL/ssfG5j8g7FB1nxBTBS6f+p+DFbpAMWLQOVBPqv+CrZMj9nThESfzvneMr/2Q5
YPbOSm+S8iYxm5T3ZRlGFQuyH3VspemwSQSwDdl7gcIEIR+UG6LMeokEctr8Aj/u2cByOxUiJkI3
9oiCG2nPuvahpnc3AnZE6/AlVYaV+RxkNGTvD1XtEel3clOCtEdj7S6CfpDPmdL724cIIghRUjWa
Q4axLeHy5yYgxbtgRWUtR56VFLIzj11OE4OiTEYcqHM0dW1bhDh+NT7y8d09RN1qaDQ7IImCSzjh
KPqiklVQQbIZhNB62FCsB7DUqo2iUXjfgcaqewJzKVcA33gcBLxv03d8VxTj9VfL5s0rBTejoHD4
idpgkM9amSZ5QZg9jW4Trq8BomNiWsrj8qJOHYAy/i10yhsSuyWHEySNzseZhPJl7uNA2JKlUpSG
qCMSR1Eym1O/hTc1aSzqNkZZM9+TalWtpsrBbfSlvi0jQi1cYAmhxN7yBBHqedSRsOszmpX6tgf0
DMvxk5N4ZqJoFYgnTgg9N0vmc1sGvI9frhrKVkq07zf5c38DRoD0YvLU+3Nc7VH/A4dB1JR3mif1
0GOyNZVafU5C308fe3dqyb41yG1JJ9Lf9vUwYGX4bKFAfXgkCLjX3XmMEQlzc+w45GDBbYwKvYMu
1usTo3+cngffqRrLF5iFdcHqCqFC33gC/eULm5IfFGHUw9o/nDhUatX3xVAp5D0/5q64RrqcamVS
CDZNhEc0CTBT8H0JIULkXSKT17FQKP+aSs2869pDmqgPF4Gqcp7NDfx5MWBiE47FcQr+glMXdqri
ZhETsvC1TMX3S1PP1vOXr4SvmeQ0eRA5hcWf74T93zNBv3gmCGJWD9z76ZM+X8DAwOkY+yDwPg5y
AkpJQKXYRSvCFxngYQ/2rrTlz/MSyd2T5O8r6AcvxhjyYG/wtaAjq1yL4z8zY2hDpxC399BHF9Iw
FbEC5WDvh5o7TG3qVhjFM7RLgDA52Kx18qfXWycZBJ3HQAi1IZOcU1vNniwVt2beBeG56hoq5G6A
D1OugBWZz3XpFCe5JF2drnzUavFX2+ygitZDy1EqhRTH+yvssLQdPHUcdy5WJ9El3Ivjc/inxbJ4
qQ7STz/HEzxUNYYoy18BlYpY/U1kCsSS29bOo1WSNm+2XtUX+85nSzDWP1/wsa+X4W+ojKmtu0hf
tDu74koIk6TSUTL+gebs1FT8VhdN/jpBGkmF09GlFjDhQbkJp9DRTXfbIM1e7loMWbTeeF7oJnX7
uy9uu52bDuPkNjt2KMf+pVtQwO0KMi2x/kt2XnTV3fV1Y8jTNpXZVePT+b5g+72oVKSeHyVD4vkY
LYg14hNErshOJE69WXw8yQgve5gRhE03KiPPQA7BGqWTMAfoWrcIx8WGiKPz4c2IKdf8IUcaC/6b
B4qa92sXSkyN7EZ1sY6qiU9r9Vaitr5fKDYunhwz+MBsnAdfBGy2Mirw+1jLnVBt5EI6ckxOXwjJ
FL0DnpuipOt0M78Xwtr1jxi6zwRTYsr3VWAwQEjZ5SCgLoZEH2YSmAGVr2zQ3jMZnrRR8dCMSxfP
KERjV49COlOMlxqFTtfRSVboNn0RMmgcufSyglFxrDuHEMgIs4PzAUhlWtTeVq+H7n/PaeooXIzn
TDxLin7HhCX/msUJMxKHGlCU7Z6dUuaPDl9/S4hbADq6S+eHrw0FsfQuPbs5anC01E16h05DbANF
ugiUkTzo8MDJ+C8lpZ3d3lFg1KoCrUR1SCWG3Bgr1R11qzpOMiZ52A2TIMF6ORvf4cVrEXqBh6g5
1Ndxj29cFz/bTKqO2hGJ9EJQnUlyKhAE2TkKeZ5PQBSQ2Qc7wD8DEkk1AYm6DUoyAQsn0yvdtYA4
0/8DdYLI5bFjc+eRox1gJPAuL2zJVXJkee7CllCv1bJyDn4u3hven/70Fv2T77EGSYj+LMfIPBju
UUSzomH6BHWGFVfuwz0R5PLJ6rChVEcV11JChkurJb9vu9qsQq+b0vzlevv3cFDEiuAX8kyZH+At
jCfYZpDoOT7W17WEmd17WC/Zsuiqlt+Wcva0jNLEw4euPrVxhmV97Te2kNjQwH7hB6xEWie+qFs1
T25NLbHp90PWrwO/x8ecdpOCAosDQrsyH8PIF3eUklRMVnILbAGxxWiMOLTdimdm45vI5TkUvr1h
sr4brmn25R25oHTY6NPK18FSy10LxHHIkXuqxyep6ROcBADUIaIK6Q5qytke2tWyl2o9EJ57NMuE
v8KW6Mt1HyL/y7ql4M4hQi3Tbc3OhP97YJtinfbKpC7fxLt3fTT5XCnYfs4Wsyp2V4pbP5tsHdWr
/SpIeQlSOhkS2MejuDtf+XIQPjkqslQ8+mmA4wwHck7P5YfudMiLUV9LPXvUVzABnBg5ApHsxe8P
YHVZL9rLKozSnCwG7slfhkCeaaTHJqYhPuRHr+cYq2qJ9mZNN42+dZ4RP5f7zaaDhLDsgL8N3zwN
WdH0Mb/ueYeGycA32i/Y7kHMRkeUbkBye3v8Jm5fLn0wpCmHJpFToD3AMMpcOazjjKlULuCwdNZq
1XSfAeyWaDO8IpKiaa76b406wOlLXpUJUCSfGdSScleEpOsR8e32YQ3EGeQfTWLJsJ9XRc1rj/bk
RSllMzhwXfuvLZpCh1pb0SZCHp9iMkhgfjWj/RqFYc8w87I6PF8Fxg4brQqgKvERLF4RVoGI0DlG
kKSE5D5edayVkaE+EX8HV4HI9lxcTjK10ufDCCo4RanCFGNw3OXUkBq0p4AhDo9GtEHC4WIriX4Y
7Ju4dLofOU5tXL5z+gkwC4EZaJPEdKdArIeqmdHW2Hy7hNh1witkdzwbD8HAhxaPaoT7CoqClhCG
qrGzLsAaaFF47QNXddXuCRyWeyfPbhDM79vi7CdNcImZ0STUcLNsdo8vb6KJk906M0mA4lohGR51
+A7A/DwVhQ56o6/vw+9yGjgAT8qxt0EyhmlkcZBhLeMHufOkH/Qt5zBU8E4dMxbJ9eqgBvvOYr6L
sU5BLXqc8LSakkNj2Kx7PFAfA5cFxVh2nJL/kP4vKAVpVR/dYEGQAk+9XEph0sBhxOwR0QKZLiWl
I30WdLLv+Q59/zacgTzvYEFoKhw0WGlPMUDnJrwojoVYI80jKQqFTQkiOhmSnyOY2OGXJw552n3+
OpYdirzcWh3yf3rC3f/GhlFNpKyaUKHNt1K1RVBsYdRHrM5Vgu/5QK51cS0VTR7azGlOSSDS0fr+
FPohdu6Z1yb2Dq98/apZNS+P4PnKq0IhAPjasDr0H01TBZcAXZaSJes747CJWP45WLwAqj8XbpY0
Z73odB43EayKLhYRCFT7H1jrWcmRb3kpJvQABj/sCF6S8i8ob/3bzXUZT8gakVCImbEDLfRNS6GG
6YfkIQwtvWEcKlfsImEtrGJHcVhcWg9JAqZTG2ILT0wrs4+uUh+N6v4whi5VZBuWs5k4P1C+dqKu
2oUxjPEyk2mpnjRhaSStuK8rCBmwtmMGXaoQ4fxNW3zDdnKdFJWafdonqPTa4irCRdNFFeWwanDe
GdzZWaCL+S6aVVWlQb4zyJGSLN5YgK7eZa+h7BtDjuSA+F2lemt/zICDSGNOTZI8HB+dTdIq3YXZ
+ekB5dUftiQ5L7HWyPdnXOgBa8roMMc+2JMgo0gc2h8KMGXlWHJ8ThY4zE2KVvSvWd8fzvLCXMmo
dwbmiwZgC4Q53YzmFEFNYiHYLd7QJ/0zeC/Ic28B7Ma81dckj3EKP5WmGRMmUS9L84VkOCyjwe3I
z14xb6VhJxiYp46GQRTIZgNK+s8FT9hP4TUgp+L+MgD38O+d5cpQ6U/BjE8KgBBnsiBPI7ERPPcp
x3kTHdzbF3B/zl3NHjy9yjIQRFag060jzI1mxWcf17WRVZoHjIKpZjLH0TNBvKaeq6NYgFoaGGP/
hbvGVivf/PE8aFcpRu7h/i/eMFYaNfAIAVwn7eJz8BFfi0FNBmzjO3nFDeR7ikxjj5A6NKvQ07sE
L1ZS4/aG4iM1qGs6Snklp1saNzYy3/3yZQWZUz3XJRUDxlsPZXDFAOF6AsePWTIh5749wK1KeEhc
cR5VT5/6RH2PqyfNV6cugM5mN8vdyI1d92RAzPOUhGr/ZCnBTSkbKLfQTBtqHYRPgOmHJ0M1I/7R
2GsgkqMfg9D9xZm+5BCyHsb3Ho/BxIoq+dvzl/JnuJofkqy83ySFo2rw8b+SK68nh/J5dmXIDCk5
f6caBcNogXMxHoBJShjSsgzbrXx/dcHeL/UqpIzoXPbpyu7T78Klfhj4rHTH8wTJc8dzNvKIO/jG
W9/KrxxTTdJW8e/XmZrCzsWJHiVE8l3pNdOyuSQ3GzkyZchmkTorWySGKR1z9WTAojqo4EGqXQlK
B8JW98ZfHFeZTXvBM67xysHrpL4KOqhx6Bt+fvkQVK7KjaIjvPZeI2LH6azNlR4JcRxzvwUbK4VN
8cEtM76R8tZ8QNab/+2+hHqJy07BugJtfZPiLJ8AtzvxvGGVQZItdyDMA5Uufq3waaAhShHF9MT0
gWNFuATDl1tMvFvrzn5vsXJICyEKLaVzM2q18ZckuePZXkH+ZTGP+lUXnRCO2wC22uzLFplVMdQq
Q0+PAAB3+7DufUtpkKDd+2RC8n3kb1PQJTY1Er3nmv6o2M8UVpxmxz/0Cc0a9nnDXzUlJEaKACDy
x/JtHaaQCGUWDibvUFPJKEmgxLba6b86pHLrrFz0nJkMBWNn4oTWsTia4jLgbAi3dBavnyKSfR2s
bi5JqhUawT1EoocAJUOKC6RgSDRC2+Uak9Gxe2PWtXMnkWKqmV8AAol+Y2fynUWkKpxfTdSxIRV7
E1XK3QtrDRshCJWWBKhqTLHuehXZrIALa1bwLydeqIQza3AAWIhBjqNVqSASzQrwAYMFM+45Iqac
k8dmf/uhshZhhixCB4sl2DxLgyaRcUx6fBPkC80ZUHarAC3lWnSOb0sSVp7hrC/rmmg319RcLqMs
dBsiHOqZpVg/fnV/gB1a/KivS6ty8Cjezl44eQ+b54/dEenMUE0a42lTQjaKuN3QFQ2cCqh9tzfk
B1+0bmtSqxJNgvIwiIrZ1SYFHvjMhQUNMkJA0QWshel94luoxZWVc6AHv/CfwtVcQHFgtDdxHQpj
ECsUAulk+z2Vl07s8JJyZW5d0WWWlwumObAsZLCnVBOS8S9yK7RgyoOGX6r1WesQ5xVbgJjU7PsD
eeJLrWLBopykXNAVlf0wC2u912TKXhrAHQssdZZuNzUn3vfOwDYT7RaGmyfc9u+CkfFY56goXUBU
q1PxsfKehrb3lsR6o7Vbn5LA9IbpGNRQADLIN8T5UZMWXQurH33Nwy6iPukYhh+Fl4PH6baNykQ2
eDeuCyarqxIu+eZVceCsmd6r74CmJ5No4sX8q9lzR1EI3k73QJi68HJjNd7ZOQamDIqiFBUWNHiJ
Fn3lGQJ6jmTZERPthCF27QB/ciCN35mEsd362eyXMJcam7rgYHb3lD59AWd5GSkuN2EMNWb+bHR8
ryAOMOEEKLGORXxbxqYNX7VMErWyGo+U9wINW9iCX/3LE0qMz7r0Hh0Ez1RBqLdBeFsiBQaYwRda
hEB/3DoCxY9Wa8pUyr/C+HWFVbSeyauEWx9jmvptgf6T+847Y1lz5c5HoVl2ab5VUPmoIowCxZVI
NS//2e1IduX1eZ0Gsdw+kN58Dq0I66iWKKef6PloLSRJFmVAJGyrGFw7LyeVnQU6wCQvOJVw+Lzv
28b1/KxK8MTYp89hEAwABPntiBi2ghcuoiZXHYugfOh+yg3xKpdIzGfyKCQCFwiNbkkZzGMaizcz
ajU3kMqz5P6OdqJ/mwM+hMgMA8WJtd0UNC8I+N9Wwf1mRP8lrrmhMkZkCkw8+9rvC0nC2HpIlKTV
YQ6dHQ2S9G5/w3F5PqUjuF7mRi+w1P3DPHxcmLJYBHiuh2s8kGCU+F3fFVz8jjW4zAqnfzahU5Zi
Z2ExiFAur+nT8UZugg9yrPTbaI9YV2ETzshNpvY57EwHUydhHeg76yKW8jkNidPNzMRUOMWvr3D5
hwSfsAjZVomlRw3KhUX4wp/UE5s+iTKwQnS88V/65QsxXqzbQwM4ooWOlInKrG5ARqiQMHO5qbBb
pTetfgWO/FUEi3NzddNydsJLop67OZ/nh2XWwWDJEFeMTAjzptcIEzacUNMqezB87IcJ+Z9kL4lN
pWp2wOF/DayKUJvACtGNHIEEySS76ZOfQFyxsblPUCsWOLtInazoGJsD80iipFBq2npg2kInKzty
/+bB+VfLMlFbnLf/JzzhKRqVEtrWfLDSfFpNaxkqsRhf9ZPM55L0QGvaw8cVkLOsgl9UNFgVUnBC
MtleH9AwVUZOxCET5jj5F6SBTCCiX/9+5rjzhi/EAQzuzQ+g8Jz57j1qnb853lXgiNOXdBpUtwLa
RCY3Qs8R4RHjNGhr7FKFhchp/rmYt9+4u9//Mrh5QIO2Lmq/f8mojQVUzYFtwUrbDclzq43XXSGf
H0NveILR89LV0Rh4zaQSv6hTXVvMPIgDoECroc0lZC7PdxUMTn0HlPnpp1IaERhCWORKXy5xFl7t
72/R7HDlWHbybxvbe5yghksWa09xuqwobeScAV9xo/Q8V5bQVIaK5DbJXP2TQfhnn3hvSQLw78DI
ldVCsSA/6N7de8YEox2JiCIXS7UvJEegGjnbpyc0/Eso9Bv3CAzPR4+BHXjM28Ww+IgJapxP23AF
dejmqyOwIY9GxgJvu3fPlowsY6yahYI4R3wW9uNFZ+PRbZ13KNs8JBw9dKHp3eQocXWEcJqzoRkc
riaOEQLIBXxMxTkqORmpBhn9pFoA6pEUxC8hHvdPrEz6L0GbylPE/QfBY3UWPNJT5CtwclaMhW5G
nQe8oBCJxBzdGwZ7IljM8Dc785yDWPOx7hR/C26at2V71fu4J6jpFfjfMeDRx8je/gOFrznMlySO
6S6kjvz6udAyqEZo9PLAzslw5ndAp48hUbbh/11sMCMZ31dQvp+F+qg/zR4jNZaQTXuBvZYr+IB1
lN1wb/m0WD7+moPicIS7vjtJpZUTkOxDM+qSTFI4oEkF5+fVNAVBK8pgwgh8/QnEhFhyq39u7sfI
F6X4TlwPUBCQsDDDx57tZKPflQqkF7x7R42RDM6bVZPn9y31togfPlLnxzop9luwZZUN4FmLprbB
imAPonL4FjxARNhHdIXkMXeU47ZHVs6VyGpXVmZw+0/Lw9svgeM0aPDBOM9yvTBR7CEa18+p4AFE
UkPls2EbM973kZBKIjTGa8/ViwoDYfPaXZ+Su24m/dIFDypH3ZTmlq8R21jWXwFUzMzzW9VK69MK
J1j+dIb9+vVoeFEoUfhQbNY6If1RDlJObWPK0AbBctuRee63qir2ZKN7ZxoI2jzG/z5NSyM9wPr9
gk0XGkQ+Ct4Rn+fSUbhsZOK97fje/vmu40jCCcHAAKy42cXK+82lLbRuUebje3vvep9cxGXXY/f/
yTwyUUhFteVIP0U9lKGj2j0RXmnr479l8rOzUexE9uak7dkdd9bqhoVeO+Iu7ZuRClGl6Pcsw7z2
KDDIXEuKg3E0cLQvXSBSFJc9/sRiPPb1lu6frBzTGgfPD069BZZJvkWzeHpNMuX44uiPW+EhGD13
CAYLqNoOwzf951zMBe/yUq8dIY43SzKR3dqFdyRcCSvnk8jE1CG+ZLXkl/vCqdUaHlBdI3FyNjkA
hdMh/BI9q3bEGwp26h37kcnT8J3+Lc6oI3kl44lVKAFNeJMrfaCXfOI6QBe4sQjzRkL6b4IgKrKX
SFHc7kFbXGVYCGg7Ecjg9ZMHlj1djjxsmFw9TR6piU2NafHRKyTdHH8bYcpyp6NSz3UlZxUIM7Wt
N+im9DROzwMTfPhzl62RUrVmYIEFKHuFZM6GE31gFUxriGrkrxdvIn2wYe8eBygw1pBAUxhyvTup
FOi3wgyT+iKxPxtMBFpMokHI6T3T4K6LoYqbf9P739uBFXJp14nEyVBh/Hr+cPLQHeXNhieFuq/t
X09JQZ8kO6Ks/qxAiQew1qvWOnk6VcrkkZmHJBNKc1C3EVC8VJQAmNc00lpotvn+k0Gtak5BhfD4
HTnYMJCFwXTAsrAW0vwqc0GTH1NEDvPzDqL08Rxmd08GWj/GuLbNUzmTbJxHtQwJmTw5CybR/ldI
ljXKMqQOHhUxkl5n40zwbPTdygZgu9jQbuTecGTTJ4cpD90QQzH27y5o3LZK/zHpA0ZWms3vMwnB
THTIOr1Lue3YZkcDrEdmuC47tjZDgaMaoY2kvU3O91hDeS+57lzKQWEyvKJAyJmL/e9Hi6KtLU7W
kzrgjZCHYUuZYzuOESisbIDvsNbLECyvOsURorHHyU2/YCp3Y3BAyXxn/hsiSSz0RvtJtxcBgHnJ
23R0ArcW/uXVw9uMw0SxR6l+u+yKecMIpOOQnOpb2vZdlGCSqsw4aXIWro/cfzInhEcxsxKW3enW
XGtJJbtw9X8XWvAMSFvGpUoDl+xZAIZ5l4qJjGQ9aPzIis3sjJGu1IEFWSk94ogR92W1AFeenTde
shGGKZmNXBPLlwtIWFiifPETV1QTyadu++otS8u0J+jyHmISSt0t0Zfd5C6+BiudlP6exDiAHJqW
BTy5PyZMo7DtuwV3WaZgeyx4L3nSx3SDcwUedTO9Mqq/TEp6GL77MLSW6XGXbiiridJqG3bmiAfG
alC9csz3jwGm2g3CV02PWLdprgn08DsvGSAY2npMfVSCjAh6E5HJWoiyt0AUwij1LBMHH5C6dNfv
ZtPIedWGotpP4LNtyFIGyi6Y3JXIU4eNZissotbZRN7zCBmzcS7aLSJ/DQMmEwb3zeTL9g61q/yK
sKTLezzcetJ9zwgfY2rb7dAc6YHb8NOq1ak/CyQPKq2H6cPrr4+9Ve1a7EnqhLc0pLK7+r4VLG+t
U7NDngoSl/7i/LsN6tPO5GVQzB66ccq6HP0Zr56siS3wxHEagiClbUIhj8ZWA2dtyjdSRHbHoiyf
dfh+xgKKUJVhntSRjq7gneNVjScpoFeTMFD3fnAENRN7eEVxDcCLd2um+uKnMl67wqQxaCNofKwI
oQMHgPMKt+Pfje3+jlF0cAC4OmwtOSZD0gdDVD6iAEI2bgV31ZNSzAKOi/CNPAyLfu4GFwKZ2smF
o1Ri3SXgIg8T9kdCX5OMPWzrVWPUu329AqiFglDISvt3daya6yP/s23svezbX5drdzaER2XMzBo9
WfPLH/WdJNtKNrnTsAtSAso5RBjj7+/7hUKajnsfGNcMX/J/spnu4tHTA1+K8rJn/QRPLiHD/14S
wTEyOjcg2tAqz/jJsYPc4SwyKB1p4S8/Up0ttirEhupIjR5WEgOPu5nxRfhc7g0+mtXMDeaIZLHR
SrPC3Xn27kgr1RpM7AY+Z7v75qGyYDAWT8Ct23xDOXljBaALLVh5beYZRs9XlWhfhKzfJryleUiB
FFrUyw8k0/tZwZSO8pPjjjUMLm0DQM8O7lC7uBDmUBqNMxEyf2Fgjjdza9p3G2IE+P+/fmmzczWI
Bwavax3V38IsIJI4Fhc9/9bnp/Jh5C87Q4uocl75wOHh9PllDtPqFLYtLx0PNI8Fb3znBJAqdSb5
Cq8kgrVx7zupq5F8uecL2NwdBQvvCKAoSj7wbZGkZnQyDGoPHvpRpEAx1TN2vxPQMeGzfHLkx0LS
syF57D40XUNbqygArI71jvYy/bAd1Q4kLO7dgv+qFKAfowVDYLBZlsiqnV+LzNXtorjhhoGFEum1
oDzrqCPMhvAJX+lQuI+ZoCTr4/b9z1PKhkLLy9yO8u/gu0kVeiIT9wy+sfPdpofuyxNVtV9+MOsG
b20OEEszYLjPZXScEsHcaZGX2Bt9OxhITffysGO6DlPMHz+FhmRzbgwF0v/IsTPsVBHWzFTbcC+v
XJz9AN3t1w+HBqaGlaj9113S6QoV7z1l935iQmq894FYaJIfsO41v5nkPGRj6nPuMv3zCXpUcaeU
WDveqFLD8L25QWsk4kmjSz86641ChFUQD9BKdFgw7C604cUk2DtrUICwNQoVs0rLfKRUyZEyxKjd
6TnM0y+XPHAsE1v31OjBM/IMx0kKN5MrLzIu07mNKYIc1pYBcCQBes/EJmVnanNgsk1VrM1RSV0J
YF3+n2xn5nHUB5QkOvHT6COKBQEpEam1aT/F8BPaD3FCEySUVEg9Tggym3prg3MpKetDbl0pZC0B
qP5hsTpt6AVhPyxilibxPB5iIcLQxNAtOBHZw3u+5tNiBQKYPVIAOYfO/P089alSAN6XJ5aIvHVL
NZNfZji/esnb2jcoCXVWpm0Q/FNMncKPwNQWpFwNSOQySs3iHJH8n14waRUOnXPRG4QMtO1imYgY
cuY01ojptx5hkwauHLSoUbnDJqg1uoU2nJ7HM27Ye8lcqlnR8Pa44TtFiQe0ax7iGCoEB/S6FTtJ
9yFnxdVhzNJyEaYprvlApT2gJIgFfGrC8xE0pzoAe03XJa3FypAQqRvhMRru1usV8uQ9H6RcOTeB
C4p6wAQPgu338cQaQnmVhN/1WVMF+MjW40IAkFMDliP72oKaBL+ou8tsvQBPy47O/LuGgqly9LXf
MvM+cJlkHl/+LY2xGPOlSmW3O8HO5agUK65vIVceYzXVrZjJOJfKIeATHwfGd9+uDInsuarHNy5h
LXqSXtpnfXWimR7z+DUlCkr5U9xoJ2SuaS0n1NpiFpc0UqvO2WpmBr/aHdyCWN9XvsH99e5Vy7Ju
xYpwraE9oyqFoLGtPeNgHs8RbVhgdYvcL+JOR7xRAXo0EI49Pen2sQelfAz9aClF5CM1ZfahQK2V
5wAOgs7UUapIhin44ndfB1SfwRb8JUHjoEOYSb2dWsYt2qyh2m0EBoaKXMpTBlQMOxvlcN3LtS4R
hsxxwhqt7xKbcsExqfEOMMD/4eDCq8CPhNkyFn7GaBkNOHvVXJh0+LlCvZdmrYhVQbZBterGT5Xz
YhzPFPWFAWkbI/B9m6/OaUKgu3x1JyxzkkmICnPHRalXJVppLDyEQHBejWFUVgDgAZKchuFH4krV
xqCq+w0VyQIorgVaSWsyrf+A0mCnitNXHL5Wc3+WFhw7nItE6v1w0HAbPSjc369QihsJgIvBJiDn
odwSbNQHtjsKWOaWCAAFB3eEYU7s14Mr54YsPWmGtvNYi6jTxOimbJ2Y/9UcNSWfLFjCEhPitilR
HEFSpn88PLzMxPFzzhvDHbNrgZRKsyUo574xgi5pkZ6S7Mm66sdINnLP0NbMtRY3m27DVGmfFJ7T
E/31WnvHxHC8KnMwF7u0MqcslPtkP9K4Acm2dRjKX6QQCwJBtxeGNx8Wb8Wu0jeV+sX4TypO21oK
MjlUed5fS/LOoh5fZuDIvkzxmNyGwt+xBQa5OH3rdrO7FKNyWqXlfqLFIt9HNgywb2Wtny/4o9vU
gD+2GyipUO5JV+GcdIa4knM0h9A9gj8WmvpN7stq4m6+y4hbgoR5IHER4O1wPBBLwXbfkbaihzWl
j3Zzihza8A7kpwjwL1rB4CSO/PxZo/KPUqCLlua2iAYR0AM1ahlOVAcZ0xCa/lUYFO9z5bygHXO3
XsDSFTZCxqA2FgvgdDK10HM0x8yVZ7VXmbioCIzRH3LNxW4/4pCfCYNLCWv44XBt/PYhF5YssFkp
whI11q0WHbIK6UKsw+qpKo5zeMoYE5pdhMxS7T6F5P5gsR1dWtmWXxQm9y6VNXFRXUI9R5uM0spL
Rn/qmpeJm/wUuWkA+bDC/dfXVFnWl6Qvd1mKp6S9XbnVThuM7wwbxjZ1zN7xR2XPLJ/QrY5AyfpK
e/NDAkrJhpVy4ONKuPKO3frs92twKyzGroq+OkyORqzIVMcDvncjCiIDF63nTGGRAhRnAQm+dZdu
uq8cRXjIeuyXt6QL/AoX3SYrqsAMvhK6+4s+qFK4eURwsfWGnMedUv1J3nZdFcOuMmhnco5nJsrg
7BGSOUMrj/HBLqQhZQ0B1Pgvj4EdJou7odHaHKKypFJp/FLbgibCiJ3G9rFWvwN42fBRVkACO253
QjYapqcleObnJfc0LmKkzi4TGQwTHVNzmsUmjOBXPOQ53mvf+Dq8c+fa2Ffaq4wRT1Dm5a1RCvTz
qTcupKZLu52r3OIEl8dJ76wvyy5MdFRYiHceALyE6hrqADYZRviZY/V+OF29fMleYUqtGxGuT/11
+bntJESIPRo1EXBO4vBY04eHA8vqHT/y1RtxNbiKCiWb5afdoag8KQL1kdrfywuFcXxywvZnyuXV
eyTuIzQXPLrbcYI2saGWTtkq9DRoJ2yJqhuXIolYEMSbSkES2RA8RnOoi4+5QKwDYFgvqXGTMUKz
bk1Dlk7dfpD5u8PF23RMv6lFC9o1WljOdalyi6Lj9G71etZ6knAbxQb9Sk6RiH3/AdD5ZtobFqqj
+Gg19Pk2O3Hcoc3LhbvH5nxE3exRtvn16j3M8sjYVlEey/Nv6OmPgK1RDBSXhIT493MUqJFK8zd9
+JxMIbiLGxNuvml6lWyAI1n56qWgzivKIC6U9as+wyqi1Azyz6XQrVHSW5F+W+RFJls//+nlm/aB
TEu6qv7WlXOdpyQvG2xcORJBnipSr/watTt0FYBazoK59KcuYTwTV72/Xq9GGM6+iwq/Wlagxlfv
v3Ckrrk3ijUijAlZCJFz0rw53BBfHGtWoz0A3vl7iIOPTV3DhrZG6qHf5EMf6si0OcIvm8ZGw4AW
QOME5Ot3XnNR9G0ViNeZTW6+xqc10huPdf6kMld9UxkzqyJRvSzAUrEBEXaedtUHw0QJfdCWDUd0
RR/u4n/Q5s4GkWsjrwz9Ds7UGiICo2ZpZWV2v/jEwRwduqRoODW/GPO4JOKEQwuNJQaKZlHa0ZZL
qij227VmvGbiKMDKpbyRRSkEntv1YVtE/x6+lMbTTg5ZWUc4YVR4x2NUROi3TKjlNp9BzWZT6anA
Uy2+QQPaIHjUVRWZaI5ft7mfVlrN7PDMkK/HCQkMwygLDib2wB2IeSoWkAG8iWw8FVnpRprw/E+I
yACS7p2U3Is8+3Yt3/CfNLZHcK/rAHocUIUKl9KxJsExhe6sYMZS3wYq92d73APr67j0ZjOjezUi
Ebp+++k6CJBt186rvBAqwa9hIHWcCQY+sJRyBAx4dOl2psOE0IcBIlp98wZMUGfPo3cp5Pdy7Hr+
AErP1DKC7LR8MfO9gsmeA/nSca6lKueEKF4MFQHcK+QkjWSXzwa9nlDpYK5g6uUPz73y294thbHa
nVOlatGM/zMkbwFORU7FY1Fh8RDvapRZwD2YenSrUOFLoalz+30p4gUVGZb1HUcVTVF8qJVnorQ3
tIu8QyOjRMYZxGttvvL09AoB3dKiL68jT2Y7XyjDVUEqHtiI6lZBtTiFWKgHYfINpFXRf/wz/U4G
xEV0mIZtjQnbUS2XWD4ylPqvtkQDOoPwh0wFOPRu7quVRXvgSI9SJgIREM8suOrImOFbxfmHVpM3
7g56IRbmzXai2uZUPrZ6qSG2xeRtrMKmroN7rbPQKdlteCK2WlGcXjCNjOxZwV8P6ENDguFA3BSK
GQz0Pz3UAuXliOFmvsobBdGoBQtpPobwBZji2v4MlbseoiiquvjjGTLcJmXMe5MaJjJsA55aVOv6
zTYhm1vxydal0TQDDVc6s5SVWOZqUd1Je9Z8c4T6CCiTEc7TM+DFn9wHjb2OMhnCgL6y7A1dbnth
glJfIlBLhS/KQlQLJAKoirMNlLt1D7y4cnNbakr8j5GlpxzkJGTLRJeXukqiXBd+yEX+icBC5+aw
+FhXSQE1eM44U4DzMSZrep9+KdTiSa12NQ+lDMMEEy+KJhxPx9f+h+Wb17JbqMb8NMVuc6nnq8bU
xrn7WkMFnkc/yrznvttt3T3TypzRoJiZWSblObLtyB70QomEmhsYTjD5NkIqbGKQHhTYFlVrJIpC
H0AtPUaspRYokaG0IvVqjgcTVwDwkUGX0Va93gyNcV+0sIuLdnTe0goWv9Bz8+esCF8+QEzim2+X
o6DskZOFyQcdXkqLXQYjKP/yjmn9+dhejBug6brVQpaCRhnvc8eqn3Wgp5u+NLr2hyPsWXqM6Hpg
XIrH4yVa7/oDIDggMbHqc9DKuwrWcRRxqZet3V1TJBiNdxOmlHlc5Q1dZZ4oZn9/Tp10PTo0ELZ+
WuzgNv/KObi8W1t8oqFDJ0lX4ftREWFSeboKa603P3uzOq1aqLJDJyLDDdNgqRdl5q65SfPIacn7
GIf0dZDVo5WzozZ8Ue21vkaoOe8HVMBB4oSZ+UdTqsgvbNPqNBqen8vaTK4y6mLS1QreMp2apGO3
jPhpveO7iFKkZLXG0fZxlxy+O5TS4iCnJvMY5fc+p+7yF+kLzHK1GbGswFEd/ASv1MrVFPQCtp9S
zcDG9vhoWxNgYynuso6jCOn7UcRNO8HB3itfNnS8Zbd+6cnpAP4h0B83sT8nf2+vZbHfmPK8fc0j
Eu6HPEN7xeE5lxtdpgpNs8lUBtzztdFF2zreQk8skKHwRe6yUz5XBTCIiPdjqXgxr9yw+omoiuzi
Odg0/Kci7yL6BvJzSO020rjeChbB5xXGpZPbFd1jPQEhorimt5GFoQI2e5a9ewNXuyFvmhrN/4MO
Ri/UMMSeuZPVBxnHsPd+fqMjViQC+LBLEWas+gFnukTMBVHus8HpD8rkDO35Aa3XrnOmoZkvXt5m
tetrzuoJxprcaMaqiRe028fyaHJcQzBpr00k0ZW2nCYltJehEG0mjAVX5zvxDBI420lHbkCLoF0T
MJcHI9TEvfJrqK+84eh+d60IA9E4ErCQjkuXpl9gHplNSpWf/mObB4k7WX9ALuwV5Tlfz356Y0So
gKxzVVd26bePIVXbaD6uzcWyYMWrEzC/V8W0pSKAuuRtqacYEDopQR+7kI6shL0Ib8tDrYqd/TwJ
X+UV2H1JAoJJvdae1xYVO1LTQ79M32IVkQPYKVxXpiKI7adyZrACIFgftvj9PMokzMlG5M13XLYJ
HMOYq29etLUc5qmw2nTLMVpMAnzsLbYR8Agx1OkU3u36lXoaPPIoVo60Tk8aiN7Gwgbo2aMIIeLm
anNa4j27ZTdTgwiVRpcZApjjKI9e/Sj1V91RAbsHm6MJMXVlaIT6kJuGGw2XVdmhg0eehCH1+23l
Rg44xTyz/S7J4RDhjLXQE2MJE9pQZxVMyujAgQcBeqKK+CmyGioGZ8GMgHHUkY+7B61ERxnMQFD3
KUIztligIUoyG/rZjm7hP/C4yROxXWxT4axoFZd6nqaQ2RHl/HVzZJLA7pSrRMOACY8Ay/6l6cUz
WAmo2OeMxaE2Jryk1TGJ4y0O3+wJZDm2Vc886mjLsTWmz9z8fuCfKkaWwhTyQpeJHmI/xMr58WHJ
+XEyTgtE6DJUNR12vER1nSw5FY3XJt2CwFsRyM/mhxpI9zMYPrINLO+BtkuQ852lB5uINHqPMXQ9
pFvLIEy2vC1VEJ20hp6csYVy4RyC/8lpiyq+FupbOt4iTfElidMBb/dp29lM+zXA3nEPO2R9/Kvb
LLAeg3VJdZ9e8scavKH0yReFPMx3UpXf5eRryRlNnfo/3UbnFg0iBIPhuXKsEwXlfk2tl1BbJCyb
3elxDG9b9LDjDmtua5jxX0dPmb3easM5waFEmlK5J06X2UYqA0XE/98DPpPKs3VpMGr6ijiaw/ET
Hgerg4MipBhakaq3A6X3X6pUwONZALcDDb9xZSmFrEuN+2Mzro2HON6JhvU86ZzaPTc0w3zG29zG
7n0WiWK+KOtaRd+EjRPYdT6W+uAaawQJNTRUbZNrF/W8lkfWWYUHiAr8n/5AOU/3OcakGFXTtAw5
pDimBzNKjAmBdVmrH3v1RCfFKSIXg9mHCEZQn9F2vqcY9rcVQ/DIwuAJx/ezhIyEIkoAwhVGLaKg
6FGlc4+hz4Ib17PpdgWIk4NIOi18SSkdtSXOmOG+cJZx5v6pyDhg6ISIkPpBLlNR7+9cBImtm+iX
pmO+pQ7b99Ncgs1Cjm3/NyJDKVlKdiwD7Dbf3SJnabtql6XPZyXciwZQTeOh06lotkjIFrU3jKWS
FTHVrSFg4HlVpslmuTxml28h0dcXtazmpzgun/omw33F2eTsbaZfBrk5/+Zmi0Z3zTcom9pEV9d4
y5199M8PlNR4YEoYAorJMxPt2wZq+bX5iOzFs8s2pRpGVP4WU/zfz0ILIM6keA+M/RygcpYWp0GF
cNYrlebH90N1XnYyQd48m7C/vVEZhsEod3cFezre2ZJ5XklUsPNIKGPWdzBmpfrJWO2giq5Q2FmR
6nBuUgg5P/lzhQP8Wn5fME0/xMy7yy6o2d3IZ2+q1DYi5Hv8/pTVRsr3yZwlKoKcWynBcSeI7Q1p
0nxIWQjYG+8HqwI+JzsJV1K5MCaUpHusf1IQoQmAa+BSt2zRTe6OsWMBbyWA4QmezaiHrWkoEWfa
wK+S+fhJQHAo82iydTLl/U8y7nN165upCCEzfYWpDH8a1T4rPPy2dehhoR6DWHI+brmzF2JjqDjp
uwq1KU2H4uzcN/ClXorcPjMd++9VY/6ttuCS9Twv285Q+NByenzWKNCdDGrBjVAtDr2GWIPFWy/8
s3Wzam3VX7IBP8jlWIDZaBguKofWg1RAQMnij/ZslJPr/hcLyBiMtVkogGIRulSvVbjVNQO32Iht
vIPBUz4aRD25n8N4YIj2y5tHO+hn33vL7YLTED1zEfLp59E9qfS1LucSOH/PycxBwEm/h38d2/US
0s7TzrXqMBlQbeqwTCqB6MgUohY5EIn0WSUUs2/GCIsM4Hj6dYoNkc+Ot6emV9vu+VwEdvoVCAyJ
vXX901qegiY3qK2aI+fKSFCA3pBjbwRkm3/H1aNvFHCxFxdLpYCCCr3y0VYh0nZqoZ4nVn9Mr1UV
Vt2yPJrbf8d9bUjPXt7Y1FpwO67F3WquyP1ARUFs1me/BxsjwTzqCjCUYnxUr2r40E9ZCjE7A+pL
nmQilsCpoz7Xd1NnV/vAqKhuX4PDujM6hCkto8eeW48/Z1PeVaqm5K39L01ZJEscHbjCRpGzVCXR
dURWjeGwMpvugxwu2tQRYXz2q0YZeBLD80dxAM4fZa6hyV+8I1Ks/r0h6HmMpwqh+gYUdc4W0Y4b
8KB3MiJiUXG2uAJlzlVxm0FsJDtRhSwnLqm68xw5xGEDfI4MAhzk1fdEa1MYdC2FU2XItlokq4zq
RHKlCS6nsW5lLQ3zdiyI8jGozgZA4ru5tBBotp6w23/QcL8wzalf3X/zgG52hnoKVtUCrdngJXZL
FnocdUXMp+vThFmF7/D/hj1n+TNhC8HVqslicjlxcInBi2h44fP7uHTCGPecXHSpNXN/2C4jKUgt
yX/i8GH8vEIwvsbml5mdN9Ok1sMIGvyDIKO62qgW6tGAZMeHVATv0DPYe6ZgDV6Cx2fO4g2kdkIS
NCnXX3inMne9wHB7S9bv8SU11gSJAl5LvBRjHW8hFliQkvmj01lUWXKhMhHp09ZVmNFPxA7SUFt2
31BZprCZxFYtwubedIOvmd7L6f176bcaCiGLuyIyeAMvIATi8YNUkgfgEnDbvwklCArlJ/NfZ6N8
8zo7Squu0eopQPvixjLFfMysozYh9vL19gH5xp8wccroCs9Ekd5oZ99tC4otjQD76cmFeH8AWmzo
kdiVMFKepdtbLsrZkyMwUrvrqkRHBo5iHImAzzNMDzSJcg5Qe7tqPi19jKR7eKCsCqZDHaQGSgWM
+k8AMv74l+MkmoJmXBJLv50a2Da66yjjd8cPbzfYlmZmMDJBxaM+BccbVrJ9Q2AtwJJAiosqh39C
xTRsK7DC57mjS0xze+LRPaKKxdIDsR4+AsGiVMAjX7KBKgMzPfzelr5dJ7IDp8w28BhY+/0RZHO4
OLsh6WTruq1elrbysL+tDrCPkX+85K6L1Qk4IluCrx4GxNw0Sm6jv1a9l4b/E8vot7DZOCruMQal
y6qRGPIoeSmgMlHkH8x5hlLcUCcivFwXnJ38/h4O1Z34lz5z4qqS1dldsKheZ6nmZ27II0fpUfDG
x7V/rE9ywgdJLLjOZU6JF9LdMrQH7ljnaSiTaxat9rzT32J4DAPuvLgSK/yAY6/ioDqLAkXIMaaE
9rWjUptmqTfSAgnd8zoizWHMyy9G86yztowoXHvAXwYJDmvXyPO67uSMi8dAA1BZYTY5ZQSHVnn1
T/xTSkPATZY+0RZ7sQNRcg9g75IwY8EWMaFJT87wLQqLiBU8uxJGFVuzyM0/Bb1Plcafo4vSw7Hh
oWa86rbxdOJsVid3E+WkA8mOSMXbWDIY3JLbeqXrhqBAZ3WxhWLTnSdx1s6BFMIaGGTa44aXWBRe
jI2PPtsGEKOu8t3RDuFWMXvkLLX3fiDC3NxwuaZBnWagZPzAt4O1PO9TipiaIYtQ9ytJIl1U7kyC
UzBkB11rik4tmZZG2TKcjK5HWcC/egNV+nM+ac2KrUs5cd5UkH9ztYmip1S7QJeRWY35qqPBebJI
Zi8QTBYrq4cIBMTELmQc9EavGsqWmQ2vnH8wPHP1ukpKY1eONBozpkMayaSW8IMzF5PIGuXL/s0d
7kTjViD+VYOdzuLJDayta2SlfVjRikieqIiPdRKXiUqAGBp+vB1RovVhtHjQy9mUHbETON0Tac9T
FQnLNwA6sazLgWLJ3txLUP8OEf9GaHeaKl7o9yMRz/mlnrTwL9JOYdqTJn8lQBngVXrj4cKRX1zZ
CZBFWnLNR13AUstE0QBlBq9xjCts2qG5fEJYWhTRaRCBdzQ/5WTPBnsRZg9ek95frIvIAh+uuVSH
VGRn7d3BK8G5NYZSTVN5M1exa8hr5pRhBXv4RagP2Qz7JIwjgOzem30cR7MjS+sjZaLV/Ajz0sDW
JhKfXwTqTA2Gko0qeXlT4laDuKh1/WirzOumpIQONrv5X7Na63cfLEUUmlKFnkJGbL1R03Rk3ghX
iGbl1cTR2tVefrX4FmDNOXkOVQTN1xpU85LjTq25R8/4a9H9Pc4L6IhryvlTVdVTWqRgt1CUB4/N
CHkF0kGlCDJh9KjCEjSE63V4cwJNs5QV3NTFH7bt9d/7v6dpOHKSxqnFzDK0XXRlHZjf+SUrz9Oe
qNRj9er/Tqp3im0TBvWe4BtL8QoRUpCE6U1qzdhu3aqmEBhcyMPIF/42B/yQbZOttCye5t97lDBE
6jeNRmnBuXacvlKOtM3WFih7y1JRIhm43neo/Y4gW6EhghZT8w/2H3cvfEPahy3oGZ928VMk7MCH
BPOyEEO2KSsK7MS6BHgp017T0kxpAyfeVPYTSkpG5dNd8Jn2SF81dZ3+BqQW00vs7xOM8nOlhgQ2
t79+Pk6lI2xyoiSKtjM3mvuD6fULR5BWJyPRJ43u28bEDhh2tZ6nnHeliJLypUFlp/+pyKXlDL8z
Rb+dM3Kkp6jb/sBjimty5CSTdsWlmf/fM+DhBGo6xXYVN+vYrjf3qmvVoSgyc44t1174cAnojTH1
0rgiEP9aoQm/OxQNNhyNws7T+JqDhcLIeABEUHN0e0qYqf2ZBbb57XQniEHMg8YF2cGhAnKqdC17
nXbqkvqox0ZWDMCfKXiyK8txMFT6jJuXSBSclbjgTWSe6sBNDTAywI4UE9Tfp033Z8LuqIP4uUYI
ywyOh3L0nk7meal5gn52HZcOJN2RY6RZ6jOrzkKWTZiBNuIQgCiOiLx4xKZVgx1f2dMdgcWKWAYe
2ALKj/OJrfSBJSb3KYL05R6YAkUbueUHw8Xpk9XE4LfK9sbh+qJGOyaC6gwwS9PiQyFKLd02Q8WC
Ftm/aWnVbAJvWgZ9mZE6pHLvwRPVsTnGoS7ZKTyngNlOCMexR3pKbpAHekF++XcQhYRViz3tii3y
88iACazOCIoQ8YsrmTKEXTyqPPQyCVIn+Eb9rRdGG8Ti8cnMAV5ydx5FRyY1on/4mH61oEoBxDs2
F7cX9pt5QL2vVP5BHvHqmiZw0rpTmyh44gfm8sqa0ci7D7RoiIQ+3FMa5pOZyUeFFVKjNENLKzZD
cCoPyxl9M8NvJ8zClGKkaFxxFmT90+YEnOKRSHOpoWkK1TVOX7arS+y9ySjW5kyw3Ytw6mckE4hu
eGmCIE7FZAAvviPDH5xFZufMv57fbQx1kGNPz9WLFSWvZb3d+kJ6FYOiMQzTmeVN9yUd8O1NeSup
qaRH+EkaGLjdxD+v1ji+naWhc5WJNX6w0kt3WfLM4g7ohM/cK+ksFsU8EF/WYOzDYN4lTK1OlkhE
iNt/B9fFfxYCI8AYBxDjYx02OrUfTMbVqwL05ygdYVo8wJ0HHAz6ikR1vxM82iiP1IfADf1bBv/k
DwE57d9OFM6uYNk2ymmQxoed/6NG6E/sQZm7s+7ApgSYupXaNYs8K9Z8/6SJFDOkSiA80F3ZiXPa
32Rt/mXRYHcYOkNmAQ4NjyguqgYe+vRfSUnoSA8jzYr+ups27r4toAbSyoc7gy0wkz1PAxlQnh0Y
r26nvHOREnTmIiEp6taFHOIX8ts8TH6EN3tDRrdj+eFlrhtUXk7Vp65lgFou3BBR4rxMYhGxuzfI
595W5rh0xY0lKClJlaIl012gw7iLQWaE4nwIxRdRsgc9WwRaGzV5NpowLjvwyMn3D/tMe0o1+YJi
B0UwNJ7Wst1uzJeKsBs4SEx/KkKdTlHXvbuGbDte7PNrkoGTm3WLQMtGf06i8js1j7m+u41i66Zq
9jL46lBi3IXx4JY1XHgK/wUBsO2ioAhhLtVaGcGBH+F4+MrSEKSBkWrqId607VMWU/YjKTWW1hO+
N/8OXeP1gRk8LTQwiMec2T0OHvqiofvVUfebcJxmPjZOWFWVJ3o5Wmn4N7C+6Kf0jvv2aP9yRpEq
ESbs5cr957RQ4l7jLzeGJxKJHYj/xQeoudQyXS5Mi+knjl+8IEyId0zd9HEIZcc4wZ5F5G9C+sUr
wmspLeeCw5vGiV0oGhIfJAGCRsto7xhxyNLloqAYjlvQiLVBkQ8bErfogzEaUz06v9Ma6JHxws1p
9/GKWKVGjGk7I5LcSth8Kuc5uTSVA/JhUDJm5h/VnnLEaq8zjOduF97amWocj/BQ7wO/KY706xwv
Gv+YSFKaB1uauTCeNGzt81dmMd21eZVcyjGTXR9lfCa8k0eO0yDbRS3lizXx6Rt7+K1Z867QWvAS
WzTSBWMyPOeiZ3QSoTSZel2xudvgcPUFX6EM73cijrOKFWLGaaX0r63Uxf5I2QOWHi9zURhwtucU
4l2pHE7+m5DP1hV2CukzLDMUPuszOhe9swlAi4oO1yFtbqvC4RHw3HI1iZGD5Hckest2jVXKtB7H
s/T8KEiRgkfIZpAUXaUp2zc48BwqNUKM9RurbQuPBKYaRglQWq2MsU2WZ4Cyu5aqPtAAlfKuuURt
O7HjYB/TRpe2y/Vy4mLSy4dVKHiMN9cDlpeLYfJyhdkgT7kxjm25X07me2c2BPj21Zamcq3yY6Xe
LOgWm1gcO56iqPPspQuYiX7mlHOft5fdQoY2aRqdeTm6kLFCMetRiOo0d/B2mSUno+naMazUa/qd
96xDQwOTJDT3H14uayXqHsNHkVk12j3G5EkeLnHObyCeAm5D/0J5CcqTAokRPqAaBr34HoBpMKOb
JPJYylPRuHT9LCoffB38WPkI5Le2hhZNJ3fqYBPbS+6d84iznqHeZ75g31Sn8FYRnJ37qLZmrZRf
5+N0XAYLARruZbMnRkH8jJNFF2Mdcwhb/wteab3yfBt3FCCi/r/oe5i8XZNyow0r6DdPly/GHnpB
8IuS44kJ5WbHdTdA1FTjnD/c2cX5r/t6eRl3RdpmgH1ucbUUygslPHfxpz4KTskRCMQmUUEBppxV
+Xl5D+q8dH+SvYOdFllZyccr0GQO+i6Hv+EwE7ah10GqPwuD0oTyinCDr17YSJWlDyYRK6HzU9cU
/9O841Jtzdj/rVym8/JitpDSTKghiwDEFkWVN2XA4wh714koxVgDe0IvXZWKwh5KIvHPiDf8hXZT
Dt/n0beTVXAv5++O8DFP36M3LeMdo24GrajKaQ3pySoMUa3cHl4e62Rnh7At1ASBeOHBQ3bOSeyV
hKcdk0dxjDhRfPA+UbBO70clkbRSIobV5oZae8Aec4NYkDNET/YX56d9YhFnlAdrnkEPHWjvKoUY
Zmd55+yekiVRtCNdaoUFeN6EPUx9MEl+Eh6YLxn82L0w1ZGQBmscWgDCCBIplhxs6RWZKK4Y6psf
HKZ3rJHusilvOKB8E6MMNjWteMgeP0OsuJMMpdq/WWgQaSfQULynnKR5vzhqGGQTMo7J7wv1YxG+
knFB/azrvUCEjLJk2l4Ih2arDICUW/12jWhw9NAqhA/kSJzENVNCjeANWipcka/aX4v8YjZImbLC
KuCfmedT91WVoo4fZbfyTAtGWlNwK4Gzdmc8gEx0yGf8DYY1yCu+4C/7XX1/0dS9AlPmlMQ2DxAO
2eBBBcC0agU19G/Y3epL+xrA7+kHAgxDElmoFUcxLQDrj882ge0pNcr3g/5l2aybLqH/TnQnlOpa
c5OfkPL/zBN0GIhTsoFDh4PUw8ZfrZ57TNxbovM/ufwtDm6lC5ZtbAjDsKgx3cMumWcrS1GUuVfI
OeRcOFA8Iu7iE0lUHX2KEFkezQjI4nzesGNDsUCIlf0O8Qhi66opGPKWrjp0dvskNfWG3XfMPnk3
ToAjxsl0WEuElvgU7mXy1RsL5b+pDjDdEUI1xORa/wzQo2lOFGn6ITT/XUMLYICT7t/DzsuzPH9z
35fTvH4gsxoXwNY5oTQqtutLgxSmWKaqxnx9WNxvts/tfau2SRjtZj/oC49kqmfgo+8RzMyL8yzH
gSw3KJBSS93TSWRoW6kXDipLVZpSMwAImAaEd0yj3rpD4/ajUDn9cDZiJab8ONGX6DBjP+1kBDgn
mVT823e7vJImfb/cm64gC1OHsV7NgSuJVS5IBybbnGgAehUispo1hLeKkWSWVbiGUWF8zrBMCcs9
w855flGVeuS9IFIkbVZoaIyS/D3l4+Gjeos10CNStH9hwTteh6e4QGsii8RdGzMzA5oP3Fsq1Z8F
3PW7Nk0HMM0ftCOVX3Ay2oTJz5hRYT7sy3C5nSLXs+4NKN2nsA/ZXBnC8n/2oilwebsJQXt2BUtx
YJyrmRf88FGsIoxmpjowfyp1F9khR2ZvBN1G320FGUYNdwGNYcPlK+Q9TSEl94cPNE3ol+wutN3S
ObtH2UzDleFcKU4RC74XwXzjJ827vIj+KXtpSWlqqP6sihFI+PnM//4k9swGzVq1FHJ18bjf+XRo
MMQMuIDESshFv6lIYDSjWmOJPJOfVQketHMIAQODSpD4i9LR7RF4F1wJlSl481oBLvXg5rsa+9bn
0np1IObgJWcKs233EFH0pqqJfxUsRPJDeElG+ddP8T0xsQrzPTCtYnZYFleZ+Uu6b7CWvbs90JeG
M+1EbLEI/Pa8jkqUMo9LdmTTya2fFGUT7rvkjfAtJ9quZdvDZXNR2+DGz891bPXmky9PXVVcQYbu
pdczri3GaC0xqoJtzOc565glsjf7ZbY4z+T2OM2SULHHd55F2w19P8rb1fC/3RPd3oJPbNdj3t+G
P6UrnQrfRiunVH7ntUg1IaHMw5tXEGuaH8FOyvoScwwWqU5bVnaD2ei+id5esvF93khOxtmDKnNk
LlmevRvkrCzvlm9xL6WadxuPalIQZ4VK+7Yl8z8O7UgZvCpLTZv6uRTa/2BLsiEP1T81w/45LL3j
5jIp1aWCuGXbWthrL8B28NNx/KFkvSHzmemALed490SHqyvpZUjeD4ZCUDKhYJDHH1SrRJCb7ROI
xw0nrvnNJRHTRbtHF64U3d7neZGgmJ54yi19AEyUANx/QeoN3vQRjV7WVWEQ1hJmIEUxCOtVoNYg
iDzlxSw6m9KCkuNazO0AmLLkk641kpnwcXJY8XKaIL8+0wDZvzbc5MfwDK0jrCfxIMxXhUkxR2Zm
2drwR6vFXQwlPBH4Zlmqt9QZ2tIjYr2ws1lT6GaYGMs2UYbWVRPKI/9fBJJ7TP+w2/18PQBxHhiv
cRRJsI0YfV2lTCfxBylJXgdnjyBuMEHLQiUvTrK+y9cZ/F/SnZAN+4DYzZMc1gsACPa3K0nxjSrw
eYd0ymX1NDxv4zrDhP/6V6QAC+HC1xQXTmQ94pdP8jiI+IrX8QNg99tY2/mmMN8nYG2kggtTpUjN
GnrqnugsNUTbPgweWsU7vFERZ+jgChGmzTl6yDLksjn7e61rqhVlcE5SMhjUEcxZVpQCSRtHL4Iz
z/P7RZvjTLEZ/rcoG0NUZ2uak8iU26OpOoB8vm5RkZvCuCPKpq+/Y+13LkDOupXOrJZW5gCgrZCh
gc9fedXIMVkaHKK7InCRbh97+5iAyhgdQRbbzfKBZuCl1/OKhz5y+4VjAx0CMgc9kV7+lLrq6uzH
Be1WUZDBor3eHLC3/1v+XKdnsf+HCfccGmBuQpuAOIdm3DqrrVXLuSqWL8nAu0NGZrsn0XbsdYbb
lXAInGXTz1hJc6n02/+bmLmFLNIvHNcFp0nJ+j+YDUmmXCRyjHrmbk4ILFnxR/nIZK12YPA3oVWf
tjS6QBBQTCp9NW9S0csRxiOVN0oCXoXgeqbCFLyz2DPDjymAS9CPYwXb4jSnQ+IX2UMzz+Qo3X1o
im5bEckyf78CmFyWsec8WuwjXtp3I/cXHaARX0nZISfsEByYGA9M/CnUkULQmNIkdwRBm5d2N4ip
hTRMBJA3VQWyejaE3o0S6E2apu79pdll/ArJ+gTonPWTbQS81xI0GdCmQZAOk1dOGrQk5fohz4NU
f0fwnh+ynKt6R6Y8vQeFjlXZIID98y4/JdUx7vBzbP8k+ONYNpZ/qPvQStq+DBjzCDKwooIl7eld
gQWlzlCEJiAvYaj+yVOTJUKXb+xM1C1wWmEa2nHv+dOoSHdfhobg6iPaMBBxh72gX0QiNVav36ug
gliPT455UvM04ZBLeXldIvxaQvK+t5ASkhJ+Hd/Ni85ldetR7iaU/D3qvWWV25DNSS6ZotjqOCok
V1UjKj1oOR5njqSzHKO5zaotTmrR0Z7dM/HeO36LrabTSYI/UVVkD3EBLz4FWLAC/g+2vErrkiga
JKKSfAIeCXUrs06SSLFo3bXbR8bC0AdCv1ThMbz/XlTj4E1Vz3ztnZECVq4N8Rb/v+uZJO4zV+vX
AKi/K5in6hHN3Xyz3bww1rtz7dWUyYQCjqx+EiecyP/1YY6JtniQUA9uKjGIGQEJCSVH3T2bQkK3
scVKcye4cV5Ly8A3whxnwr7iWOzHyATgfoqRWQ6sHPjeM4jgRsuVrtCOqYelcc4Hp7er8atvgY96
h4M6W5f3LlJP9kKHISw1ac7BFTvtksq7iA9vBpAMPj2cGQzfKdcs0rc4eJad1xpL8Y8F+6u40Lul
ffFvU60EGxJfrG8yOqTROheZBZQhwqMYdR6DGIQRe1mcXc9nGFgPGh37vibsyBOz5h6D2OwYTqwO
nIHu0EZGo5KjtdQDNgd7pIukJwbnUT7M6reOWy+phObdIhjb/s/GvIIH1jdhwBDKayMn40aWNBmi
t1yujgYjJctmTSQKicANoIzkPtmBYxQxXh2Fj6zy1uRrlX+KDzUWYXyzmnAaMSfuUhyxnLp5fMKU
g04TQxgVbk1LGCoggbLHHLL4IiO9i16luY24jzis6KqH4vHv6+jaJma9DMoUrkI3o6jxBDBGkUlG
GOu3QDdlVPLma8XabdxHy4rdu4a7Tp/A8JmDyPUUZJotJaEpX38aCA6GVdPy/dI1dzCJTaKOYMJX
TAvaGSV0Ty0KjHGTiXg74oQATZAt6z0jwhCEGckoK3+1ALU2gKQETQcyZCPtcf4bFH+fMKbdUmfL
nKBgA1M3itwOFjk+j9KZjzhr/XLRhnuTtLo/UwwPnZEqSIs7fwuCdgR87XbBL4VIcWM9e/tZG2W6
RL/WbPcZe2YUfxnM+wnKjjOEd1GczTpFtrbt75v/rDAPUh8gt1Z6sDiOOd3es+xv60RjVhkvNL/b
VnUp+z/PoLz3ksKJ5MwM5Gj1bU7cBwSwsr2CrqxSwxC4uNkdkRgobduqZ+1hKUKBXLh9shJZGaLT
z0S3qqOOHHFkm+KroGCFQRMaDES6qRgMzMdt/WQ4mnZYuY8tV1t46ImnXSBywCwMbmWnbz6dzejy
fNkIQ+J3yTRMx3k4YOf54ciK8UrdBt6HdhcTadG+gcNai5Xi7fI3cvgMwy6gd5CZTMpI7NKTeK35
61lxNOt1vqQwKIfKVyFgGf/yaYnMx4hZ6chbQGHlpF75QtnQx8XnajgeafEcjmcqTEcetnCv1UNX
Ygb/NY4NGliTjKdGmOSwnqpx7TlBHs12FMXEb7nakdfRhv5TIJH3n+oamt1XAAppPPqQ12NqFMqH
BTWMZkwc96iriqvndIuc7DVRKHLMvp/goOZ570+iCaVMeG2SOJVydkM7m7xoaYuMdP9BxAhddBxp
4T13LYvirdsUf1m2fCQcFZDsVfmtTEiqYMtbQgOS5GX3/VwrqnZfgXOEy2QeZbzEuYRchL6EIdUE
K8RjLttJAWzCQepBBgowsRgXW7Hz2Scz6OK6rF1782ht4lSRwGgGayPBVVsYVd4WJSD6O94SMBbx
87wK9stemm8iUW6OeibSnPhbHUbfLnHO3k9/LTOSHH9H8k6HhK7SSKw6ElgbUP9As8kvehwLj5U9
z7eOx+vqLrGLVrznoyzqzzELsr0seRHnquJvZP9U/PuVQoXMysiJua8/PuTrmoQc1iyDnwUUzqLf
vQ7TqD7vZO+NKmVZ5WzjtnPmN3lcY8zah+UUeBJdsU/avm+Nrh0l8QBZpQrkgm6bxvaZaZaKV0yL
nWz1jRaqpSulIknzM/8Ra7cFxHltWLm0IRKw+Em+6fjUaTfNj9E8lePIyyOCBkDRYlreSoZDhv9P
HQQi9ej9buSAuPKPBNlzfn6cEA4EBq9XPB59VyF2Bnh5+aWeBgftnPjP+Ny4c3El8nc4k5fLRRYf
X6jOiemHar8zFEQ8clW1UCeTu7Bd4GgZuHCv7jlCU0n3Y8QwF/EZ/dzErzH9w9q5US2QaE+viWDA
PhFqRa+TOrMB+Fr7qMZkQWkvstFFW0QfVXB5BRNmfss5BqPp1LHb5Q0y8xeItOS+Kq9bGaS9loqX
Df/bO0d9DX5Y13p4QKZ+/9H4rvzBbttItFr3ODTM0hbikMWCiIIxiH2qPqKygHUBsZHpxZ2fJ01H
/XFaOpRG1Fnsxr6TRO+iOWyeGJ4LhXPJRpT9X2s6eWBgwe0dQsVlrEui3eLUipqem743BTmo945g
6Bq9OMBBH7ulxB7gWLOWWKQUKyuL8NJ4eaOlTpVAJMLSF1gBbe8/eYTtrE+qmwFR3AdMIIqV5jEX
8YlDZaNXHNEbO9DxRsJ/ovlLhtLtLODTOx8n7jbn6/YpGSKscYqAMZW9aUReJVNaq8ARDe56+vm3
iXIUnC82A3t8X0xBGv6xnP3I9+P6tbtCy9WctYUowa6PpwjnqAEg3IzF5RvjzDIlF6UUt4K4IDuB
aHB7cA4Nd1KkHXjGFZzmc8YXpsiGaWzuJ84Bk2MoM768tYwNIKzWhZDZ1RyWSHiuOztCmHmBXw6j
QX2cPrJfnkmEafPDCt537pjD0zpTX2vS8QJd4S1/AwOaYNKY8gGKTS06EHS32J/VUTuZsUZLYzpA
FiSljHf3aMfKjSGegI2L5X5T4w8qcL8vueuWxNHU32KQHEEvRM8gA+qqk16pjnZcU5ylakag8WoT
TsF5fQBaWMVTtooqEKHr12LMAkP/Y7Jc+hGLKstUjVmC9gyqDI+5iPrI9wrXT0W0EweVwhQZQbi3
rMpkpoWwvZSnM4CL4PtORpjXORRwwToYCbUiTDUK51Bt0zDwdxg3sqIbQ72hMgDFtNJ3c6OJEs9F
ci7IY+lIbgzuR7PXy0mznGFYr9bshUKrkZ5HVoJI4WDlVsGY5zl3F/MQMXVV6y6mcYiLv+Hq5YJa
DIFlELFLtnrG0kHIzjff4QIUdHu7ZW5mm7ZRKn0A87VSQOy6Afd/FAegZt/XmoZkD5CoZxn9YM44
M7WmnUqHlbcfzlk9YUWs8dZCzZ/o4yCrVjcKDhamiypJLr+oo08Cus8j4yqw/rwZvGMDx1/Xe/o4
h4qfscBAGic95MOdmoB4ztZVIzCfTAPUfUbldrccP4ofyundmlVS1o4/RqWvzsmv9AH2cRk/O2Kr
atZCxPxV8n8IE7ZGKgj2Ru3690dD8XGtZ5bRvoLsv/6C4FykUjqo6TZT7eR7b8StZr6JCszfRoPN
JtzE8nobHwPd4faec4cJMMipxRLRhO3HjqrksBPsmDeGXRy0N3OkmZXMVjT+KblYwYC+ecJkXoMj
d4uS0sY+R9tk9lgMZL/AF5/f/Q+l6+cpQEZtXq791ELpKkgP09tjoyEEaYWKeIVGgOJ9RLBAi+C3
IupXWJMqonimHvSAfNjLz5z3HI66dZFitsNBPRzs1HqgSQvI96gHirL6zShzaysfhX4q8MsexwY0
r4+jthkBmLvGRjrcXAXVwVdl6zvBF86TDpbAoLrGrdUkO68qcuOSvpLB0g5CPdJ5LIMRCQyS83K7
kWVKPXDFk7Tdi7wvE7MIXDFaz4kOdQIjiSaIq+bnkzrPsvWVOCZEiBeiZWxDA7iDYY7A+b4KnOXt
Mzmbvu5FdqdYXhbUh5VA0TnRHiQYbGYClvOih3bEbl7pHowZsxkuk5HGK/frshxb3ceipolcTiXI
KcESxF0ZaeznumNGeuqBaLbRniG7qe08I5DMWWU5Igji10qq9SkYAZFxmtQmDpyWg7vctFI/ZbAC
Qlg3P3UWxBNrTEBsylifaSrbA1YJtnZLLXsYVcA+mXMAcpP7wIdO/oJ5XFEtVwVoH3eIAyZ432fU
zdu32ZrV9GiNUN3AK2lRp9WRac7doOMhY3OC1N9j05GpObFi7oCHokoJEobTt/gfuU2wLCeVA5Bf
l31fzhyiQhbAifs/o4wvuj5V/uL7Lg7GP3Ux/H4iw+RkxVAxKwU7ogsV0ICbmvhtgx8ghj2GXGUy
yEy844ShmIbsn+heljZeBCFdQdFGuCAWo4ajOF37dCozP+HZTFyYgU0G9UQIs+pjbhQgcIzWVAF5
LkpM0JrJwkFAOxm8V5XRhdFCtsTQA1YF+vQ6devpcaxuGJaGRWTP7tJZBMDlwfBaqNBLmjKvrj0E
wCR0qSmqR/D1IL5QD0gETJrrOO0dg9sgl+nSpmnEuqVsji4Nw4dG5XFj62NgcKVaFRJojzucQH89
GW9INOaNatvQMeyJoIfRRAa/gXE2EpN1NkMJoyEurIeH411m6cyPST/xXzyWJRLVnf1AFM+uqYyW
jGY1ktNf7lzws6wrItTMmriYE/JCLe7z1kNTrv5Iy0G/HJHy+/4XtbYkO9lWjzdiZQSrL3dN6RP7
8wZtkEbna3gzuvg+Cvp77i6GLAczjk5QTa+VkB8KvaC9Xq/bRrl4IfZK81mLBqvaaIGHczEbUDro
C2VRy7HUyUGyJP5L8p5Z9j1cfwUzb7T2XMp2VMKKgKcbP+fpY9vJQMkJ2OE6cwOIxlNQIfJLg4y8
AC0k+54gUfN476QYBWvSNLD12rz+tIB36+0/aukhCsvkU66fEwUiOsimOzZeIh6VzUtM57eBLF8O
hN2ZJdlHss6Idvgo+DoUckhKDmxpXi1Go6UhIkGNwjvm7F10anDXqxP4BthqgnKHWZzKnkZbeATz
lltuZIe5P3pWs+Ri0HuGqLtv6wGoiTNiBE2IftsOBW1o6y1GHCYYaZdZu0Wtn0mA9q+E5DmNgmrC
hv09iU4cCHtgUrZikHS6r6jyVBIud498uw2drPidXZl2RTtwuKaokeQQqI1Dt6SBPpT8V0VYOO4f
DCr//+HVJl96XRt7UxnspUuKRvTpx3rKGklz7XgjGqcEVm7wTE0y6Z2sP02Mr99cM/Fy4foD0aCZ
4jJOn7W8wqwzXjYoi109hI5AymeRIQfn1LvZTy1hK3rcUNmV7v22HhgNaZdFjQJHHzk6kPpiCgoT
oBEzlFt88jmdeII+oOLCukaCHilrOUR0azwzIGNpl6ncOjrOoS7hhTB3nEw0lCt9nCyf/wQb9Jbo
lBIhj/qD0WtDjb4tkb2ALno7rkz9mDzgrqR1HmthkqEJbrVppL4fRXz2pcE6NxhHm3nQyA+1cHEW
YbwcnOVif6JYa7UaRMnY5NAOTqJmZFm3EFBfxH17OrB1NC9vPcyXkiNMI+mokZtdpZcWO1SJKtp/
nqLSG/vsSD6ITe+pUSktp5mkXoyRRg0BWlnI+AOxsAQV/VjSdREQJEmRMytxaVoskXCOuistFcQ5
YEvAi3EGe4xkn1POUu3qjS+pGk9CnoiLfCVk722PQ7a1dS5AeR+9Ij9fkoVzdYobqDCib13z5OH/
qspkbwr9H6oi60ulXGBqdHZmIEevVCIepknUIxsglJZKYUovI7387oH8/q+zdxi/Y2uONQOwkSTm
0XsGNWOpgFsmho/IjhaH6w3MYZaESL7/DbCZ/gS/DdKEhdo4XYcfMySu/hd67rVq9eArTQarQ9h3
sydgHQ9OfHTrdimPRt5coUGzBT5z4p+tBqKCDvYdcSnD0/HPYbOQVe/jkv8O4YkxDebFZKkl4xam
3Ax/lsg9AS1EAFKJtK7QsEQVJ8Jjcq2tP/q5+IFtdps8oyiN4FM3NJbEK5LUNBuLAl20PFrDm2EK
9SbCbIbhZQUudUnpHz7rkZr3dKZmSdJp9myGSLfn85o6vKycxuXz31OMDc+I4hTNczKm17yULEMK
0efS6g2obrrUvmI1VOviQIbXAq2VDc79SUX/6gBwL0UnUoMEdj99Umm3ROJm7L7l8N4CT3XDmFf7
Oekcn4WWSMiF81C89jCG3wFHo+LBc5A7TLSqR3fIf++FrgYMvYkbvHPbiHvZEMR7c3+EPZ7DI/J6
8X3iKtH5QTV/PRBp+6HKCdkK2PupgWJdoslvrp7addlqZCav6VjFR70PloAjQTfhacEB8JfqiYix
6BpUPRQ+ZacxTZ7dsS8mof+zFNaGlpnFbZkX2h1L00Dbmc6Pzmnju6+sFCJR7VZW6XdR4k1af1JV
U4Kvmtjf3PMU9KnK5RjIDwoCl1WmHC6mPLZiSL3GdMzEMrkVuj1W5BtxbNRzRLE3lGz5PpBO7R0l
62bab9DFCv/dTf8mNlRO/xt1SiF2JWMkbumZlPtNmwv7Y28VhDsjVvqufhOc7I5UxOyTjDup7L3X
B4dqq3tA9fBgyW2rM3dHfkTWPiB2ZgG3molRD38YeoQi3+3hJJgamvRu9ukt1o1omF7T3R9+Ghgp
MbFOBEWCURK66hinDyEVzk77y8NlbxTb0O0RfsvwaBvxbX2IHLCybrRA5jn3KeafbkIlM75EDEgM
NjFn3Gq2sUKSy5nrPS/JHpJs5GliBYvBkSA0mRFjUDM4+FMpwSLr+ug9ZznX6/tJlWqdwnK40WZN
lyQRUaD7i4WtXHEFRzjE5krzLiPLd1OzunBt4cxllMOmDLi9URcobRTvfLDoMncHTK77Sd4YF7kE
eJbbkUUpNFP8sf9ZQ5lRkuAY0+ScsQDj3aRXiWFYhKFRWFmB+b9zme9nIcClLhFrkxPs1JnVq2LJ
movQRy1XKgSWWr6oGIfhWiKg4rHeeokwO41EvhmTHByorGICfQnK6LAnT/La5jb0PapDP566zUzM
keCAEoMhfjpfUeUIWub32Ks5e42cBfarco8XhkYAQBRM/VVolmIP8Qb3T1aYsCKz7xDjtjJMajeR
DQ5hETHCcibeDrb60FMPnHphru3/+AwIoSViC1NojWsjAA4y+Gvrm/MhQA1+GwHzmwAGXtB+FQxb
BJfsZU35qiijToG0Rtz9L7MDv9RevZ62MvMTmfUjk85TeAt4PpNX3e1kkEHLu9++wDPOyA3Uy5x1
PTBUOJ3uDBbfUUqRolWU8FXmifsU9h/GZSP3aP/IvTD3M1jVmdsz7J92zMOIzgY0HPpW0ZsIMYCi
Doz0dRlRhI6KulFMvDr1+N2bZOP3y+gkebXrLM8pKrq1CtCgg5wkkJHPipJZOUpwTQL6JEb6Y4GR
xkM0xE/s2VCNp+y8pxHUqrsDoa+U6E40SIe0cH8Z1h1tCdL5dBk3V+tDrpKnMnj54OTHmWvcwNhl
Lh4FVXicfnpWW/dENKR4KjCgPmOeJAhuJ04GFqGatHpwwaNirVEUBY7fWW5Q9XHFVGlqvYbnxX4u
jqL3aJ9OHivnFCT1oA0mr9uzy42SLNmPrk8T8AKvNdXk79Td2f9lUH2mQrT0vlSnD3czUgP/kFO4
sI/jJm51LCSFqwwgGYQCvM7uAiAKnyxgPphsSXCg+xbDklghFBaTj8AREbxqlQQLYtd22RdQqW/Z
5OtmRjorRqzacq5gLPa62wC0Xs0EVUpiMrgbNwdSnpdtQpfK05HSbLwnFakecwUSsrwBOCX0y8m6
7cWMAS2AJfDSX9iElYOhqTdMPekXN9tihS/VleeXWPVQXD60vjV5wSMC3jypAEc6Hx1Jl2BVPulv
K+YsyMr4TpLHD9lbdK64HDn3b6ekMLmoO4ifU77O1IZmhKTkeB2zmTydx6hz9l64h0aWp4t/C2Ll
BiPeKhBcmRsqyFbvXwBvmgbjgHnkd8u+p8qJC/Tm0JalJ8Wf9gV/44fYYkpO4ITKbhd+ngzcE/6h
DCi67/wX7b03EPTS4/UOSY2b/SF3m07Hl5ODPnZmhPGYbo1N/D+swPZ1EnqX0aKOa5mJOZWgiUOi
sbXbKi/XwleAB3DxCpZd1aGbA16nE0EnZl7L3ssnafL0eQMTvwK5NNdDD23OFKn4uwBGyPm3qh07
Jqnzcbwx3ucnXkHofteOIJu0SG/etSSosaiJRL5+FYkfzxSCcichD5Bydr8dE8wIpPJr3agMiVkQ
VzEX9l3bEaGnyCFqQ5HSwPmpLDjSeAO4jRhheoaLAk2NR7gW7wXxh+3mNfeUqgZRlhpMpCwt5Nxk
0lFXpRhmsI9laq4PzF62T+EOGv5rg537NOB3wCtWUtP/tvyQn3lciubOV7KIcsgNjNx7QdhDCZSR
XMzgfL3HBg/YdTe8I7DtjSPpOoSmcSs0CUqdcVLXpOSWwMv31+FetBJ5g5qJ3VdIbvecuYG94tfC
O1xI0uodMSQscKR1KCny27Z0TT0linO7hEareQ5pgvRsBGl0PzAHEL5Rjk+lyxN3F790gCijkRpO
I2YAmMjL+SVUYu784hfjOxsq+tetib5/ba6JvppIqpXJLakYNtSqcCWPMU+TEPMXclIke/2GDGgz
zl1WzbHF3W2RJQvUQJNpdkim0BKwbXWwzcQhTb4QgtUg2jhK1DtGNEbYieaME2/5sLAZigpKvTLf
7EJrDqhTRgx1fol7UpmyuTVkYt/Ul6B68jmdQDpeX5WEM1BAMoB+VEYnyuFqErX/nrT17rXAPGlI
lcgeX7RUaUULkD8q0J+fiOcdoFtjhGrNvfKB6QfHTy31K9/WYh1nXG7r1hGQikyhxJZGKI5suxnA
KbgIRlIk0OAbSX4QlmK6WVwhDVd6NR+zxcuAqFiISGrew4tRilZM1EX8+ZeVd1VBVtO75M0qZGFE
2mmIaQA+3f5o4AengZw63vYB1PaaXmFYTVyS8tevlSXkGtbLUnGFmjE7/FghdGKGHjgRPx8yVD7l
qJ/xTGwovh6B21eZUWnqRr48iHmp4qyRxGgOJk0bbtDAwA2KK6nMf1Eq6zE4HdbXVGyhPAt5RTGw
duE0Zap8TknExpTKotwQKtMqj6ARPGZDYy6S6jEMqvRgnmnioVFAnNdMICB3W0FWQBTLINlvViKf
5bygmli2mnt/7rohUweb2vPiJCM+QbdjjPNuRkgCzZrm/ddjo75H9kSD1fM0JTtyHjl+yhFTSd2G
7dawRMI3RQ6/iyCsua9nSGSHPmWVLAf5HmCRLt/2+8/SCnosAK5QGWLtvdSLkw5/4sDaZR2npLHv
2hADK2DNXl9j3qNfA93rA9ZHJrU5JUtROUa8bCEXLk8A/Jea3zNsNKK0n8AMWon/KI8aXy0x/9/3
kBvyJ8Z5cke5b+sI8AzQgdOLBY6PuTbatLqjS29Kn7gPldVDMI6Jdnab1U53gt3qLULGIcNzcYoW
HPYvu4hq8g8BfhRRDILd+K/11Ql4ZT5rrVM5L0mgJ5cN2tZEZaC9aqpsG5nNunDufrdyIurHDgqW
fpVV+TzKXmJGHGcWE23uMnfA+ezpKs3cKhamWmX37AiXBTdMCs10foGYEkOwiDOTMrCSuaP1bqDy
kuGaUrLR2HmKlEf/bYErPZYGgo6uPlwq+98uJn/+KaD7mULWHIru+JPHrzKiv3JwuD09uXNe909T
gcRQsDSKkDVoxx8IZHkLqEz8KhaQW7quRcxo7DD/92C4nf66ecdvmHiSbiwgMKypJ2G3BTZrcCdN
un+8hs2e3ZCrgBD7/EILprUWDSsGyThHtctCbQy8s+T0OCzQvFxpHXyW2znSEAv4pWgA1+dSUxk5
d6VqM3pCMeguNdHrI9h+mS6HsyFFMijW1fulR5+9aQduZhzhnKVfuKaBQzj915dw/5GF/8I0aGqc
zYiZ9Ap7XyG7ari944T9sf+LcFb7IUGAOixT9lQ26VNRSdiPM5m8KMGHGGcoagJUb5OC0XgpGZll
Fs/LAxCjxUFBct9gpeW4ge5HZOAs7c6EG+P644K9F1yIcGJO5c9fbB+1VIVw0IFXAQMXLqC0k8HO
o1DQa1iwBNZZ7DoEx9tagSlhQlUijQoxIQ4fmnsEYK4bhPCJkOXh0WGc3S1Vo/kLRB6ZvSvZpKaU
+xRvQ6c2Pe7atYL623ygr4ns7rjPAShpNHeUnYcOS5uIQeOW0qPD23uey5hcqZn3QvDwsQZPtS2M
7EVtVKvHVOZjHuOv97i5IyGKAeo3DkvffH7Kldfu+8PVpQlvnd/afRUU5o/Je7mBkjXH5I+t0HUC
XTS6wjRaH3AhLiewEMG/vD0SeoX8KYp3V+SWCmQ5pss4b/tami47dCaEug6BCVaNbtHc+AWF7KI+
LJ6WTSErHTtHzZ0GpnuQKstxqstW8H8MiF7bq8Gg3ctqR3VxdQmEDGwkcirdxkj2+1Qi21oQNJU/
f1HFLw3HcIOlWp5pgVM5ldzWrS4E/ownWbs4BSzmoOqssjcXBqmMkqoWWKx+4ocsOjSQ9GZGDmiA
qxa0tx2RGSMVD2oOkdDRbFFym2iR5senteHorKeyi/+XvUdDMEkhh6z7tNiRQplsS4oYiHZMHjci
IjxjNDebBXrkPetQ7PLI7XxJCr2c5tHftpv1TSczwSPu4OVkrqyBFue35XwoEeZhz49PoWo4lJU4
nKS3j5gPCTpARo6t3AWBVYZgqUTsOgCyJuyTWKkJQ5i4m+L1WUqtBAQ7GU6yHSKVJErScETPH05F
ceNK5IIoz23eOhnJGDA3AGj1brrISBZ1egxfbOHMHOEQGvjEUA0fCaWWyqOWpukw+HlxBmSU/Fki
3336cLLeAJv/U4HVWD8KiZbI+tqQZQrpIm2n9A24mPP5jXMD1kzOxIVfBM1S/MrvrSUTbwIanKvm
As40O85j3yfC4wiTAuVADPUhVe6+HlJc2vZxrnrkQ/Zz/47ve2a5WiYYJHlpwXAbaYfCIHB/tobK
Ipu2O4XajaTEhncGJWGUSQl+ugHRzM928QgvI+ZOjUKG0ubl7FO2GWOqm7tmIXLlOKMjRKwAF7xZ
pFJx1gojhHXObyhB/KKkWaoQlj6xyDVAVC9PA7l9REdR3EqqeOqWrLyLvdOai+bz2krGsoUl1CQ7
RHbrpl2RsHduolgvC00mfYvWWge5vkEAmTM3XmLkLwWN3Gqa+/yGItis458p8GWpvJ1Nl64TibuM
PqMOtWt+QiXkfEn+9RmI8kAJWtcYDF03VEI6OHQiSezet63dXyjqJIc/BIhVpTdax73IfMW0Wy16
Wfy6CHdlbvPpa7yJ1Hum4iRe4KymfmNHq9KCS44S9NbkihtdMc/t7q1UpnI1YoRMI5GfcRUKBWUS
pzs+sw78dJI5wZ+SdJiR3h9FYvhgFUfJWvWfuUooZKmgUzf9FANzsEkabGywP3cXuFl3L2Fq6sgZ
cJRV8b/CT2+vq2r1IKEUpI8/hoQiITFC4Pp1l57lR2s4lKBRcIR7vTYzGdUtnNyvXCrSluXpTwX+
bbfzjx3u8hADYMfMdEhKpYe9B8KbERv+CM52qOrM4xzjor7AF4l+E5HH+uAWBpXRXS1bl5xkfkqd
OKf9rDuad1oU7J7WtfL/JWK0DV248fU9Ut6fmo32vXv4NThH3+L6RaABIo3sMDD2+INWY9F4L0Kn
drHsuCgo58Nav0RenKLbGb/7Q3aYR9+rkzl5yTSxs5QXwDKaIp2jP5LkXjwEWMV13jC2nQH9FVve
+0tGG2Te8+1YAcuip0Zmmy5eDVTqJNvlomtmAr83356/FYo5O2l58INOtZlqdT07r0y/q1jurDlI
m31b6zgsE8SFFMjkixHz+WHlAHE7z/pD92Df68bjgkZhLnrMHPQTVC5wVzOy/yXXyEtEl13esjez
TKI+67GgxJd41KDDmBWiBMz7PETEuo3QQy2CefXvu4ZVeaAQnEwqH0TGI4WwIy+ABDKn7db/tSEo
AmeLoEeQFitYJHr2w+TVk3uWtcpjZbdRHWqvIdEoIE9o4GAQMRtqPCaddkqEEd/54LY9Y4vEua7Z
50CaAuJ2fDb/fo5U5yp88gckmqmcSyrECUgob4ZaHmnjCE3iQYcmvfFgOd0gkweI+4mO7JkEGdQ8
6JWVCroSQFZxNePyS599rfJlXGUC9C3S8Fa26HiqglV74yfs/xi5fVwTmkBrENKy2N6b35DKBhtJ
let7SwUNNYQNQ3cqqxJ2y8r4q0A9kMqeRi6Z38b5hWK63kwd/5qFzOEfPk/ZjziWVIGc4FMgEs99
w9/Z++bbjiXi+DKPUTNk0kLWs6edNJcZMrO2y8JCeCJR1mXXVHlFP0/UbuIKdx5Os6t0p5ZfbqYm
A5GR3ISmtDlbkNZI7SJpvvWeG1WG1P9F6XsQ6uep+fK5smtNyR2dMZWPVtxIHowCiBKkt0gvGAJU
SYxjvH5sJIq+31imxhPO67CjaPRSjbPfpW96QZgnush1Dld+sOD0+7g4eocCpn2cBMKd4zWAmTAq
NVkTKJ/iFH/SSuLVP7Mjabyms2WpYyY6xowcJBpKVVShySmTWXQEfyESlG1NcJNJ3TlHfQn/mr9q
hoigKChco3R8FODocxkX8Lfwo2qJJMyIN5c7+jd7ydIQI/kw29hluteVd5Hezu8euqGDVlHF3nT/
ZBG+fUkCRM5X603niOLWs8TqXQsXsLiaMPPwXJQLj+HozmutTRwL8MSCy+uYjQ23Dt4/ArPTcjm4
Surz0rS3qp/iKeLZCPdq+A+1bfcOHHxoJSBruhF58SsuJRMO2l/xj/bn5zE1PJr4g7osEMmZ+dBB
DvOfR58RJTFby26LFepWXL3LLqvUsYXL7yrF19H78HSpFrFuka4AiNRn9vs55pvNSNFBLX+uurqb
AkmPhO+sf+tGA9X/G/Uvl/a5Et72zkJEiU2idnUtYpCuNpSlzVkdwxkfmX1VltQtJINZ7ywlaN/y
QSFI0YQ0oT5jPeCo23s8IfUVgdNYnyR6ny7pRcRo3nOgKz3UZpMlqAUt58Pz9TTx6wzd6Sn+rPzv
RD3Pk1/VH1ou7wypnVbyRbIsq9pcK0iNP9pSODY3OGRc4tWMma3gNAeBOhTTMiA3SWxbOR2ooA/z
01QFAF5l5BdGZ0YTHTSFVYULGdw67mg9r3WPIG2yJeM9aqGjk89ceVcQoh2kPdVR52nMj4wi9Uua
J8vL87tkOmv3djUuEERTfrcZdXQnElcDc5/Cs3QXk93NbmKYFBSF5ibOwP8BNklUcbBN3wMhhlu3
dFrxG/kss1FMBpL8kkaBakXZXjv8XlKDw2MTwO4ggkpZN+0AKKnbBALpXeM4PwLncAByMavRjBMB
4vIHEOVpp5PNLyoRVhbzdxzzv+0a0pVnZmQtj+km/6kXgeIeoT+j8CwLh1BktwNRq/qXBltFO74S
KHlmJ+DuXqJDF5vJGahYDc9JN6006MBIbPMGJaqdMad5cCpxRze2gh3L65UHBqf52CK3nVak8Hyi
6W+59w959aY+m78ht4d0v6F4V4Psr/kDB37xCH6DgNLcGb0ewbXiIKZjh3JsBt+tY+tD0mb/AyPv
Mlsy2YoA/0JHdHyHzqmJhiicsd4LIRCxEGCD3XGSKaMgRvRD4dYtcZjcNpGo33+LDqu8NjxRg+AO
4CPI6Jielpj4Ql73n4/RV4UNX/XXs8T79l4MXNBH1lIry7QaotZNZQOJQJvvtXfHAZQHDsfhis3P
6DifP4MRudCqfQhwovXW1rAWlT8EtreDL4+A/skbNkLJrWc8yU26K/U8B0u+ISNrI94wrBuCz5pH
yFs9Wn6NRsWa7BgvnZyG1VhoNyL15gc23Qc566n2trTOy6UA8RQYeXWF4EEkLUR5wp2n+tjNXiuO
3xxHjt3gTxAPlXfBTsl8l5bWE7A+buU+Uk+UabJWBHVo67rQOrvP3yZx/ymt6StYiimpY31Mes2D
gBa9nnT1Isz0WMwtZOVobe2QJnz+8fCQtTlKKr9M+nZfDoOghLojBIYRkUq1Ygswc8REzDScYXAN
FEVPz8c3FMYhS3BfqjtXPicN34Hcq6ArnCINO5/HWMw+P47JSpazLygLUb+Dna5kgFMA6ckAIy+b
NFmRoUhAkvmjMcnNPJr7I/ODr2hmHF6eTgZ3+LC2A9wwpMqwnsaCJafYFU0UCwa3cxTub3RoT+wJ
kDc6VWQinDNYeY7npR2AK2qhV2NQZVMZS7gjVCzPCWsibsEb9F/R84SXQRJHCOACQ3LHuqg1uhaC
jj57IiyEYZEsa3HCaxcjpDd+the+4044wo6JMnJbCjOi/HFTDYKfcy15ET7tmM2pbsbbh1ZV5n+X
G0kHELRzGswN+e4sGV9UaZLlKGGSjSDtksq7uea0ud3jhA6iOYR3uQw3AqMIg6hnqjV31xLv6RnV
pxAfNmjADo3M8jfIASsJDc6TgcLa7wPTJs1hAPqn/nkuL5uv3KZdijO+gekKcPA/e8wMerONIfay
IJxgIH9Llzxm7ZtrOYFIOO1Pins7w/X12VDQHdE7aU+LEPt4gVQe6IYO9gFx7/UjLFVXp/hFhD+m
8PuWXOA3NrmT0ZlniM8btg591JhtxzR9uGZv7ZJDpD2VBhbEclHa8LvvA+KwzuHkdUTz2n2JX7c/
/qWKnVKCIgvpwB4QX05skDpHiYUOyJ5nSS8v4cuY4+V0uxgfZ2WSjG4WD5+ou6C82MHTT+cEsZ3k
D5UtqxeE/xJlik+UT5iXDYjWNYgaQNVIlVvCkP4qCWuL/JAEuRZ7BIf2bO2hO/2TbcOfVTpTd/qS
H3nwU3IE4dhsukANjoWSXa2YoN2HREeiWGTuRmAlvwG9Ifdw8GHzqQAN4zUOAD3GXc1dX4tZbGSL
r1Ed9FLoD0b6/t7CUV5+KgNbZ8ymIL9dZlVXU9jPmK/f4kd0lOw+wTX9IYfZZ9KwP/nS2z1WIqKW
xmQLJmW613ZKkh4+SqDTm39qf1omVE5Nc6x0hVs/76JfowBTI0TZSEwFHtvso2/UgPM/OEgHEuW+
uCMG+O5pZ7SVJ6RCtRqBsliJebTcp2CUjtyev+b6aYBgpe2sZlwnRKqfHgiYVzKVWB4zu0eUENnh
wEo1HxI6Pa/byI8RpEkR12iFRtJ7raIR1gdmGbzYY1sWgjytepLRKhe49pCqsZcqRwOYJVI3nwbW
Np+y4m22UAsiAiPGO7QHBOZJp7aiA0BWSUTEYXlzBnhomJ0NEZ6Qkb8xItDIS/fo5OVh95rnJF6Q
7o4XMg8Vb/UXHAIDiE9bJTulTkc2C/szfvfttO4yjeQtJ7mL2mHdyZuyIm9x2bXynfG4rEGj4KuW
lvTisP4Ql34Gs4VGHjUD2mNOrwKHWWKYdOdjGi7/mEfO0k6AqHcWgyWG8ioXT7Q3M1Nm5NqmWz0e
eYvm2+Qn/9nOnzt+/HpSS/qUCwbNQ/47KnBr7ioyCeFUPcJBJi1eK+MbHk8hlkF62OMABvNR2hHO
BVrOJ/SM2OgzjPT1ytkYOENPWgmrdJzrK+4mvuzwR6v4AQwS3QRxigmVgnrcQoZSSP46/wC/N545
A4vIZQo7uD3T0G3CFk6oFkMG0utUl1vjHIuKvdVYr/6m8EyphNQxlPkStgS8dBNQoGo0nDU8RWBg
aOSTAV2N4IDb/Lv/Njh3+NYHnSUJshV1dL9t/OOFoVRsQ9UnEleKc05gs30oYlIAZCEH2iYcdM8m
3dz4ZukjflBclhAS6gidhyW1QCpz1/6EFWw8Re7Nv7vaJBE23QVfMJNPMoCXaCq1Vri5ucnrZqDo
pFyJeHcFkAGUQs495hdzgyICdmJWYzPMQbjtS7wJ7DD6smMmkSPPZ/2+yIwDkj4c9gUuYVW4DAVc
ZP+UzFhOR2kis+LaknvCjQUJsGpebsLM1tAqaqlclslqRGq28Rdi5odALo3bIDD/zEcxorl3t+cK
kLt/eUHDTyLYX3gr50JlkYIgVvX97rQaaQYpmCA+fMZsYhzsIAhdr/KOpeBBotJmMJUvzUY6MmK0
2wjiq341yyVtS9cbAQz3ANMxJvzJgSetKYqfdzxSlGSEWtLgX1yMOZbTRKrgEhCbZ1HxfDsb04by
KisnggdYooFbEIyy0AdrbxzdZdEaV1/7IO0iC/tYDlbsmUTf+hlb9B5MA9K5QMDU8ukSMSW8zQ//
kEfFLQnrYB1CzxdzToPV2kh89NM2qYFv2pB2/CseA/RSIFpvF9gZijIV+pG7ybjuh2o06tVmmVjR
oNVrg3DAkMxWIfbfsH9+Pd4W7oAkSecwZ+oG9c0HB0OAjOOHyOWx4SVokhwxD8PN9LOakpT1l3gU
6eUmJIDo1rNyqY176Ipa/AmbqPjy8DdL8avc6Cb/HPWNtbPeqlhT5siS2TPFkWbxu0l9IME5b4t4
FZgraV9JjeYSRG+J3KxiNlTlVSaiVw5ztJ9uhkGKb+P0lZPlsbUZhwWUhQzFIl/vtRPxufGwrpJu
hU+5JpEkWaoD8XTwm8QwkjnoYZ7GdDqw1wareZdkrRKVGKjbYPRlwRRB1NuYBgy0vnsAtP7tTI4r
RGagOXcw0w+GPQuhUWCeqSl+T0OPjx7PJk7lrlsFTs9sO736zxbHgIez9yvFvet0Np/iYWwgNrdK
UIizvUjnA4eCk328ijx9hR2pRUeZ1SayIbHVgEvMKR7bLrLSujOgd8WLQ3IfCBej6IuK2Tj7yxSf
CMX4+uM1S2sanz7b3OMd/qinxeFbl6gn1aWuz0/N1/qV6cfqcIDfl7QyD8nwfLJ7calpUYmLBhkk
JHv9MRrg1i/PCoOMJqavPRz4YFhu6FAe7Q2l9GiOEhE3lhNXjY/L1hGTedBnHEZ7mRHVZaObyFA0
0F8gZvHXDPxsVaTASYA8udEXQuJFQK8mteFiHlSCO2nNYUioLlpF19quxeBVmP4CARyy8FuMFu6m
nSvj8tOcT+ckETgaVAoKj0m7ISZd0Jgl7Hg8R+RhPOpw+XaA95CeGkvpsA//PzzvxCgn1N640Im6
QWsa6pf3F845EPqILIgT57vH/X0e6BjQKqIKYchD8ubJbCn9hyyaFBnKfpao4vejb7zMm0KdeP5F
AP8w1bXTq9nM54lg7xd7aA+R6QO2rbQcT190jeVe1d/dko5laf9W1xU9eUr9dtsnNV6/MwpkAsNZ
VDA3iQvQZNZ884Aq2UfjEXXZJ9+Dt1ZX3LExO02o0lNPz+K0z+3JxZ3RXVLTJgFpXSCkMlE1mUSS
Yf7qHXLXflh9hLTwMgzKcv/G5GSBhKLNBrJDi2Csy4p5XlPF3lYnv2lHADQ0J600XL8qXelNHPsC
aIqsc2lfSLq59W0eoMCMyxzfGvchrhywG8GW215oI0m1StDHacDcGnKw1OxUBUMN3uhSE9uBrtav
o7aNPUmOd1GPMGgbXyc/yb8YDfgczwzbmFeEIyf9R8IbE6NTIJe6QYVD8VEWYHhqf5HLMHC52dtU
BBh67pURfIFxlUKMdoiewCedjiE3vCiVtn3fHp+gmQxTXAkaRTU0JpBqkvyPy7IEJ+/YGKp+yBwg
98nWF05L05H41hW2hMBhgtU3pLycs+FY/8PFNx0JHrXc7HQtDN3QdIPPTD0lq9misGJ3HqbroBml
WAh2/cHP7EAs5CA1AtXj927KYw6OC7bFluklh746ZwSf7WsCOz9XbGjoajtYPe66jGD1yp4V0k99
KALeX1BltgHlXTVw6g8yBWCs/YxOSE94Mk9TLZtKBI8yJ+crp9GULV3SHvPeY/t8iWTKX4T07kX7
ujmMIejucJwEBBV5QLFr3p40w+iydkaC0RMKwMLHBf3OMRwEZvTsOSbxrzN3DuKAeZS4pXXrKUYw
hvsYsqqbdde/CdW9BtN1hqr7gTx4dM7Y+NRRhuFiducGwpuzaP1euulc+Kn9YIJXNVKQT6E0vxZ5
WPHmp6TFX/pj+MTZ0h2F0scXfja1jz9e2KLQVZcN+2jHbdleXY6eI9ArBeYuXTCTwZaG+o1hfqiZ
9uLLViwqHkNvU4slE6AYU4JUwT0kySfceCmRSfbvZtIz9mvwww7/je3xlqERsXt50fmvWT14aBs2
b76os6zO2pSSghX9KKDLGSgeUGO/UPTAhKMZn87XBfdIm5MkCntu23CS9Uh8jB+CYrJgSgBX6qQD
DjGUsUx3jzX9pRu4rzmLl7KjPpvXiUyftCctzrELSzhVu31F14KLEgqJlFZ5uvLA38UT3rFnIRXf
hZDT5FlmPOSgz0rSLOcKeZt+azEfTgEiifM2rWhcpPg/41JUig0M+oI8UqWt561HAeqKM3+1x10g
bm1uaZzaCDCaA9v1cLyef+JRNw+x3795i5KrBpGars4wBqJPiEddqoZC/m6HTxTaROWHr7Ajtjla
WnNtvRay9Flh4hWTYP2eBebDaRBfnurS8Q8vI6bTyZbCo2TvUvcH7uA1Bj28lo0/5aPKt1+8djG2
eV5FCH2X7ZTeORP/0QvaMZUzzlPSRj/xQR1MeRvYFnWcIUhmrud7nhBPUZjLLjZGpEb5hxaYXMVH
8bd/cVF/rxbUsq36G2EWC3gNzh5csxyy9YOS/fFqLhxdKee3E6wS7MvAeqJRudkzEXq7mWcaIPck
mRCXi2IRqK090aHA4NqRyVKVeTMDLUaQXHLHAVEZKGFHgveQic4lNRVwXCt/3xnKZ1CzvrEGuP5k
YWJ7sHjKfTpAZY5fMukFabpdkL+0+4aJcsFuzBRr6R3+M8qYDhH/8qa+7/wyP1H2U512fHz8BImi
bt93y7qSZ9pqvEYf6B96S9dzjxYdjpOCdR9kiwxW5nNriRTPcCSDqJpkAvmo5IdBrMykfYhlzAKK
DRcmuj+MuOihgD1Zg3mOkrPtcouXB+ztCyiHGR4ww2c18iuaKxfYOjJL8na9JsY1IWGHyNXg6IQD
FAbRn+Xk6eh/fMMf3HEbowJdp0/OIANFXT91+MkPxjfvqp0w6w4ucUgRgA1m0Z13wmU0wb8veXw9
Q6c0JAZLVbekqUJxxu90zUAo8sRdo7H/WKtTNnqpxWmjDDSJq6NCMrfrCnmFC+b0yErZaW7CDKvC
/nyGux6hVWd6HMtGsMkW3Efrz0eXE2YsJhUDF4mhGHfPf66+bxgdt9gJdpzoVfpznr9EvXrbXnK0
/Ay/QkzllyMs4ffLXUX3+2m59pUcL/mOM0uwIdTLF2ivrhSUuWIsxC5jbItGOhSmr4dG4sXGNpOE
99cXb5uNrblzuxP92Qiubs590VQLBoHyLvJeT7G/6q11tSzRA8GTDefxymgZ0ddS2j1SGUPpVv2G
Av/KcbrRkKOSda1WqsF3mra/JFAJYjJhI0RCVJuqqmiw3esjIgfq20nL+os8HIZK7wk2XyXJjSgc
Sw320tV4bMSnWP7S4oGxvUu6+oV83uJKnFvG+nqwN0AaRBBku7DSmUkzBmAJ2Y3Po0jH//uI8jcf
z0hFOg+0bU9uUjLsnW3raNEY1+kmOq949DZ8FBeg5aQlr0lQjgXYxh4zEGLSg5yF69FzZF0fwQAZ
LthbX2Csf0qG+xgcIzO9AISKj6VLRn/ucc3zWlyO8kTM4hLd8E1gAO8PJw54k8PAiuO0wkICUvXi
xL2sGMw0V1ekm3O3rx3OQmX0BuIWi6UdJOnvrT7UZQKcPQ4Zf0WE4+pU+4gQDsW1g/TA7ApeUL+t
k18/EkXAP80/NWa6bxokBSiXAA9iGUX1YUZqYWH1HRrKf7pZZ/twnvKdu07WwMrB714am0SX9Ik7
BiBoUnEsQMuuckIfld9MnK7E8jWxvzFiDJZo5XSuiAvJi2yv/c4mqEEfz0sk8DkMS6ZQCTlnCHwq
4jHHnx1L5JJvv3KVW6p5H4AmFMd5diiJEFMysQvyjBE84vl3e5iV37fbuXX/VMFlDRFe6Len0QUp
umxhDBprvnBr/bS4ALgqVBpu7ibn/6eVqwP66svXt2dCVZeV8YY6bUEqD3L64ATlIkmMRVgx3yHB
LeBoXcDG2s/sil/jue7Kkky0q7g5i7wAzGYWLdRIs3sOTCdaM4EYvAP2GcbgWz46OAfjrbrKX6AB
o72voJEqtAS7wKCn8op7xtXTj9o8ENfjYB4rP9yqeTq5h6ehZCFxivN9nh5iPkTfIKW34CeBWlXM
RP6Zp49DblBdZ6W40uKCfuVhO4YfGc8I2Rs7EQiAvbT6oDcImRfKANXDyZy53dJc+PT30IGyIXSq
kjiznta8h/gmQc7Kn7eMXeoD4iUEUpJsrP9lHjshOisEvAlFXS82XbD99zXidnpv3vvAehuaqzqE
afyCBcc74Jip4rm/XdylgUVRHN9KrJCgnP3zP1Pti38PbktNYfhUsDg17cvFmtNUKKRp17jeHNdF
jrtc28nUx0BTQbViejUonTxoSeWpp8LyPcUYHjuVlAYapSsNqNL2ybtnVW9k+wl+j2fdBKm6otdr
n12nCkhfaFdkZXZSnp3/BqEsjSJ6G9JFcBpSeZ9CIYrKjHL3DgDQ+kfaCqNENX+hgO71okaPMmPo
1VRm++lXZ1EHktK+H3pd3aL+NcouZTVl85gmlMrmQ4uOs0N+Bs/dAEJnIktz6IPyC70VnYEqhOOo
eb6GRLnrtvKeC5B5eWc6P41pAeyg8iMreMX9RYPJMdk0rsYkr8y/JUeaQTcVQEW4QnARKTkrnr/4
Ey015om2tpj+Xvgsd9LCCr4wdrtPDbTzReuG9/NdYH3NypcjTXVis7eKIFW/KLXikbVx8muYhcOs
hUFp2tkypN05u72aO76k0/eZH4/IHfWoK2nTaMWdZetwPPXmmBqIxSjYYXzD7EdhFzMxVdr92/AW
XF0zyiIfse0RagK2tE9xJOh5VqwvbUF25ItysTAa5RDJiRkkTCXEgtL2ryhov2qpRE2MdgD6XW+s
aLpDziZu/LCGdABArC3pAE9ZzBlvQnYNKSfK1iClSBlck0/PcZIB86SPEzeT6S25z8dF6RtN5rWM
YVJT3tbwCgNuRpSD+rXUnsya8142Drlkso2BU0tVZ877sYi079rrsDcWd5lPAVZ1EAEie5bMJMKr
H10XX3rsLzVuPGDnsXpjcglvSdWcqxh2v3PTJ9iuPPYQ1SH8CgfF+VMTG2dHlHMEuw2Uq4E7V4zN
scZaWaBIBghdcjvXEHPm+MCBxAllYT6s1W4lhSYvCs8/ow49UjIed208h6p/la/Dzyfuh8S/jWSj
AkinOfwL3bQ07SyrbKMt6aeNHswlrfS6wt5zm8IWJNfhDvpHx4iUqqFHBH8DX9Q5oLxlLrkMwAfy
6pEDDedMmMO6JulpAYoe7kiCDwfszHSCb/RhGsnT5I5ZTxrr28Mf5BmqavvtDOgkmHhVst+ZoSkX
3j6o1YWVgfjkkCOuTDBjMUC9eYRE6K8UcU+Z/yyRBj88taSo66EQeszxz39ZIas5FmAQjPLoV77J
GpwHeov/nFlLD+LHwXlPGwIZfqmeXayt3BtGs9v22xBGagJ/4vN3xaqwNdb/wzKJRA1kK1nxuZpC
jUchk0QA5LHeF37B+0JwXoJBvrG+RRACLSKk4EKNy1kaC+asQbkdELXt01cYZnfbytdSuTl9csUV
bZoJ+6Ph1FOkxbsOtT8diNFFns2tw6dYWjMorfJHivWZ4Rb5iguoMdD9WDvtg/Pge0KIFkde9n+O
9OOOixctZ3xiJu9muR5GQBopZLurzx1cha3oB2qXKToYi2P+/A/KsoW480YxQsOBczXhtDsaa4IE
sUlEJB+aNOK1dHU1czWh0xkd92KRC8jy6bxz1Alh1dh6zgxz7Fn4D99YhX7XFyBGBFvJDu55LGfJ
iNI6MWCwilh2R1nz8tJ5mu5B9OuD26HQxV16gEc8a9JVuMobspg2JczJWtxn5lbZOaTQ9hVCn2XY
ELqx77x7WS6CbUwuDcpZn4RmHlzmq9bES+yG5GmUxAOEjqOIUviMfJbfJAEWZ8OWbjBg1PR3MtZ4
I44egwMs5ONataQomCYO7oZV7PHr9ISUVM71vvQdIJxNYOxbe3Lz3HMfup7MwvSDwAaBFSMDtxLF
Ge7XIMezgYselDVVKnnhUW64GkPeFG2qFm83zJBfY9IWw5tC0Cq8+y5jDZJFdGrlsUX+pQiKxxPQ
iJOlYmwh9RcIpyZR5PdzRjLRTQRRvECcOWrVuWLHuP3+k4qwWPR1LeqrU0Z6MKFiemJqytzwNFLJ
CGDsVczfarbWD6gOx2J2pa5Ic5iR8L07DPyauZfMFjc0pS+OiMksWd+jn4i3IYdDUsFbJ+4inF7u
610Eg0PCoaYxjEp6SuevcBiCVbpkK2qZcYPbMIiHbNbnVsZdTEWbe/bfMmtKcoqMUlf4ZiVDzqO0
LraoAnTd+IQBGtAbvUnyyKODHwuWVwwfpKO85hUgtQxJJ/61pf/RISDBC+bh1geMB2oZkpwcMr7W
MqR0AF++TKjZ28BVtFq2LmUKEmOb3/fIBoKMZ+JEeQxzRGcNRdtHhTXyrmKWXt8o6aV8h2Hp3x68
xBOK53oLk16A8NnotFda4uQMIkBqPbFjH51fj08Vkg9/2+sLVV+3QnPjxawoJ5KZhkGibyoBPubc
uC43J14Epb3MBtbypI/Q9XkmT791t4ruQyz6s3S+Bh4KBg8p8jgIOuQl8NN6GGvmRSwvBrNM8d2L
EW02fr1HBkdSq7ztspfi1nyf/e1wbvoCXuZbqqMZSovIoS/fKGahWDIzurePdFMPsxQklSILdI7E
aRdmd9oW5YfMR/jsTmHoNSfHHMkJ4SvM3Y+nxxl9U5lBZUPOciprsU8al2mQ0P+cn6bgDX3ivPpx
IkVKFkwco+gIDvB24GOePfr0hFJcgpyi8+K62pMv0tELyiAIXxzGd2BIXTmBmNsGJJOLPLpIYPdN
/BRMXuCur7a1rkcz7z2ooVY7iwfyreMTybwD4pBftXIH9vAfLU4pEz3YH2+uYGKCCnmjqI1zkdVa
vbHUKITRTfvVQnUHRusBnnuDU+3E1q0TBehZgIMxdHPf7ZNGWuxMcA8zonCIy8gd/V5CWH+PFYbS
Sd+Wj8TxEfym8nYDioIWOAj76sgiO9mGTeToHS9X8HeCPMf5MnNMWz1//YTGcU1q3OZLrUAAzjlV
lBJW/FdXnX1sJnvyFZCfknvsC3pm+sqJlJuXhSK3swZcAJKaxzokdzzU4qQLMhyJmy7I3Jo1ac/9
aJrfR1ANeJBy5D59jFD7N+0/0YKr92pkuXKbTGXrF7EtloPb0AuvvDdak7IsmwaE+Z4cBdrfPb9e
0D3R5JFtNZjTupk/RiEBYe59HcFUnVHhQgOxmicdU//SS7viTBZKtl5JP5a3RiQsIbSSLdlj3D86
3AzY9ZwtkiFXDOdPVsnLCD8b4hKVTU2164P+fIf+eA2VMQsWgChYAcV/MMaah62Tx1/eBP2Gf3SF
bRBDS6XFeNMfVeMw9Si732l8WJvl59jMLMJQfGjoo2kURjjookRgWlG8M35caE4ChkeztOmzax1Z
jHEorAhge1Ctq9dkVEIUDbZ/3U+qv2JEHkM7IJWSLtsbhwhLfkPPoJrlJotjGis/DyDLcrJC/uhb
mBdQjbLO8w/Bnq3FYCC/+Iu+bm2YYMyoxa7S6k1SGOWAgy+eES6FR85Kz138V2uApRjcaPGvSm9j
pT4R2i686EzK55si5feKmZvxchau3th8Q9t6rew6UAtqKMeYX1ePogX23IQdpxGTj/1LMBLwZjn3
YKKib1ZcJ+QfQUqz5YdoDgsrgfm7/dJow1brbKyqPvsSU7tjEPiHQW5cM+VykIWzYAKrwJQqA/Sw
4H9F9iF3RKMsWQwmaKpR1OmTJl4SOqEwh+4EXIEtk209H2ULV9RKajF/ddzhwehGimSB10o8JS2V
bqsJOUB0zNQCOsNdttDegEy1pxUXrViCjgi5fG87xBI9rmeRGPen73h/EDFpbkmfeu+nmtf3BEdk
g976V1AgVWgkQgArIHC6YWs+g+YtsyIkylrxfLKFOKEij7vqHCYWxENl+MXB3plXgTF205YsenQm
7+fbQQ6XnKzlyig8t5/xt8tMIYljzUhI4p7exfDqThWwE2LXI0M+592d6cVZF9AcLQ1rl1DQniqG
ls5nxLH1O+vLeHh1+tmFoclOPaKD8ouGzm2iyXSZLvFdQOZvOBTRkPcC6ReYEfB3d+iiB1xoUAU4
XoE2jY2Zdw6WGR8cFtVcpQtMIE76t+rmuvOoJGijwjc3lPlKDHGPHPKUTvS33YvcV4pF1FlqLD6K
zVOgksX+MK0ehEzucdxzbP4//F8v9EOJ/KP1NtsHIqF+z3ZoH5ytQLJnYlE8S6xzDxFunqWrXlMl
K8n1CPysVsoNfyNDO2A4KwDmDtED/Jt4JY5+USTiFfFq45JJtsoLtUz8AJqpxFQV238gA3v9YNCu
6EXhd53U17hENd8McZHsEf6YMT7snh5RYIH0GskZpDg+2njf4GsYJ34zThiDCpzeA8/zPzgCsYXM
2ogs/jjPIRJiJ2/XSaZPl30qnAcwgW3GfcTgUcQqu/cEpoQyjyUm1RhTPceU0d17mU1eQwv8qz6t
ak/UbI/kNWKpjkWt66B+s8akA+oD3Yr6aOEBMo9lpZePRwVkRUsQnAg+Vlmw8Yiu4ebBntWj/4ZY
ghkUKAduNT2+hIy9dx1Jg87ahdmLOUN/yKOIPdn9fYJv+BBdNWDYd0v0bwyMoaYcrG+jiviTDgLT
mK6ASs7f06NV6JcnGaituGARojYMtTsWnFyxSuv5Ln11gBAxy+i4UThKddQsCss2FHjnSJcqM2SF
cQrlksqte7cxc5/6KEjUkhKqwNTR4rTGuKAEAkWms8H7rSpD9N5dABqNadgQvL6YSoNqH/Ik8Bm+
ObtT5GdlwIduvL0SIlU4hk482Kh36gwdbl978LgzqxMsh6i9Icr7abPR+lpLNfdaEzoBJ5uZ0fYX
uQkfEfwNtc1vI/BwFxmdEbecelLCMYTRiYJEP7GbNyk2/jzJeHl1k5w9oqwFlCFHe/FIzMrRO5dk
ft5Md206FZfydP9aPQqAQla3pFHlxYsQJM/8Xa0ic1IVRshs2IJxfhkM7OlB7VwGvjXmluzb5pHY
mKLbeTnECwbic/eVbY5GdPbQxcaeOK/5lwxod1t42pcATP9kyFdHnIMU4VXGh0zyYqOVdhMTKT32
6dqDADAMK7MmDt5ZF2ZkmEUAxMy0hesMlRR8nmF2wnTwf04E3FeLYH5oJLZigB8oVcth3geJTKzt
E7/3H/54QLipsPaXRgW9zzgVBCifrhXoT90+2wO6eM7PSpbtl0XkX8UudT7nk28XH3rc6haKnv2y
yzzhcr9AKPaJcX2nMvMVF/q/fu0KWPVBIiBUv32rNwR+YUn0ZXOWB8AGwo0jyuqttbPY9rt8+8lB
WdscJ+JSDtmlaP8nZVRWrTRX9cecPfGERdkpzYQpVZCKCZ4e5MMFqqwhRWAcjcim4HyXQqEe8ICc
xrVqa+QPQ9ZQxuwLv9yzYgjvp3qX0QxIGNC/FIwot7wj0lUteh+tr/Ujuv572HqnE+vS7ECJwLPf
BKquefxQPfHuLDPhUWhwqfl2qClAyiuCcceyVU2FtE7Q7gXcJbKt5bQjr1D6hdsazdv5Ym0zmYr0
ny8OOGDd7YfLnPvJVBu43SBdz03p5Xqrar2Bm2gC0WzpBmX6zyz/eVgLpIbjSYHsoknJywQmX4GK
6Bn0g3f1Jk9E1KRsOXCUQ80Vm/UNVcIGKEVQ72PZGcIssp8tXVOW90cySRvmzn/wcxnniddznZ+c
M+uOJr9DI01XdamA/iwklGaDOW0YUygzIS647GnykxB9BOpnZHs8I8FzLFehalRVKJ1cS/in0RTg
4TnP4hNZBXQn90GUrOsbhf9Axyq8w+uLEnrRhjxyoDGlHVrB0ObCVP7EUzx+t81Gm6y0JMuIcOyu
1jVAccXHGHgPdQghXifc8wxH0cGuyWmuxIkEvQE2LJKkJehC6IL/gFqSvawLH/jxnFBz8B9yeuqf
MxcXv96ry0XmQwmZ5aouGKNEDKgQFVBheidibgEkP9GB+i5xVflsYlyDAVU1x0q2fOnPp6fpI/uE
63V+sHM6L2ihw6KcxhTw0NXYWaHxtCUdjxwRNJ6mue4kAfPxFRHcCVHFWyHyEbc1CBKnigNWz5JS
bYVKDWVskq/4ICRJmxMvfUd18HjURT8jJM32lBbsLLIGMnnroebTP+IT5/5vNLaQkXGbKgcKAMre
aDnXVYoGzt+8+aOJLZ9WXIYJCf15Bruw8R6bmUnyU2+elJcfS0lnBbk6DJ6YPXfdIxF0Zvt6HZWZ
bfwNYlxqN4Yk81/xdgOPMxlaeNaz0yuNu8G8z8LrInGPSoQF9xr/YkYrm4WYTC6FJX77HT5LBFTu
0qO+fep95D4biheMk3rJBAWLAClpkf7jdqvSBvNroRrOOd81zHZsl2Re0XcSoX0iCCUiyvQJVY7f
hOKOfGVhmGQaOwG4hkz/+gN7CBUBXCegreVxAc84PRBCRTKcNb9H8rKVv+9Ly03u7pJWQwMaxbA0
MgXw/2H+sbuuj/QNkW97BHSQnCckAlH41PV4VXXsg1h+wEKNAwuJAvnnvz68T/4vcUEi8VuAOO0G
WHhRRh2rVomYmlbNMMfqn/5Eox/29FeXviebWvccygwt/VVUCLF86MldBAR2kCjq2O+orOOTat8a
m0xV5386TP+QNmcti6v0XIhA5LUEQygBW0y1632/GlhrtZ8D+8gQvD104t+w+2Y444dFscd3stTR
Tvqlem784lDwt+HcaQst/IMaUpKuRxr9rQ1SEaTSZHSTIIMGFxQqkD3lqJ1IpEO1BSFaqSET0Ups
ZzLOiIrXe0vQwbGs0bcL3MFWe9O/C0t2PKFxnhVgnk6kaIrPtTfEkjI0RoHsBik872DtsWQQlzYe
aPgy+miuc4eczKMX9jA1RCjp7LGcG9bSJ1JK2J0Wj5roielkumnLXo+fbLq/LSlFvLl/dW9VxKBg
nt6xnuqh75siuTWzdJRF7Ia5wUfBhpoAZmcHnuw8iLbEMCGEypuAuHLsum+D2g0+LiP6PdhMdSjV
Gc1sNxSTv2e4EHwqsHuBcjKoZhoVeOZwUZDIc2BrJS/i+P3gx0l3ae3EOEgFDWzC3wJ6CodCTKtF
Hn1aCnl2++sQS7D0ZSLmnYVFpivVk1RnhTRyZ0m5zlT55lXpNivYVtwUniqYGqMTfVJsG8AZEXpy
fRJ89vpevU26B9CX5K8Bfy6H2MCv1xAW8uN1X+tSNTZpXdURQuUssADifI7vdvGS7rfmEKqkVFeV
OLcRwglNcTk68QiQdY14B7Bu6JC46vCubOogYWkh81oL406aQ/UHMyRjFzkh2AOP8iMLOqjqvdbM
k26/OZwXFLnZaFCBvuYr421bz3vU3D4TJQ2A2MeibW9yw4jI7aKP4hR7y8bCVdElIr57NmQDs1+z
ENN1gNolaOrY8T70Uhg5wvZ5bO6pIFVdigHc1Qdcqp4TAtuUoJ6r+1v1mvR8ZZv/VRxmXJ3HnGyF
MuBSlmV97BELds5UFVav7v9kmrWTAoGBGz7mLr+gGDjgeJ/GvZsHNGvUbojVz9fU4zn6UOfu5RmO
xteaYabOITnmnuXBfBcP3UlHSrtBsIXFIgBCoGnAxRFWHDPDjoP0JbyRzXtgO2fn9a5kQ1s2IbyC
H2A5PJyPxFIAZtHJbJ2pq9hoOMYb8zjZPPIxxoob5ThQMjc07zJuynF7Xg7mdUFT6WOF6lnsMk+u
itTfxYp6jEOA4xhvfBEw7lQ5v7lyd5UU6+BcNuxfowgCtu/Xvyaw3r8wks26+Kd7THb3xtFpRamH
6wjpSojvGdWgS18M339QNST7NoEerrORW7MfZr/XxMr/svCrLhw1BilKcudFB3VHuDs4dytUVG8k
pUbOAFwO1w9eU8yF3lidHT4rsEn8wWwnvdOnCsnskOT6W6Aj/OMVxlyMsyAkkYR3o7LT5SxiWwAR
+zWBdKFyQt3cR2+gLNnJN8I9UJgXehSp+7FGbht8TljvXYFo7QhVJqDhAMUerOYVW4OkdHxWQRHs
YxI5V8rcowZJwSO6JMZzSWWzobNnyxFja5TtFQtsQZDEOtsBGPwlSuZRqIrFBSBCuW4RNGR7gOa4
+VZAFwBfrBcVClCoojSAdGdIPHU3UzPtmQm8cgeXgS60KQzMsml9XZzhrJJr5klqTLXhZr3PQl8y
UqNmsgE30pzeT7tiAlravNMDuLllBupA3W8MOVHQTyNumgRewPblQ0/7TQk3yuPOREuckKrZO/kG
FOfeIIBL63U4urOmReh0WfLyT9HJblTlRzCaz6/IKsRTzZOxWi2OJs8ShiWuhxYqQWM9JPYFnZ+l
H4RGDMEAXA+j3e8uBoZWTuL1ImIWQK01AV/Uwcs9Q13EaOeJXzoIfsOrPM/phtwI0zq0YbhBy7wP
a2gRsWEbSb1KBhOZycF0ZsHb8BljE6pqic0R8wsMungERzBquHbtpzR+pH7QscuIXr1PHIcYzpCW
8Gw3UeXQJmxH4QnNhkzTMuFup8ztmlQkUc/n1VLrV6HYjEIi4kMIEePJSGXCxvviZ53p8fzLlUhQ
7Kz0TWl+dSTmNNi6/STWRI7+afmeqOhbJi4x9kHSFdBez+M8pOHCM66CKCcbj2qwhgMC9qMsO4Bt
Kzxf9mj4Yf3zcSVdBNec9bOKK3Fjbj/Lxztwb7vHvIrZGMZF9wUySgIRaf0GNCa94Bqghl4/k4QZ
VypxBbijcWNbgLitCnVpzFur5+y89GNJI0xSQocxXND7zou7zIHA2b24ZOfes5lIk5nEKwjitwa9
jymuyyqjJCXOEMxJIbxOpJxrOquN4yDzUGk2wAVlZdx9dq0eaGAc93ImC1916LahRq6H5vb4gRHs
OaDglFYosMoCw1ZQ5SiPoDFY8kRXuQcHixnuHf5sgUs+PLuyJ/gWi0BatkL7GcGPqW71dBxKwbnE
iH1HesbCluXDLwYe59DJfF3F0WDB76JO8xFuAkbPDc9offKzzFIrxkLajbzDsxM6sL46yY/vrtqi
QyqrtcgBzVBFCq1SatJ1+dKY1fU+Sx1+2R1bE3TZXNzWuma/5ehxbV0fCfYNjtI0k4VI1cNqpXzZ
RuPfchTX988atjDY0U2v10AWW+iLtCGhgdkilQCjeXMYrhN+RG7H7RHJgxGKXYKQnK3mw49alpJc
HSAKBhdCUi+lejx8LrMfyOfEtA6vsPbIvtNPyKMkFzhtfr0sQQ+wqC0fHrZjDmDhEblZLDiCmgYV
3l+MGqO36/Fuzb7e67QW4BUvOUoylHQwJxuAGw+Glx78KshybcotaXspjeXvwqf0QaYaNeZlS+Mo
RsKLiNYZu9RGU1XmgiXwpRbrdanNqQz3YgBpgnaDVUlLptdHJOkcaPFnobv4Cy95jRJd/pY3B5Ub
swAtOzX01iDyO8BPsenm5LSowP71B1suEOZCEvzAqz/BSrTFLuH49LJGnfntqImlcNmkdCVLtP8C
xIATmPYvTtWvJcQG8hOMbJ4w6011CyrwXWJHX9vmvU++zVm6NOSQzOOfCIgjLU6yoerd9vh4bG9d
Rl+MPmpE2B55heshgI46UAVP2kVgKG+2n9k3RCIhrYAqiEpfK/pKRFPdWQZLn+YN7Obgpi69TsO0
5gpY2uipXrjWNqvXp0KY+S67dgPwmxH9cQgsSUsk1w2Bn09PIz/M579chLzN+x8WxLrV1jdXK9Ry
XfHnL3s5Amjd1iOWM5Yb3+IrAdI+tQbkPMJCxBaD14zsPiH+/QyJRTCc5WQlQL4ZX6MmYpTAqLD0
6w9ttRdeqZTLZQp/jXJpVkjUzLBVDne/c+uKigq8kGpGFXDObfQarqmv1R2ufMxT6eH862mchKVw
Fo4a+7B8rdswrGlU8vKXEmlxmNu4h5aWqN13QXQ+D6l1M14nZ/8/Y9mdsBT3xiO7y2MVw53pzbCn
bgb/h78Knx0KtY1iEkY692094uEGO+JbDN9zIOsxjpUa7ymHhW9be+UwqQnLhY2yGUtd8YAQX46w
GTNgyp6KMoDS2eV8if3lB56dYsKNIIXl9nU2unqTtgnIeAuKDwzCjpnQpwOzwzi28qpDQ+AOyPRm
XlSUv+CLL0nYd7sY6vc8Fwkmicb8UcQtKqWXn2+aRuDyJRRscwLLoQFGg0QzVvZkdxhOwl9Q2RCT
pcc9Xx6BzvAZYNxeM0WGnMYXyhg5F9B+lP9WSpFt0XBK50veBPWgWwgaKd1h1GB7nFNYM5pktzNW
DlRXuQu5qr0W8iwDanG6VG86UFTuu3dSfYAMmiDvYivVbGgpztPcqq+U6tE2JZDpSud9Qlha88Bn
EEyEOt+KBRgVXvlzKnb7GHl7pZytq8IQqW8ExUDvNZLl7EfYGNN7GZSDLEguTNBh/OJrvFf2LFwc
mBk66Ltk4DpXhTy1vTAhVUXXY4H5Ik6Z37PCtjAz7ZBOHy5TaOcO9Zz4gCgNRxcaJzrjKp8ukBmf
55viicFUkYKC0UUYaPznn2jD4dUqVFCV3rVfk+16vNtwqkNK86lfek53Ow3j0u1AYxUd6cGTQKAb
p6wCH4e0SwVrUcQh80mbODrAPdi/PnG+t3bXDP05vdBbOapbEkCXoCTAP4LCPbQrSe0ypxQIVhSq
1yedd9N5Qem3hJdswRdOXUh6RDLhsHqhNKbbhePx3N/nNzwt+IV7NIJMKuk13xth5axGOXdDezye
nbSPZPiYjVAdWKQ29gku5uBv+ykbEH0TVQRCtk3tu/sfm/7SeBOEsMB6LUUkAmeCJYK8nqr5Sjdq
UJmdiOFA+CWdxIA3iL//Dlk6YD5QaKyP6tKuOvIIFTELkiqnXNYztQ9nxPfHau6+93jNQ8uEP3Ol
F5se+EMidzoXYWenOgLQD8rr3PvhGRU+zfNziYVQ5ImGON9cfS20I2j5X6DFF2PhVPxmlyEWs3ml
SezjC7x/9isRU59n2ko3UL+aXWi4eMAXI2cdERrUzmOstRXcgOxHBSt5fdvT+GrdmkQI7fZC5aUy
vTJBDwnDsue+DZEjUkU49inUvL5gSVbM/sI4H5DXiNLzSGMo+xK1QixTkn05iqDM0rbOGOhuGOle
eOtIRSvDbArtcTovLBYrMPgLi3GyhBntCBoRUNp79x+V6p76eIEVO/Kep7gGF72oTcG1hqIYN7o1
GHjYHOIps4V7TQh6C3sXZA16Eo1GpnRw09NItcQVwqYT+XO4T5adZSpRyZQ9CFZZpM0AVE0fkP0+
YWwremRe5fBDfja5HK08tAe7M6VGXuoDJdT/5FxhUoIXwh48BVM18r7+zAcy+AI5uhE0J/adu9Uv
F7qZZHAIgv3WsWAwbrAzxqD/pyuMFF2UUzNshYUHREvueEKoHIxUK5nGrGYRXx6EDvkSXDXlnCyt
1GyRraAf9gB5FNxJ2ovqhZYy+Q31Dz8i33tMP3E3rxuH4vdNCnolRbPnhpwXN75O4J2ZGdDhla4V
WWdGszKlcjxKm7BUZLiuyH4/Wyknlw6VjimScFAY+1jbqjj0yJvYHOH20fX2XDMD9L9oQrCSPHi0
wYE0/X1alnvYz4AFAA/EVsx+bQB1DpJ/aJ6HTybOJ5Y9/XaNcB4fpdfhW8iGM8KBAcf6poSa2xLX
Ie/yo4UOsvsMYBUc0qPCkpm4iVrJDcQN8LDrnZfyeZPBaA+Ljl6N/A7Ntstvl+Qp/fNS1EI3IELH
vuf8O79tQDi53xJ/3m9d9T5iasT/1/5E7aWIdb1ZwRLAgMw1W00QE5TQtvUeEcuE7gE787skTpye
qXmtVSXIHUx9aWqCt8cNkVrKFfDxs4LAE/5bWSr05DagS1mGarurOoKBeDHJYVCUt1nm5KvgD/JX
NIzoMGHAnarhtcUyaZwRtTqkz0Sbl7lmds0PH8lcGc25rIdgHsz9Yb7wDpDXTUVFiuGN9bbW0v0X
t564yuTojqgsxybrizRppIJzDyBZL+MooCwVGDiR5iPDmXad9Me+BkZqoJKQ0ZJdPms2SUBRBSrw
vp40t2JJYtapR+fwfrIShKrQTRlrHuxy67Yg3qR2I6oH6LIJV/Gkr7Fd4FLw5I8dKIUK/IsePv4r
hV1Mm6kTs27t/ldK8qWgHZPEYP5iMaN4VRY1KYCrPs5WqhR2aVfHViu3SdoIo775yIHXAyT9GCc+
IXmybqnX+HjzZXjQg4IqSFGe3/qJLpXyp57kdKOVogzalhy5VyC7vvMqlBzmkCV+ZIb8YeB1FdCP
CZXUa6PoPIMRzF1oyuosF8MUHFG5pPXlfgnKSTsIfoBVevQbRcnSebVoTUaSIZpAdcCLXEDdiVUg
UyS0m4+YUSeMRTNbLpzDXtxgAI1HDcedujPsIfaezBTHV6nVxzWBYw24UhdY2bLxj49rAKZKgk5S
oYjX6Y38svnLOY7vKlr1oxVGU4pwhwz+j78tk+NxfIwLhcew/OF1PW2SRcJdyK1hxcFMmJMBb1gM
T0+MtpEXERHugC2F3nt8ALQOjMO/tRMhd6INswiMjTDd4FTFaAHRuj5rpFWKGWuH03V21JYdfTwL
32FKh+xPtyFJ/JtYZnCQk1odXaG6pFEwnUDT9aFr1JpG/0CeFdNjQFLmN/jRy6mMYSK3SUarsKKy
Cc7atFx1C6wawT3tUtpbv6EotJIe8ia/+56lqyLD3A6T9UMC57meFOpLDZ1DPK2MP3qvvx8Kv18F
YenMDfzML16AXHOwXdX+OY/xggk7gfOyei8C94zNryxMP/SVQm527ggpJQxToJ+B1BtkFkoEjJEa
3CxC+1u2SFYvEpmASVvUkjdaAaGXwKWuqfU45gsbfUhbmWESiUey33iOpGSVEFE7OwOEa/0gzw9g
iTZW2L+d29XAdOitvBsgfylbgMDsjgugBQ1fVPvYaDkdob6NwokhfWY37Y55yvc/3Escl/byxqo5
2S46x3ZuqLhSeOXjlFqJkdhbs6Z8aPEOd6rIGbZGTnHDCuPdtirm3pN+3bkNm3grP+TMdBSllAwX
Qo1s2GuEppg/fCXT8Y1pVxWcnuVq7OYNgEex9WWZoRdhfKwR1n1hiDxE4NVI+9r3e1HUrzTKHi3E
WWxDaBOek5eZp0O7VuURfGeGJd3xOsU4GXr4MCdqFzdzt3QyWYs3Kb8VSjwqjltAhH75/soXYstR
v6xU0gkOwGZRNIKXMw4sC02nJz9GB9EM1R4IHx5CGTnJijILqiADPdJoQimCRJSzZKE1Gjrg+0LC
Nuy9TuGN1pe8GMBsLepnPqU69Ozgl2mDVIo3GN1lR9F6bo4pthH8XWCvF7FRm6+csse6knA4KCzQ
QcDkaCDsONxqwkRUZe/qeWcRS5jVsa/n7R5ocqD5VsnTpN4Bz2Bm5KbDyYgRAMg1ms+BbF9HnlYo
eq3ypIMuZWl9+QfFR7qM7Rai3U/NcJj774gJblhHszRixE1dzMDwYVk05UPCMLqG0sYoRPvZqePn
1MvDwjH1hSCD0GMafIjoe7Bp/Elnth69OIyl5gknvXhYDLsvFKOvNn7h+JMG7jmmX3Gcp/Jcwm+n
SyXloADyCy8xfA4SmxBFZ12ibOxx4kDYPIwZ0ROYHiPKszjgDHmGRAL31pevSYYCCWBJXzsYqM3H
xm+HfySF1MVn6nJymVBR2QmjtOR+9erlIfZpFgGgBmFqZXDl0dgNthiyRNp4WXSf/JnSWwVCWXNY
y/+EPVcamOxkUdLW/oz/ArL8lgeg7eMRa5OYkq5jbQXrLwJghq2LIzJqUBf9GDHt/MZjhQ8FhQVK
PNVpTa/b9mXtxQzXwuWLGmrYfMvUheJ4llY+2fK4uOGqPNNT9TS2wMiebM78IHkyVCbfdXXdRo9h
LKV90e4zK6mTKOhadkbUTaKw2vhZRLSh9dQRoQZJZJQVsiB+a3JcMUy0cJWVXguIbhf2y2AQcC0p
zdsdg542ZJmNwd44vhaowh9aIjM5OLoHPkw4tQrLRodVQx6faVQOGKaK3GjC+W00O95BwM6N12Sz
nUmkKL5CsLBitxA0SPCoErsim0RbDC6MExSgdaS/lnMq7h/vI5Jo1CFHrUsMooY67uFLFBR3SaAo
h5367nRw64e6Lk3vn+iAkQiSwcyUwFi61ij9QSUsV0m38El7Jg/vVOlGXNCEH9/kmiQYxaor0Z+1
T3MvWevQhXYVTFjBTJlIzz23objTzHh0Bz1iwiL5Bsla2UbEMb8haqM8I/YnqEaZN5bLoxrmphKz
jSeR+54rM6UCZB14AtzeIjFpbvkjIR3f+X5k+53D3CKARsy2M35QpwQGIKgSgEqwjuNOWrRpclN8
JchGpNM4ekH/ESvBDMkcj/NyRT7bgJpEYUhdv+FW/fFOlLuirN3aAw/i3nXIAu+thofEhnJT6n6r
O1NNR3CjQw3UIm2RZuJ92PG21u1cTFjglut76ODV8nqS7YhgKmMY9313ZSijyhETbwWq3mPWw4M0
WSQ6bcOI0CX6HYwFtn7tzyrIVwNg3LNr3dkMnP5t9t7pXiwH+o3hdDoDeH84ohxjBpURO6IXF1aj
nuP+bhjlAiuuxAjMzn9gz3Lv3iu5HfSEI1BZhDcg+f6+9G8/jkxRpvrJQoFclx3WfpNiIQcDaHer
LVAAeg7Ws3f1OjwrrJ3AdpXoV4hJlXg62L4M1HNkSVP9GPkPM2BH7T7e/99+5C8CK3eYvV37Olhh
2EVHBEwqTSKHoYv4iR/dy1D5Ean7GpDLcZZfcy6+aGp+6IeNUWe1welwcA90uajgxe2HHsRdz9tp
XOExzzfziyC96HWJn8kHRrx2lrlEg3SaNo/D9eO+xzn+vUQXHbyL+kBbT4vNKihvKAnoErpDd92V
E8mOvhoMuR1dkr2LVegxdzDd+KD6MHyUrHA9IcRTNAHHgXcg3r5U8C5i+/RjSa87IEBj3zFKzDnd
ZjMvzbgqmD95zUXJEapTulvCPYds92bOyuR4luxDzOcYL/oaY+nuhXTRIaMmrjoyl30HMFmA+IJz
G2ZrTkmw5Kf5YSSsSMRPzcWYuqhv630UXAZG9K2WRZXVoMRYR/jSbB6FlcWHNenWTPBtPeru2oDS
5UuQwmiool9WyXc58w05gaV+l2yp344ehA7hTaUglL4XrptC1q4FERD7ygWTswgxHXtFdtQCxLzv
0o+if/U/WbQZRbUH27tYc4yWutyOSDldcFCT5+PixZDbir9DreTjyvBsAKEBaKumiMlL+0UMYIkV
K4KC4u/KG4kJOGnFpdp1aC0PIr+05HmGqpewCoNV5Z5gjrsju/vXJj2dBcCmnlwh6NvQV2FwnGhd
Mu2J+IJCq+FfpeNURF/TR34GV1A8wMRxXjaq0WDAAnFZCJ69sgzpR/qmtG1LpdF4znXaFYaMFYHr
xjJlFGejFCIw3NZ6ZUX8swe+Cq05JYgNpvCDUA1Xgu+D2n9xkLUrq30nozRzKdgWk5Jp0bUaGjn9
z8Pf6KxZxYTuGyG1tUdbxGygf8HToHEDnH1n6UWnXfbKeB9bbZE/pVfERuhb7Xp+duplxX4Csnkc
1jZ1MWML9ky+5MyhD5TXtbi5pTmKpwGuyadokvMtmdlA0NVjM3GFzQUInRuoLfyJIkCckW2MDDP9
cwl/vwBqTjHW/Ho7flsPfkpsmUwHqbDnTg6+9oasB0PCtpfZfcpXScwHUckkr7fC/RQh1oXvCN43
MgnF6hrF0Ge+hdAOXSbyg6UsngifxdMI1ivLPob2/uSc/khdjsybD8j6LID6Wxi8wSt47falQ+82
ndronmeksbKI5oLfzWlffl9UgZtgnvPuCPnzTQrbRvjkEPyl9F1+Dvg0SMtsoAbuIMhMmM9TfVCt
TUAep4Tap+GthW5gmx/Mx+sI2uXIZLJgcfE9KHE6OcshVYCfzr04LG3mS7JqNhKsoU5tRcmVy1IK
jobOVYGPa3QjcXcggt/X+vOBR/UDqC2rayoMhwifHpn7gm5zgaYn4dOyJJ6tiziPQJsaQSIcX4Ed
4dMjEQyIOVkjNBPYVB/gCG0ARlCMaA247R/ePB+0oI9UqhjNy9HwURykoDJUUIKSFhyIS1T3fqxt
yqvOUnkZ3O5f2y2Fs4A4IJEtkSokLfjzVK8K4NDwUJeFVVH3RNmAO5yty5xrp2hpM4kIvR0x+/b7
xS3I1HI1xFGw31+otXSciyp45cKLXLbmJCQT2CPf8kHak9KlXZbpoYk85uzQgjYhMFB2KZx+pOk9
MPGN3fP/iDo9VHqc9GJoll4DPOTKiOi2escr1SHvOSKI5V+Wn+z2IsVRdOmw33myr8l8VW0Biblv
CsCCAwCmjwO/cx7x0P7oIfxqBVcszApO23v+VA1cd0zt7pk7VY9LTUbghvrv8BzlhwgOgaOBze0H
aYsxpPNyFsCVLrmCfJQx3tVHWjo8xk+weacVjeDjg0iCllFR02284BBjqpIyDJMl0m9qIplewt+I
xlYmwzU9nlm4d73pgi0PwWJfmS1PTSeSHMzaanbERZQfd2/rS+blEGRFG7aPqH2+nN78hckrHLod
oL+TNwCAfqp+tPLyIZUlIIzrExMoBmuE9lldtfUEmPRhObdy21KN/+Y3HE+i7EvhLEjE3OToiRTP
i5k5Vk6CXGRXErH+WLyvtk0PFhXTOWiCaLIPdtHr62loIjTf9ykupzgYZTScmiRWphwT5say8xhu
gpDpL6lv9WY1PQXCYtkuT5rY729xq9VghT5AUBir9jDHHSd/NgdPTKHWf7F3qJFIcfKT+JlmLqzu
4YopQlueIzZSDITXGYJACi7qyr5DnnXGOMomd6yfVU2Uf9dnv61pzijf6a4ca/5c1fMxbLZ2kt8M
zx3m4sRXCM0SExw11kyIof5M5B5zuH4EZvaz5XdgyZ7QXlDhR7jbrMIlpXHcihDtNnrJt/J0odFj
OYUstddauEIUnNCv6tHhHpC9PzFVgXVgu0byWyQVhcIgJuzFwfqtOGRK3+d2suMlsxrGWP0/mb+y
5lSmTmvLa7mG8f3dB7TrdIkHbbPhn8JDSoLNytzM8PxSOBpz7GqLYMVct8ihFOacqGRYmAxlZ3mA
2QD/B52kfB5f7VaSnNcy1ScgX4j/w2SsveQNMF0xzt1FjVkiF8ff8olH711pXtY/TkCucmxBk8IM
CYevo8wXF5tusfrLvHeN6UromoE4J18In3T7LRnACbrfQb1JIzXIRxGrB+KKaPPpktByye0oUL9V
C6Tp1THSYBwbkTPT2kNEWF+K4S6vnbBlStRzwZkz6cRERwulQ7REkQi5nd/ucKbBseyCjORAjMkA
9AS11Q/wpeoSOgVX9fne+9wufMh1UZqh8+nwRb/iRvOzZY1PspAA9Ijuk+ayKc1G91m+aWkUxArF
lBMCw0YocLt2I2QObHeFTJmmhT2q5gtimUm/q7ETO/jJCh9Cz71MYawI//XzNfDRrwDp9aCO2jtg
xhHJUxzg9dKE2uxEnKMT0MOHKW5FxEHo3p4ekyLG3xY5hjdzlTldfLAeUAoXVJsxzuoF1+u6qeVS
1PGZDrQvABGPHyYZ+ZGKUylvqL4fg9jX4bkkY8K8WAiD4P3GI5KaMRrtUrswOnki/eosKauiSjTE
w7clzhhaGMJeDOxfPtbXFVAbUvHYz+fsX+Gqm4JJdJ7LdihfNT1CtYQvRb6k0oTJySNy0nFFXXxv
icKbGu4/RbNEgJMXbPRfXa/VJ+oqYwI45cHIJbJiBpaOgxLC6MkTLyszqP6ipMMP0VVjLNh0m3mw
WTkfNSS5lk9MKfVGhWRbb0L281XvIMhfbyIl5Pknj9JzzUnnowIUmVA5Ke0X1jeKQlwcJ3ns6GXx
/0wioz79ATkbJX06XgtGFXcXidgy7TFq1N+0akGovojlZjsbwCjBThuUpooSvoT3A6CUB6ji5s9z
80r6efYUjcQszWm4SJJCIlhd0Ad+g1UGliiYgZzp97u4MiaqWDBpr1A1AAw2ygFke/8c7rdzwXqa
9hGZkyQqXWsV3fH5VTt/rZNzBLsbVY8IYP6fAWkTdVirerbLbnOs2EDKm/ql1QYgny8vvmtafp1J
FrcQ//drFBdSX5X7ltGdW/C+xwzy5n68cnGxKEf0Ai1VDbQW4kvRwxXAEcwEzsl9g7NBaNrYhMqS
//0vBVEyXJQicSPiPdypv4GhURzaMkMJyoe4BHq6V0lffXnYqckVbXTaKLn/1e0ao/7ExPEDUlnY
wv6GRX/7JfrzrkC/9lwR4W0qUvDo4tmE89JHm7ua3TV0s3Bje2R9kfFtbGJ2gvZ2YqtkRWSsNEzJ
9RKYTJUhjm+QQnPXEU4lDWny+q4vC1PY3RO/jrWQkrmNVKMU05macMmQuL4tiN7Jm1z+OfzN7ULu
FAHfal7rY2TJuM2Hg0DtYkaGGxFwecQ8JWeUTLFw8wzzZiGLRwT6y1zoglKfGyr85THjfDOFGu9D
kgFTx8P8uxkwiE8a4LGBEzAlGxQrzqIx/1RB8fGQ9zlhZrrgmu3v3SbLgBb0kqf6hgRtcHEkJ/9L
XwdtgsBdP6WZ8bvVi5sym9RUMD3C382maTwCf/JuM6KF/KmDZAKyg71Fhyng0VaJxpzTPhOs+1vE
zaWRHLooTSdx0AfGqCWtnUMfNQpOO83yMOuHpjjWKmzCjXZa8FHFKr+gGgGXEjmBy1HnAqiWsg4x
g+TDhUV62uGnG55c2fXj7rTJqEdTCm9EHiJUZtH6Ayg6gOwr3p358ZaxZGg4weuiUcco9BLFDoDB
PiI5cB9Z8qJGvFck4tH5cXpC2CRIsQ6nriUX0Ho+r6Vkrzvq+pdJru+c/E/2UlmQEKZ54p7ev7oh
ohlByEdTaAVGDYOzMY4jcj9a8lLmEwU4gIY8Eu3rorrwThNljJR8Ce9cLHO3otN6vivTqCHYvcwV
E9XQgarZDNHwVsYJ0Ebpi0otwYFTOGt8SD8yiGhkYhV2hpjAzbnFPWLCrhWCR7vaDpjfKHNkMOT2
2LZ9Sp9HDszphVEwLTTXyp8ykpkl2xvnfsm/io20StsJ/MKzoEFKj3YTFv5JBqjum/AFn2msiVGa
1CwCw9gydbBmb7lmYLPEipFEZ780kbQzbKzWp6GFa+KS7rzVS6ofmPx4UkxaH+wcebMoJsEEkoZb
2lvVcNiu5Qlzgz1oOTvG/1SWMJ4rQEeHvXWTN9TX5PjVWd30j855Nq5CQnQ2a8+u+SRqN6G7bXTP
Cz4axQqLIR6USQIwfvoZxJISO9I2usqwV6LKu0mm3dxP5G46pXfhQSXrHYuO4j2i/eDCvCQLjkYu
0G4320nFfhkxDTEqhJsao8j7m+UQpQ0KHYPOYx4u058P1HVW7wezVyEr70QVte/oomCdOy2t/IO+
Pujg+nbZ8ZggVJ8v7MK5c97DKLzWIQZdtaC23urvmhrk/Ap9RRF2cPXUJPK3/d0FmuODtvax+WNF
IVLcuw6n2eu+EJ0JnX1pxyltyUEdJ6ZzhYElUJfaOC5bnC0pUMBKzX6u9hhI+Pe9vO95KDzvnNd9
AMfHiAlajgRf7os+o+Bh9zQep2slNhMzjnvaRVWbDPvkK2am5uOqXr5o/7YxC3d7AyoYlUfq3uv+
aRd41iHy1mSAHrQQaFUUiQfYbaVTgXT+td78i/rsnMaZcjqOZpBQtQj/zaI3pP30sM5vNcV6jgxD
7NuWBXZaHwo+a+C7R4gg6S82tCm4FWZbA4qaVDVJo3vVqro1nEgPiHxCapU5fUMLN0/vPel1ewJ4
+C2eNPiA5Dfr7Wgksy6E1vCD20PnEIV2AjG2/QcRD0AfWZhSIErSEKN8ysfqEUH+lZWOnn23rIcC
wFT1Nb4yZ3YaHehWPSCdAvePXfQuX2D/7dgwpIqXL+InkFxyi/gZQJvm58G1okIvMO4qTQ6qm7J3
Aedk05juSPzZXasLQBBoOyJ9QgJt5jcmMWld2es1gjs6IURZxrB0oqN0mrkYuTo6rCPiB5A2TXN3
bJyM4iRqZCjwFCIBNMlWmOj3TPFyOKeSWsiZM9qGCwtitjPFRc/MYsUgoKUB0hMTYJibobUsu26u
aLfx86/qHUAAm0d6wkP+SMBLX59NzotTkQ+XbdeaImoaUqXTwtmevbF2j6b/aHXz4vO8NZam+oR0
L1JHV9Ft8H6xdwIyiqyuaL34f+bYqOe4YLNxmewqGTlGpS+nwHpA6SrtISyMRIoeIFYFMZkVS09k
yv5SvoLMuBPnjRrz34JyOj3Em1LMIKV/TzmeVKdvunlnjKa8zPtREKsFqvuigi0OBDzMtUJsbUXD
3nCv31NQMtvhX0+emais7QKsQ2OOcLKrxSM4QgOCe/Qap0UXb1l/5Pi10dqbyVJJAj8C2Gn4HMrr
5tyMnsGEAdBL9U6hi41pW3bie00c86EzXC+MV4cz7y22IOl8Ci+tye11HpfROdFP6FVTmM80Kvvp
+7e5wFkqOagNwRIxKp1nUs1snxoLZpThNwtd5Tb4MVCYVdF3b/05yfrLDZ6jUlXVdv5N+KxztV09
Jj3j9WsgS+K3o/Ohpe8uaEzaRIcJmkNe7tb8kXku+mrG7n//N9d+4NVEzxLHyrRxMJz+H8RSnFVO
U06SYEc3oGv3HhZNnlV2O2yOS9Z7q5Bi2BrRQFXdUEwY+aK750y7eEkdVhN5duwvoqjfrZGb1/lN
JdWj0TFVAy1mPv+0mSDPN3u8GYSYKMR9Awc6bm+rgCTdOMIxteN2uwCpeRHFNdHb4JcCk3kWw9Xt
5oet2fszfBNcMR94qcXVyKzqifduozaDHoIOmcq210B4JQtbngDKI87nBBjOy4nAiU9DLqowXLYY
ib0SewSVIC5/vJUUuQTdFLKLz7PnpE+UgDbTLmQNJQN018skmYj+Mi78Y626hEsqbBEbSLxynwJz
IYCVQ4fig/MdJzaB/GUQ99shkbeYPa/4jm+JmvSXC6FOjoh7sC6mPb7RYbM8IR9LB/77z4q2VYPo
2To11sT02LpQrM3k3WrNmvFUof9a+R/r6rn/HEAsYCsjpXbdrs15hB2g/xcdevQYwYlY5WNYcPsD
JdlfEnDttHt7nv+D2Rmr6omEuZTtpdlu6olpB/ph33jFMLxdL4Fp5WpmGJeusxO6+12U7bWk9wBa
Nwp5gBr8nHSE4/+Q9A/ATlmfacfymbjj9A7t6jolvIo8Eaw15zcJbuxYRRSUFUSPhJH8uI2axPHy
sDfSeHvftzb8qPSNe5uv64Nby3jtLJgQ7uQ/SGIvfBE2eTH9X0ElWZV8oWFpxPLK7X5fvxJjSo5r
AkmI4GfUdYYFt3iLNeWsjnmGO9fq/682rjyultPhNmPfXH0yKY/T2uyJwgN8ojDQsSogZTgrm+Zy
uDFp5O6+k+nTShbxvVSpechxswQauWFnvPXVTz8oazsTU8ro2gHcyIH5aPgEdpI4K4sejhFcqTKO
fjEoGWmciz5w+WbIpDlN2gbC5zsI9A0hNNOu1+L9CGYRaQvQi7vQHT5eghlSytfVVtXRZJf7JaPT
Yc5jJ30cG50ROYXSjZyyOndAk3QhhYFj5YRSG6Ett3dyl4gegmd7vLQy9wMYlZT73vYJ/zpd9NPc
7C3s+a/uNkfAKCOOZ35/kfXvihVJ8RZW9GgNiASwUHz8f9qmTt5Ck7tkHLEkJlEiMJxwMmbvuDm5
280egVV3EXNWCr0rXB7nt6hlyKODWyOHtNn4lOiqtKRXswcmegmC1ef2By3RKQ452jfeEPqlkmRf
gB8t8ueY4atpRL96Zhixeq2NIOFOzKy6+7DEHlczzRytFiOU5ceFR2yxmzUdijMD/wChikrN8FNv
PpMDkSo/YcTPBdD0fqub53AbsgGYwki/e3rZ6IyErmJnib/SOMM8MPDFP/dcROqeS5oXg4cYwP6s
Nnp2c8jfO+lJ31tdlv9ORPsJr3RqyR3ry90aXRBH5ioc2IppAN4heo1YCRSlhzec4s0DUg1k1xRw
8UCoHBOpl75j/2R35QRZlPv24Uicb7+1ONIt5MFIyrXgF/iEXdIDXEeUDerHEZCPhtRk81wRA4gC
ocP0lIXHEbs6Q5VdeokUwnnTOP2jxxgYI+m4SaWlTWF3RCxZoP+VNKIz33IoNfw6Rqj1MljPbl62
8V0/gNqMke2xbaE4+sRXY+ZOX+GMi8neEtEhLw12/EsysztX25nQ8Yjf6F7o12bggSpqMJqvVF03
m44qSK7ckD+7kZ5cNaz9bI0iMP2HRcF8v0snKwdQ9QEsHtFKTKfr5GkHgux2ngLOSKKyEX3AMGas
y1TYjCJ4GT0TRi+3DYLC1rmv9ukUBRV22imbisWrTX1xSJbL/p1wJzS/VarYAYo29wmErDXhYVwL
bM2zuyCHt64nnobM1MGqCr+tQ0cc2EK9eL+l8pkkr+2TEiB/xkebPpA+ch+lItJbR+zkOY4DsWAa
PMf+9VXz9MGRMnF7qLzV7QiIpjW0VidbTqXIZX2qmDarFTvlrl1sVVWs8YkDO5QNGCHOq4H+9W0T
T3RHkGQ6N6MuEFX/6EA2q6mwBBA1Em5hcgqkapPX7l4dWzFOx0SeD0FYdG1zV4co+gOneCEJ/3V5
cLQRdqRfH9Ni8pCELblvAislqjQCS3/PhPmKTXhkFFp4rfmi5F3wxo/xgP55uqvE1dcCM3NTXeQW
/OfuJHrx8/+KzDSRyZ+6tOs9v6T3nwtRjrw/qZQHPRaPs174G6ED2cvvDW65K+2mxHjhBAnb9HT4
yFvP0j676pAXWjyK+6WKF1P+OIX1pfnSkGozGEIOT9Bhuaoqw1GAE//M6LZ3811s+AgKi1RvNNud
rCeDhI6yAoZgvuN2l9EQ4tme6YkKtc/w1E+Zrxan3ki2EdiClMkQnqiQfc87wi8T8yVTprQGoAxP
p64yihCx5cDlH84yGnJVYsvxdf0JzmykBPO7W3xnvUBUvYh2KSkX9wIU2N+sz68kVYaM8pKoM7Zd
mBYeIzfgDxTDRVmcauJHwz9zE+Oz1gBgYhxuV0p3YgF8lA38jrer9Nq5loSzcR4o4PKv65vg5jqW
iv3yslJUoGEH3eTdkhg5roXFWCMrOp1rSnDu1YgNFsO6R51lfY7V4DHnLO73GFhiHGseN8urxzPm
ndjuADIZj0p4OX95bWVXgRacJRewG6ynHintRizFgx1TtDV8rEnWKqTs1YIsapGyMV/kzIPKd4hV
hoY26Lh2W46DGdvL68O71YXHmkg8SjyJA0Uw2cffu2jsxA9xj1CrjZScLVLBstOnkTnAuKB7q+vj
UHwpAuLWdIib/xO3H3tcfhL3PWdClif8q+Wd+Xf9MK7aob90bdw1nIn8ws9mb/jMy3OnhMH/D9oX
IYdUni/Zft9g+5iORqsXk2o+CNm8IUxBIaAnVqj3cmI1SDmo0FwgTBxsUmpS6CxGmReqhOw2Sh0s
sUZHWGFl7+uKl91S6d13vjy8JVU/l5DYNW1pnINajllQw5kn8OQRKEPHBzWQ+A1ATD8SDtWuOqz+
jsRGtVGDRstAS7Tg7XQ84h6loBiCSJvcVTW50EhHnZVtU8EXN126HB0BJTGtn+raQOPMOUByY6xF
XXMg54/W1zbxu8K4blm0v5k5O2fKlyYY/cN1FkD7F9ue0UfdGkLvQ3Btf4oGLwTDSkkhn6o5srlD
rX3UCoikKJAtZMqys5kxIP6U9X7IpigdW7bbZdtp50u5a2pe7yDMntW+eB8E6CTemRCWFmRubHQi
Yt4ne/3Cssm8EceRzjSaPv04KFmnoOwS75QnEKauxu4LFyo7ikuIMpX/ETcVDMhcwB4GQ7HAl+wB
YEJXD//CVg+P/kkUB0LBFbiffr09amC1nu+c6DFrqqJpi13aBSIG7kHjnOrJGiPAdaBWOaj7f1eP
QdWXBv+gVgWyZP9bOXoSJH9+/m1mC+DVYgGls5pWicnmnVJOnyczfakZuBhwy8B3yiPFu9sfYSqf
xVWZjRXXwQ9aWTsE6cGoC3htsMAiX7PLFshkOKa+TIHnBn5OUxNBGwKbrzQdiWNX6aa2ZkiYJsVx
BJe+p5eERYr4G5jJgka2xdddehIlsdFd7IsMou0WZHIA7M9BvHTIBKZ4mGHXMpQroOo2cgcWvZN5
duicTs4qrUPjLSsvNnm2UlzrPGi9yMfyRWBmSsfms4bME9hL+fwPc/v2RDSUX8OGlkjwdT/V5Gpt
EjkGGhe8YmQuAhEioGWXvQ/QvOCfEEsw5eCf/JrD1SYAvzqVaTIxBkAIxguOOuifeTELmcgzTk3h
aK3TxaSRYyKob7QWosBSJZOeGHUnJ2DFbuTFfPTXUOfQICxrX+h+jEUiWFVnV029YgqXlMCBZzc7
PNSUFpddscxlhz8CTVyVfObidauCe5/oASqy4O45ThIO1kFaesDsmB/Sw3w1qAGzrhwxcuf6lXDZ
9lGwrmbSBW6S0I2uMTQZkhD8DElTRjiRJcEKvw8F1OjHi03L4za2nf5/LSy65NL9rUB92zzLk55a
FqVxhqChT8rMyhqMyKaTy7EMFzdpgGfOX1Y5ruqVLl9QZBUNJjXlcGVVMMcnQ++u9ejD9IlPyW+r
7/rPULtEDmlgBmckGNberefx+ZSnvCBviBiN6/rW0WcPDerZv3Q6wcBW9jXuvokLtDyJG0wRJHEj
Z/YIWFlzKqZ+z6w7zZ4WRkmTh6S65UhvS7ROg15BS1I9xZeybL1arVWiaDHtoaExZNo1+WSHG/Ja
+PV/VcvM6Mq4AxE6yKXOgy4kDi4QOIXwFKk/l1lhjkHWZuPPvA0sAH5sCgP9e43M/oxpA1b0WwJh
h6MY9ef5O6V4T9fUvWvUFiY8mUuWAoWuOUbhTYggN1pFyC2Zc0DRPwQPqB2tMEBP4wBEu7c92wyK
jjPi2TmefSiFvYOJsI8kzUxfhAq6njH6I3Q9wlQPcpQp+g4s0f+LigCXMcGKLbZF5ip8X7NHYntT
zeG7xAASsUi0pEGBBgmHitkYy2HTR0A9reKFwssPub2zf+HsrKKU6pS0ZqcdN6kA8X30qgUTZrUN
+mJQQCInGGQCeVw01MjV7eKy8Pca9AB2W0MH+PkbdEZHKrmsi2EySCMRBVH0pBOM1nSSpcDUHbJq
hhM/wE5pLBbm0mcUbGtEGtTz5y0uvjcSFD56bDw5qgSTxx0LMcE095h12XvjFNAAuyIrJUeKwpOZ
VeCRtQQp4Kor9RkxIIB7C0MmtWQ2uEdBe6AyjXgdpDVSpRwUoxLxmNXma+T4FfYVSuXg3jsJfTB7
xJAv66nKzk5O2msswWlX45F7U9qz8BQVKU30Wrw1Y6TdLBSNs1vKM2pJErPtE8xbjhOB344bidbe
AdKgaVcWoUIxVL0v/MkeVvxliQC1eZ/EnGvqmrrqoGoO9N7SFBwpz57mkkvsfE56F7zsyJLPUIYA
/lPeOql4CNkiD/Eb+n5bhJPJDPAZmZYqXU7SmlMrRWvG2Yj+pvCWoF/cu72fj2xaKHDNZmhgq9Qg
z72UJcNLjxCHRp78R09dE4LGQrZgrtN2JZnRU3oGOsZ4Ax8Rhvsj27EoZk9bbWRO4XuulkmSAGoQ
gmosqkXahawWWRfF3xo37slbplN1gh2iHf3KWn8P6EGuqaBlC3sTdqONAp4V6v4tAO4meBhIc+HJ
ecGQlIdBk4RKGLc5Sm7WLislX2fzRRGa528nOkNml2noBZIRIg1exH5PYimlcsxw0JqEkBMeKySR
fWmWvj9+J3m9uidOKdulzTCq9nnu2h+chG7BIBl6KnQebNdDzcoOJ0CRcz+F1vhQmUrD/aO6WrlN
m/XkCt3aJVT/RX4D4SUDpueVOhT8i0S5C/t5dhCojs3gATn2D5EhZaCVe1PSVuL2NGllG84GnHbh
baMav8EGYCweIYxa5MNnCMqcyy5FiDHTVfpq1EavlGku3gBtCFIE/tV7DP7SRyKSELvttgDTiB7m
i6cWSjlUN23IzF5R2WrQOSipr/mNgod1b3jDiiYGwkJMaTbKjTPeWiXJ/nDxzs8TNX6DLdVZB15d
xyVr9nNS8RCFhcPJmenuu/ApOOQdobevo9wS+Y251oP2yMj/30GN8GJli0TNRgYM9D3TYqxKUavy
bW2pg/Elq0QC6Pxy4ty8BDdK6WaZ9n1k2sUFSql2qotJvxYKZbl3hHagAsropuA7hISgBpRlq0QC
73AdDHa61yqhv/QLH3FrkhnI5mU/UJgAtBx01nemNT9mfqkkx9YbYhIN8boPh2am1tH20jDvdNNu
/9gg98kM2+eQkdGMFOXw9ZudzJtsm09ZQmVV0/bsTD6p1mbs9b7OJ7+SzIbumZc+Z9J0cargeI68
mCUhKGo4gBICdGuuoXQ2rilYxNKVMJy8vMYnoTjs7w36knNZH+/4kARTcB/u6e84PPzdxY1/wdP3
1V9/DwqtOjKJpHPshFgHstXNmxZd5l/xXg4VaXfVrzMP/RhLf9QIU0po8IKtrWGQ/dRqIWxfptnK
grJ42zmwBqV16Z1057JbGLH+mtAoS9wA4KdxR2ykPjajDgdsmf9Spye/mgX5DloAA4DydG95Q++Q
L0CLrtt/NQXsKkaFbLmFJjLfjmcmpihWgKoPp2WQpl1VQAg7v7ouBGvgdN2nRQWPfHVzN3Qza0IQ
x3j7wqRahO08Hy2Yy646WmYN0fr+o4IPeQgcQgwjEhA6FkkhReJIPdJ4JhS8hCeu1LyGbGW88miY
UpsDo7PDCEHiFJRw/Vwz5d0q2gFvtSkHHLMAfcDnAmHHz/z4oi3TgsKf9cfNmvPNoZ+PsAyeddN1
S9I55LWKUOM+V3PWmw6Kb4CRVi3/mu03+ZurqbVOziY++OhEhZEE1ISCAWv8iTpHBM8+luSYal1F
cyxFO6NpDap5mf5At7eqc3XGWn/0SjYqNp5hi37iNEeARVjeL8RQih+nlHwvs+SeqaHeqx4bcbfe
EMoNAK50c1cEi6Y8qKIydH62HX1YR4bgxI4PL99gGJKq24OwICVbGVYliN+Wul3S/D92YfpxYxMf
/pQwA+LSB6hfJ68yS8Yu5lcuiIbL2k+AjUf4oyLMPjtxud0TXrg5kRyKrgT6Ckzx8GIcOc0nUW+R
MXvo1NbstCkKq9HayIi7fAR94kEBHC8pli/OBbW1GccbUiWgTbjGNztbP2NzDWjyIUcDENvO2aL/
k7UJ4yW09D4c7vKS+w6U1hhj/UT4sbTH5+LukO/oX1egZCyWP5L2clkWJ4Javl3/mPT5CXEjn7DI
lfBH1pwdrnrtLanigs8N6Ero8+JTodZUUrpz6yKjKjhtT+T8GjHwTNKg+ROOfH4T9t6RJAwfjPWX
E7mV8gkH2ziJ4B07hUjPzdrN08QojPubqKamso4eAlZsnkteYZmVBK9aLtN4q/F7kCQNHQy1eJba
VBWqnD81P12iS+vzX06HlRg3RDUN3m7nVFtw3EMIRVV6PaQ7TqHFUQXoCRMtGloec7OyF82Q6Lgg
dcvSDEqZA5NSDRaEAArBfGrNr4RojN5kOUvLYWdlF1WKgMyJ687pXsHJbxDAbjUEUUcWVRhg1g+v
ZOXo9IaWIrI1ke9GuWlRV2+iFqqW72O9Papu9jfLB9bi7Ho9kDo0M9UUudVzRE/JYQo1ATfnwwHV
8MEE76ENCBHmbiJez4E91MNoXwZa4tjtJb9UnlTie10vrYC/qkitz2osLAUeDLkz5Z0+4Dj72U9I
Jf36YtGwKsvkGSLF36cYbMiZWV523Io5qHd+B+UFDBAlzqOiLjJLJx6oBFgI18d5YMgX0cs86nzw
pHFJYNWUQh+yelt9lvy2aYPmbNLI4UTgJyp8tCPebgaeYQ6McbZXNku4PrBBdJudEofQ7fxPkBS8
A3nsHozan0qoxQkhIcOEGJQ3sEWqumh62OSNTLNOoNt2bKZERDz1P4AZsJyyKT0FjLez3MhDxjRQ
+4FOFggJMEnDf3TGbfC9QKrjpIr8H7/J34jTq92SQfVOuuuGMaFPVB9IsaQCQeK307KoQ6m1iuWm
yvvORf8+6j/44MLoU3HpGozDiScwXX7dJAi5jhsWInOWwM5ZB7nDthjpoRR419TK7Edarnr8ICO+
KivaoWWaiK7ZA7BYSvHT4dCS7ifKkBhHDqXngfOcKHt2D91HnFDHHjrdTFqzBOc9TamvTCn3jCTe
2uXy5+IQBjmO1Iy0zKEq3aFUqBozVjFRRhqx9CkcVhIYbs0o592kj/8Bo7l97YS7Y3/39RN0oNAm
3A6VC8cMPf9BpDJV1464QrdH6fWF0wdpNiknKOrxjE02vnmyuKivz2t9Tip7fLwmfOc3yYHmgJdL
n5xxpKN6ZjdsQElB1vpcJe9uKGi/9uK1AtLojrnypMkyX+EcKclJ6h6VB15K7UIhVmg5KR4sZh2z
AIkQZ905EL+KUr9O1pi8D940nWziyA9I8Bw1wSGizraaQPOdLJqgD8H9ca/7hasj4MncKh71Jro6
+5xEO3+D1xjhjomxuJUQWO7G299mDmYocoZZ9uPNLNGQ7pTNX6dzoqFIjCjnOUx4J52AGnqCG8tl
t1WKSGG/OCyDqsmIQYz3SQNOAb2CdM+oWxGAvehqLhjrQ4yIQASpF2x0ymEAfzeTWJ6avpLEa83A
shDWumVy6zGeakAfRGPyV47pJRMBBAPgDH6V0rPHqp28tCzacKDFVQHezvdjHVqcpdHP6aXaHSPa
tQFC8XPr+a/Bq/YdBHaPsT9dcKGSXW2SsOQ8MUBS6aumEWOFwjnTbjhxrOkjPKAgWZ5P+H0tloM5
StPomKapoRj962vgoBv6KkENutyDI1hUP66GOOtS9wanyLK5cWZ788giu5WNmXOxSYwKJQx/9Hak
/NIUmmN1NU57QTdZBmsO/4g5QeGMo0oUp3hAKJE9DaUukb9zPpKYtm/cgf84fcwNFIylCXEVm6af
QWtLwptD4vaWiuT9Ip0tMV4A/8Jo+tJOLbAyadMM0xpwmrGq1hnRwDuDkqYkxwU+wgnweA5K5Tv3
yjeE3E+xmwWRg+cL7OFikafs/6SG+CjBOcY5dWzVSWQO7p4S2LQSgtIv818yc6wtx3WrLORBTQ3B
hjLU78RznPbu8nmOett1ITgdA58Wdhz9eoUMN+EsdMkIHWHdSmo43UHHTcRS/oGh7D+Gfqydw49O
eZOc7vSdh45B4geVkLMAULn8J1tac9hetTMUR6rRwWiqIsZsZK0uKbyZPkWjM+czIHU5LHatS6ol
ZmwJYBcjabbHWGgfBwTokCViWs4vqayr5DYSoM2Ho43R8zkA3oMDyqCsOU57DfOx8JmPRiqbqDq3
9wt1WjXqM8edlANoA8Y7tmjbUyMWhq92lc9Yx4E+KNGLMWT61HMKvFtQALZb+3FeKviR4Y1Dhbmc
Jomh/SjyqOGp4jzaqiC9mqmQi0MJ6CAx5k40l5fdDNyh0nmODzw52RUN4ZaI8/AVmxu2SbJCsSB6
TBKNbbeQJ76lzw366uHnqhfF/3D/cqY6mX9nJeMTIe0aZIms4S0IO1g0vpFpnN1QIIewO+xk8D9E
NhQ15O3yGxuwcPnIfIBrAIY4IipUR8UvUxGL/0F5BcYIPYXbGUJqPwYy0CA7kXaAXhJvXBzBtMvy
EJLvO7OULyExUcORfheCaXdTttBxNYXtuamYfvgn8sKF9mAEHgGf3cn41jnLoeLhNiwRNjGAZYg4
JpBQogwzi/hDlHRDfiGKV3Ha40RfjVLkd/3+dgxQZOTM4FRsBQ9gnTmyiLbDhmlwKMreb0rh7q8W
Qb1U0osLi4f21P2a17ukUXaFelnnafX96d17aGYY9IN2plqTTPbuncanKkixCJSvBUaiqo2iVu2I
XGeJkZC/02iH0ePAIvRfn3lsTETKcTM9l4vD6G8N/7JLdLsoZG+gkIfGMs+Ov+M/gWkuCLQx8oNy
DcYxUtgs7JVM5J9i1Fqa32U0JJh+xjFpCR+7Yb06kODHXk2NWD8iZagDjr/0RwUPhxvJTG23JiHP
uoktult41iT6hvDUT/oxD9fkz2KHSz3iJH+lsfSy3m/IPWsAJKAlo6NcxQz6E7IUiHMTGUB+5uVo
xKvZkzPYH3lra0Tvo7o0uySDn6YhG9xvO4b1x3jsY2Cm3K0R97CA2R04UHy7Ur9iJt5vSHYnRLVU
3OMXMxjVvkvWfqEZbr0Vg/n2/Pde3LcbrNleM3VL3KGdPf1O0y+MPdmPnt5ESrpnX6KZhakd2GDG
A1NxkzX3QSwNJHOZC2jT+0rSYWzC1wxpvhPXQXgqGRJDh4ZPLwmGrZ+9Upx2rXGdxZEWzsFXA371
/S6MlJ+gCt9SZ4OFlgrgDrxDE3jMqwwjQn9IyS9GYc106AMKUdnq8mN8KfgVfEapt5uhpCwucM7w
dIcjwV1vzwxpgSDH+2XfQHnKtxW3KDY7l/Le0rL79yZygAf+M5zoycMJW+vNzCh2cPuI5WpTz9Hn
92msB3VSrZAbcbG2vMVs7z3NjdAdEcM806270C72LLbnUUKNw2ktUP4D4hoexUkUG9ga5NRn8WuU
wyj0kfTM/196zvV9VvJ4ZCiIKDXGSPjRfOM+7CdPwXOQa+HFh3z5dNICR43eP66h7wK4fnkFpC5Z
QG1Z4KRM66l0F+Z6GMAnmm+2Icc6o5nxqglKvZPg93bFqMTe2OJG3HekoSdWbfwOi8fzvm8dg/Ij
MxQsv5z3FmzDw8a9AZMaTVACdt821Xl4gTA2FMKtIPyvkzvCnwLqkYjffF27JkdaLsJp35YzQjD8
Ddm0rA80ULCrHsjhMmgZyyL61tvxIWBalyaoUIDlqxv/lH/dmRf1Ott46049qe0XmHJbtul2KNQk
E4ssQfhHFPjqIug0dASY+jOvdBH5i2gO4kfa1o9ymmiYRKlyVOggjV3Lyt5IDmMrAuQ5iOAarhHs
Ad9Ce5YX51a+SA97oABbTyrfFx5jrcX4Pbm41OCptOPQfQBDpK3JbgljYGK+egxu4fFF/o0AhHbL
8qzcg1K7PUaaOdtzaQu8Yd3IC0DMelFlYGy9IgqAS+UElNrMV4ImmPcjRfL3pcAwXoHJdhcUHvRA
p95gspsiIhgESRxvSq/iliqfC1VGUPY9rEMZaNTRGTu0uGswZBqztNk+tnqEkOh29KNjc8mkn9BL
KPWQJNHI63+UA4O2ALa11eW4HahBAcw0yxddIZhin2iPYqhefY//FZWCnT1qReTbdNlIS01l7uO4
lJN9lED/AC8UlMyEdPcIJS/n8YV5eZlQ52zGPikClvVsgrEQLI9zfI/HvC+LsKGWnQGCOIgAqWns
yl71qRjJ4Bc1caM6UgDAy/A71pHI0riEFk76PV6yNGtZ03uyUQQcEgtMDg9KUYHLlL/81eMPdKSa
lCFY6FUhHgyfHJRUENno6TVL1DCqgJDw3bNf7P4x2KkkZCZsQ+t8fO/rlp9DFnuBoBtK35++UPID
PyVZ1ZfV+n7uIWgPTGRW/ZLgDziNdtweWx7Sj6ub6jSwrW5hmUf83ckpz9KKptdGtZG3fb3b63mh
PUxu9qCiFgJH/15XqsZDkgZ01396b5Y0VUEfoOYMsslMZ5Y+KRUZf/K9qjZmvzdcVlSSL2BUYOxW
hIZLZkFXJuMQ2mWV26JyKdmljatL+gKZR+Px/mzwYCejuXfW8l6+rq0BYZKi8GoraE3LQrytKcX2
0/TNomUAa0y5DLD67oKiHnuCh6dw9YVzdSY1pkv9rcMn0MslOwilOK29sUi5/qao9a5MxIC4GBj7
HwslA+HxS5Uf2m84cE8rSrY3+hThd9B8o52pWsL3Y3Wt4vjPBHTIGM0YtZCNkkUBQ/MT+rU1j/QJ
262F6sn4Jzry/KqHPM34qYGt2rItSO0/dcJ0DXMjsjbw0LyuXJgTazgOTNttOT0j9ECqfq2FHSYi
gGen7w+GqiHdPFo1DfysUk/us40d3ubuE7/WFMTD9L1s4+9yblpohhuMZtZUX4Xe2wUT8ZbrKzwi
49Ja05QOMMsHRa/cnjU7k2ewNsTvr65x4dyGC0prr41xpWN+0LVJD89FOZCqu3ba+U0AbLksx8mn
g36Mg4Tb+IEhbC3tv/kaSegalFYqaK72I3FLug97/RV2rF7dLfJq3RBA93f5yLjLJqR9sF1m/bSI
C4D/bXdiQL/PomNXhB52B3BaVfZNe/Ds2tT1WLZwc1SBViKG4i3LrsufxaCKsHtuTdHa6p6gcvIM
Eni1FltdcN9FCT6DkBcwUfCkMOzjDNsj/P9WjlXYVAj9T/ZfwSjTZfBlHocxbJfREariJPWFMWVp
yDTH82L2FBO7+L66zV6TOIsCzK3uhBJRqCenFIgvFYa1x1nDirNO7aN9CndyNwGRPePj14yH1x8/
WkH9mbFtPhMD6v1iLTXLZXeZZjaYZ4a0U4DwSLermnXARQ6WBiCTkoEqttsQPuek2W5oNckhmKbH
8YBHhWHZ5NQTMMtO+OcmvHoyge3NCFvt2+COs4D3bdooAKwKc2qTpk+T5SjtO/03jfQwWXT6c6y1
pb4KtZzr4Sf/VB4vtLuItPObEhd+76MeD7tgpQwWhxqfzFTCcWio7CC1cWmj05zkgg0OqDFb/Aei
iB2binV6ybSmHmq8Kj8W3qlBBeC9lMamsgxz3QJQ7FSZa1pjSRqmbubKJI1LI2kzUHpO7GfQyc8O
kjJxWg1v9eGreEjjNfjHcJWEhN1T5S9/pjp4fXejQ+/Ad+qxpyylU5vHNHLXaANH9qfB4cgkvz7I
b70cHWEWlsc6QC+mGihe/uszr2xXXEI11928u71AjIug+AJzXatpWXloeuQLcp06jBFGumcgGGWa
/G/HyPDqu8u1NCE9idZb/2iOe4/SSeapY81OothPMlNaVgDFmSutoly1EzggPerYDWqSgvY4vNCY
RY7FVXZZN9Q4Z2ptd5/bUe/9nEX0Ypt3eGtOW1dZyg2ffCYes5le/4Yjn30NvEXGf2xoPBmYZmJY
RehXemnZDmCBpRseDh4THlcy+krB0bOHSZ6/IbX6VbWpJwP3ihpBsZhKp7r9oZeQKKQJOW6Eh3bn
WsDN45wW8A1xSWfg+R1hpK8son3OVUdavFR4kN+Lupx8i8PMbTBUaH6mZcrmAcq7kGFzXSmkibzt
sQFBe0xwvNOU1egPzPzHe9JmX6OGL4gPXUTah7YutH5Q4vqA+uzk9A3dTIvgTONlDOLj7LmkSylX
yn0noFjTPVKNiG1+579mZC2CCmQllXbVXXXcEzAf79bISrNO+ZtbNQ1obBkGYVYCFP3sr5A1Lb6/
C5l7p7tIPYqhmQuR11VBuZ/NaPZotr0/TsSYz+gRBka31eKikvhRtb/mSH5a8louo+IR9sMdZ4sm
PQ+q6fKVcZanT5If318niX4PDDu3Cp1JrngkoRcnrhcdaf7bDuGqsGpOWNurryKbjAiDUo21owLb
TMdRMiwMctEkYl4BnEYa1rYQPQqKeDFeE3ebAZrKfJtnHDad0rFRpL15TQcXTXcxzA7NvfuNnhZR
iEO8on9Odt5p0gqSy8X/mG9IEGvLI6LgMtEtMdXSrYoppoSj7VYL8zQLQcAgJZyg8j9QK6qh/Pa5
sOZHs/cuwOGl19vL9/pBEPKwIDlOdObbYkEaPtWzS2KXEd0E4zD9wpWUzNERE/GFojYUiz7a6vkG
SZEVHKYCI5uXEuMkV22Eu12fzQyQ1pPV2EmkWxRtd/5C1IqSpKOlFrhQB/0TZgkJ/7oPoaz8rfTK
TmqZ+pmqZXKux+lc1dyD5kY+02I2kZU4RtzgKxoKieBYnAmec1ngiW6WiChJcLooUVLxrIvzY3/9
pueSgaCSXfjy8JqcPBywjtvmZ8AyswjBIT7sROm4fcXa9q1aZsUYVEHBM6Xhdp65cLUSwg8KdWqn
32Ux2tLwC2qR3fIflYE5yhhWyiksMFrz1eQbSBYxwToCk6NMaCTiL82Fc3NaihxdU4x4aWtUq2XY
NByBgb6I8C4PEzcJD2g+5Onc6PAe8+1C6w2thJgWsTqTUDp70VfMQjCPEulK8oGpoPgFv6C+4sA5
jTlYWuKPdScrxseYOGne67ZLqLWHUMo0/ZIgeRtRD6yKNHQRHJdy+RMco4M59dYJWcRAVEaX8cXD
SXMRlaQIFbErCWz3r1fYmwJ2m2o+Z6mgJbezWkfZ+7MFthAY94BzxvTlmFP1qUQG5cHJRQ77h/rX
Qjj4+faWepub5r7D8vUuBOE6V5qnDw6KHEKgGyGdTKFlh9rg2Vr7Nf4P1zn/Pp2E4WF6vSXnR6X1
eyF7Cl9At1YsnR+VZ94JOTiwlfhZdP4aQ6bfZa+6PWAw64mKjZ9QXovVQRoHSiEprQwj9Y/UhLRF
6oWpUXm9T92cFCVML8QWuvwIJfeE1n/mkrpmXwCgh5KnumZOssTJg1ZEGqN2reEvnIBKQlNbfrpv
0WqeoDKzIj7g1XCUlxs/+ZXaA7lyF9ZDtQ4usY/hknzJAgJSFc9VQMx64rtK8hJiYpJ+KaEi88fu
evKsgSk/8zCVNFOj108g2RculjMek9ih9jLmz/gAMsj4TPJzqrDBAyvG/bQ6eHO6Rv9RTBGG8VWW
MuzNjD8cCUBGIC6u4h7KbfB/f3i0qhPTBjZK9txpKC/WbPWAzUXUrdC3Go1m/fnP2k9XYkP5sCI3
ZASMwKMns5rsbwAnYN/KlYAZY4XFi8ndXoIp0kWKBONgTJWbxwX/2IBiDH9lKSOTvy0cv+1zWkhR
8CrJqyqkoEbAq2LRezKevIsmnhW7XluA7cDlBLcdjP9C2UP6el46x2My52cnn4NzGCvU3qnoHWmK
xHuD+DRvKHwY7aSmeXOhBBJoKQ833jq4Su4z027U6vEZx7KnCMNR2osywUzGQyP6NqldEvZkOJwy
JT73ShAQu+3KRWKeLD5Rdjj5gQ4AJmUPe4Vntc2XnzwoyMnqh5qjf2Q2pSBYmP9S66Ku/0mmWG4H
86No67LAaF4JhVBWC85+1+WQpa0YDVVGvioGtrvcJNaGmLvivMN3jilhZ+DC9sx9WPMjkTAXIGou
10q95zFErn03nbOPZ6PL5Xk/8ySEMs36wGicXkp68unYq8W/M6lPItQZYY3iROgojcWcXt9EmBlX
p6ZnEoN696w8PJ0+vejnH9KF+wzikFJmiyMwcKrzM+k+0tOxJiiMD0wbPldNi79qBTnp46PHeFKB
HppoKQoDi6Iw3sXRrM4IxQO/+pWd9MmpMe3W6zjNXr5NBLRmnCg+QKfQ7FhipDFk/n2439fA+XZ6
jB+Yfp5rOwLDGTP81DDG7CHGjPvZBauPqxD9pB3BtR5pijm2nMMVN+2t7gRBCC5LDemr83dj0/BL
ul35t7s0eVFzjDMJ2i8OuGO8LhZ39CEU/9bGyrN5kWSIyHNpmO+5ImD+RJJNBj7yGM+5PdYUG5yu
l5m7BvyCsCcySHL2cvlAftKOitxCxRSxJeW1ZxYXIYtbm97GBIa/C1VXnPtuJVGURTotuzoPhUiH
QUNc7fJIuhG4XaaaKnacgpn7FgE9lY+7EULM9PYtAFU4eiqsXWSWIzP05yBBtEhJItyIJs0rK8TQ
+kPenq+ZY7xWSySE7/Q8T276RAlCpueqfWhmZVYMqSDjETfcMSSLf4UKTaRM3XDeYGZvmBBsyYUL
JnrkAjR8fSHG35Gst2VIRDVLTSFVBIHCTV/57cY26l7imoaRBWOlx/iA7VbiqeibjT1Yxn9PFCWs
T7VJE/r/kkMf/ft8Sjnm5CQShBXD67FnHVvBD/miRz1bQOjOnzfmOK2d+ujptEKuTqYEA8hNPfWm
GkJxBouUqIHQipteZ/GTwb3j15SyacPUO8Rrr0RAkl0ZpEq+Qfd8Wvl3XNmL/u0dkJUXoMu6+26i
FEf8Rj5cuPJ7PnAFEe+yJ0Hkj+hrCQ/oSGiDos1ivGhZ2Ue3Sq6kU/LOalM2nVGU6eKc3ngr1iJT
2FE52KspWqB/0hHrn9qaIVGFpIoM3VTk7yNJ+TnCVo86bXPs6hHBxFx7fsaqrqmQBrBMyIjkxj0+
zgZDevya1gxZIk7B+rVT/TuKDSurNn3AhNlc1cH2rJt4RduH2Sea6dnHLCqCbOC+YW1/Y+kFiC0W
fauIQuPdZMxyyEWt/ERVduOwa1cWjuMMWbE6qfPZXnOY6QGXNxFn3w/C+cfObSX/z2r1lS4DzW3G
e9dxR8/4KlKlyqKnBEaHTXOJ5NDm9tS6YlnD3+LLAuldQicLH+0SW7E4uAxyOX60RcWQlcGjgVs3
MTuudwbeyhndE++0SBHlEbWZRv3Rh5wxgv1rMMMM9Cq2XQeAhetk8ttP4XrrmXvpTMOUfX4GGFIh
UBKFbc8p2iwwipTcAi37S/KQIMJba4CDaXx4TIX3KASpMp7bo+RTlNoeRFMGzbxHdupp7pTV4fl2
gukxcxWcYYraHaZOXSOyT4w5UxjXx6+oh78mBs0L4gJ80aEI9EhEG5QE3URsHxhEDZ25vEgpLDpG
zsfj9/Ap5PDXCgmHgAPmUIqhxJ8PDSWQVwF1zChBzPaF6zKPwAn1WJq0OWroY14zPKTgntxK6G/h
/lp2qwU+mWcxUkgV4M3yjCjXSSUPDBwAZcAVq7/pcogVzbAZgeM9+Nz54t/fjbGIxxH/jV+5hyoi
dqGfBPy/A3c0+1klIPd/IsUCt6m8HcMnR/edTzlMfxMo4azDCvpbsvclzQJsHlRA1k7gCuFei2x9
dZR32lC4If96PuZY2s3hpUxWKU/CT/EfQpApxVi9hjIpOHKHdiUDDo2rrRrImLvsO/ZcYO/RiAWa
hu0u8134In0enLlkm+RrWJNwextxPFNVxNShiXoin1cGi8HjvXZ9Yy9IakYgicdG2RTBS9G07MFT
PWjjFBZ7HggHy67YURdnhOhcGfyCPuytRqXr/RLLXra2I+IlRIcXO+PqhY1Zz/vh/Gh7+EHQ9Pap
kt4PQ6meFm4SVMQ6sVkHm88Avv4UGEybvnNNfotOSyJGtr/J4LoqW/0kXAZvjBlK4MRolZi42JCo
aSyGybaRXJOMm6yI6Y/27gB6SAKlutN16/zaed7w26N5dBzL3ZEzwosr0D97d3o/pR4iHdXabPWM
gcfEYG72Shzau/cPsVGzjpE2Xi+1xQ7QjSynWjiGjPaYWLtIY7dIQXnagP0iXfQRvHf/AQqyr9WO
fVvb7UJbPGbzXNvkWJDwHViISxQhgiPDmva7ZaVJwrwJVSK8uI4gJijHbfW32JkKob5UX13zp2k6
CXhA2Ya0nDx95k/jAqVOixciUAEt+qn4W4tCrKPCqxmFd5Aw5HPdD+yt22/MVkk7BFuhMlhzlUJA
6fGhLMtax29/Ylh0B8CBJK8i1Ryy7v0Jud8zk/KlbGs4LrZKeRIvN8HEpgOIEBULSNePHju0TWaf
kp7PzsGXgjH/cMGFWCG4Kxo4m6NLw7Mmcp71y5jx0PJ2ILJA0yQUIzfZmNTD6V/duxz6nv1U2SR/
q2MtzfazlopQnoqTaQXyIlaym/GoeSToC9U4mCCFR83Wo3P3icHHufNXvhbff8M+Of7dQ6oDpsAl
bQ97GlJDDamgWQwmu+BnVrBQBpBLmkylyU/rL2PgPYBwVTY4l81Pf9xbKKDJ2eYWuVFM9FXGYEIW
5/npf25XhMlL0f1i1rW/z+s2qq8JWgWuW5wvlqpuFhVB62C6gqYgYsvIa/cVv7CR/B+BWl//xsyS
QUBUhelGeEK8Om7bYCQ6LKFAfRBN4FHYkfGQt7DVBFkroU1+osEFDT+0VTAPdwKXc/xlcdPiBnZ1
oPYQLO0TtBJUl7vwNRqahRifBNz7zZL3gxyrYZX1Z0s2rkhPkaNVxX+cQ+6E28kREIA0TnBZETtu
UJPOlii1u0xYCNIXCfHnOkBWgw/xNIJbjGn880JGqu5lxoqjgHkWn/DZHiePOtH/E2j3rYL2bylv
MId6qSVjLBM7Mv4Bfpqu1pXROFxqiKgflu3dxHy1y12qGWBB/NtuTBPhx/Uq0kiCs6wfSQtuoOyy
l4KdkfxREWdxDdrTDyzZ3o44CeFXHSgZGBqdbs1Jg2vxJmjZaDn/+C/6eoQEYl/5ZkrHAY8qi32q
oqZ6rv2q2fAeKr1qcf65seN9Tg3VXjRRCypha+szYsRGPd7PQrL08WskrXmhiIsUNeU8BKCmgzRr
tl3XxFBLe5JJ292ZI8hie/uQIHfhX8FAawQu+NSiEH+5Qpkv+NY3GFr7twMtOwjkFKpIGgfAuCui
f2QMUMB6zE2g7t79mPtkTy70bu2TZBN2bpJWrvZL5s53nfUW/ttqrxVqLc6Dn2GaI291mWsAyVWe
zuaro+ftGG5eT3IsIOxlb/5z7CNejr3dOnyJwqWMw1XSCUCH+X54ktKOO6JdPVOTs8YDqCSF858D
ZAczDlFz5/fFFcn9Cp9PPw6WEa8+5PJ4SbqtFSST4+3AYcs7DbNmIYeP4iNAj315wICed4ZSUQX6
gk15fVDQlhmi+XimTLdvWTW6TbShYyfzseY6DMaAaov56YM515y+zAdBngM6mpxPWmRg2VzrXurF
VQ6mpXNLde1q0Ssyl+KP6tHR30bsO7WdOM9xxbetmTReR1z77GAAwS0ZoPMJBm8T9hQ8sDDraag+
M/ybQkxTGXSv3mHwf2r2jyLStyA7L3QVl3Jcw7iMD9WCmtOQeh9oAqGalEGg3g8yr8Pzwh1Qi7sE
QoWAQ4yr9KFl7mljj9q4F/hrOROznOdyo2oq803KGzn/1jv+En235FkiXW6I8+REUjVUofuRwedi
vCe8/KnlCJ/R7qehTZ53rmHNcD04n67lmxpMIJRh6jkHSKQ4sMxjOyH/0YFqwuxVvnDYqVTYjkye
NTSXMuc7cX+6p99VxvTXyNH3GGr1KcFVhfDi+PR5uFzlkuV+dbiF96dISsKFIq0mrOM4PBpxLpfY
fcps5asMITW+v1qsinzYY68LTqZN91yh3uegyKRB7t7q8iY9hKN+h2x4df4ec2E6mbM11OmUwqUi
WV1aPy0peNvMr0hlj/zjet2wt60KsrPtVBJchgsdW5PyahK2TGuxv4Z32j7Z0xkwcuDs1llMthCn
PNq5aZ2ExPa+wsztl1n7EJ38QLHZxOyNRPFVRLjF+lkkfcJNGc+iuUyWfA3oi7R/1HxhYjTkXp2c
vRzZDGYwQpqDT1zbaGXbEga7iZMxmdoIIgUBglYtEToJhAvJMTeAt0BOE7KdLJshABPI8ylrj6lX
BCJJs8hb2KKkRVNZMlyNrICxnVb6bbb38QK7ZPxr+CYdDWFe7WDet25T2jOZiklwl/hv8cmpVnbT
mfMxeM8+MplwWNAPCw4HfdvUL9sCxzQlJ+a3yQHxkZHlBXUNtr19Y1hSSYOEWl8jg0YgAFgOoSkD
bB1rg3NvtcuAPfIkKgiK3pnSDAU+v9CFHy/+aD0Fl5pXfWVR1lodvMQ+XIwmDwe3yY08r9RjjMas
ufJ61lLyD81cJUE6uCrttKAsEXGRCexNbdEjx7ys1f6+iBN4EzVGo47VaVRS+UeB3jX833FDjoJL
YdRtFEkup2jMs5nV1whe2xxjQ/v0jjBE3XVxiZfazNgEmsioqXi/kfzV4DXwGansDGvp3g8vLqHG
IzNWe7feTDtsKcJiP2b7engCvf1UnYBy5ekro3xnTgxDhr/EX5SRT1KgwkZEZOT/5hvRYCnbwFLM
kKFwA/C1iibieiJu9Q6AIN2uDBCdNGx+dkaxv3jaxt1P4McjJ81xYMR19Er7irNQiVMMWhvUKxWl
cAHPRP8dpzDZoJTOB1YECd692yF2qnVWVJoB2ZZczcz6yDywIJTJt5NIju49yxw2o+UYadcjZ6P9
XcWoybd5sggb92TpestRJFk5lVpqxGKZ7CZS5gcfruDbdR0vJ5gYmQjUd5l58cwEvGApxRL2t1dq
Qq7SIIXj/y0ME8hoYl5hnbxdDqy+WOUfJSv6FtXBTfyE3gYn1WPfprFeQWhN6WWP0WmnM9QeVQDj
gxvScozuFp9Df08l2FZGMdd1LKUa6cvuVhe95BVEj5/JQiC06aXZu2jE3DHYT0rdMuPmej81o3uR
+BkIOCm+5o+1GRJy3I0Jeyp3Fbu62gDd7ex8Utzj/8P0jlfVywFc3Ar3qaXvM2qjh7haRsvz6UOl
gpCdCQrQbk3w9ib07jy6HNkAYVolUP448Pcf6aMIi8MIXTA9BmVtJymX0BJbm261fDz9uf2DO2EJ
FsECvEi+s1Tw9PK6L2BtKV7DxpJqXMvk+buO/EzTVzPlEyHHwziGIVLbsLKHEFbZhNI/xmcir+eN
+zUfn1PB2ZHiV4nauv4SytCVqYzp2WJ2TWqd9HFZha50ic9DNYf3HLGjb98kgbcfsR+OC9ZpklcE
t4bqP4KWh+E2ntisxofHjE01GLoMzU4/Uxb4XD26VUG6uhqBOOEkfQp28JxPkniOM7rydJ3MjFCO
u9O+ZsF6T3Xa6TckvALXTm6fTH/MgYiftQx56W6j9VfyEamsg5P+/mYNxZdHOUzU9PDm5u671clr
16TFZXl4moeATzjpfz+4z4uOjWVLzXnvYr6ZaC6i0TJJrbIJwXDw+DmK4Wy08RyHn0Wfzqz0UaDJ
0am0jLbNwT710T0X+/roJTRufpiUDg1gZQxZgpi6l6vw9B4MOAsrrWnl4U4mvPNQge6G4xsWMvG2
g8yDD3QU4A8NqhBGH4801qJne4oTiipJlVE4RmEaQlYXYuz4FOBw0PUTqkys+yv+uSh85gjMXeAH
lGd6hxTpz+ZS3t38oDrc2Wze1QNwuyeZSXrYUPubfo+3KLc4hzUpSUSPX3bfCumFGqovUuNi1zbU
UaT/j9tjAoGJZyrc6B3YldLFAj8gYdVGxYE7s4MV7DJGNcM60/UTZJWB9hRx7fb1j06wRtrG1RN/
6re64vbb9StAEEZo5Oo7n1r41eMHGFJLf02wZ0jL9uae0ytWh7f/ebyHzU7ErbTb1RhTgTd6cTeT
W3sHkZbjtBxAvk+yhN25Md00QxUBVdFnE7FK+eP8JXWN4Rmp9r5OhU1KLUP6yfKMBBlcwWsHlULa
9YjsGes+7e1TDcTKsIdiMXakpdSU17uZNDG6qQaX/1L/C4cu2UP+GHik1i7QJQ1itgRnNZUwPeKm
123+fV+1fXyxbkuKRRfBSi60LYmJ8pq1N6K7fIeeonzMaTCDpRUEEV2JVSmaguQ5RA+5SvnjZf8E
78R3wi0Grhk9+3h4HH1JLQ2v3TwVa94dzCpzZCfOZl6shtVtVB0xibqHEVMDxfmnEArtnv5q8ypL
u3QAc8S4LP2MmOpgq3iGJFC4PzRsdrDyGCIzd1JjGlwH7LZVdTitXBs+KQDYFDSOqpvVdyL0Qh9v
025bW7Ypq1kQepszjnQHNxEr91PuFRbjdBA7kn97pfirlS5sNetOUrKBagRswjxI+4wJe/IoGc8W
s70G2tNulZmJ4E0XUy92NtWtAubrMMIj4iSKRec9jMG36WAkCVIPUDre6QDRE+nJb/E9H9UXlNB2
0s6mlKP0qGIEbDg0lvp4J9CuJF7zcyQTA6E42Pjxd+sF/lEy6+n5ywNo8Emdrkym9OI2x7oOh728
67D1vSrO6Ts4m1BZAft4rQ1ij4Vzg7RHmFL4x5qCG6e3r20K/QR3Us1KKi5qsTttx+xvEwc1/jz/
uWyDJdvelJW4fDxcle9pd/fs8mOAWmaOPQokWxwITTi2csRDneBOlguac/OXyheeOtNv4qfwyFsA
QFcrAwQnvg7MuBKv8xxtPudmMtdnQBPUrey1rDeXWy+urDW6yQJYNTNQZEArWbLNuGPCsSvHvf/n
ckRBNCNwrQt44tdnPwNlNw6g+5q3F4re63+gZydBOE+Sg8eN+ugKqFMy579GvqZ0Ti4SYwyaFEuu
jTrrPZ1zRwl5tKMLmvkzFVcBvbsbr+RBRCfLIhkJJUPXyuq0qD7vkbne++7DCxK15wslDxcpIewO
j4ik7qx6HgA5iK4p+0/Y1Az4WmqmB9gMcMzjtaDP+FojDR2iCtT+MOMsLpEI1xagGom87ER4+ZA3
9zr13FeJGxoSFLsfavM8luwKXZCrxiiM8INfB3qWLV/ct4msjSazlE18Ra42TypkdRL7cO3a35QT
UCCnEAXEGF1gF6jBB9q7fvrvlvvrioF0zzZSU8+Zx1tCC69DWIySJRvCk9Eo5KIVGbKmKCEn/1/C
Oaex0frjIc/TWX+ewabAyijDvYCkWeaS1ZEE8qbfA27JKk6aHkqbmGSE7+vv3vHN9by1MM39M0Qz
7QMDrmXFdsZqYpzhLTl9oPBcYpyElafPSpC+0NL8nBL/kBhEz3THeuWNJqtfL6KfjKzJUGMVJqmA
wi/8vvlMxE7VMhnPCrEibk76/qcNQ8uFvy5ohesndBTB4X0u/L3pdS2DHa60vFEmGuNEC9SoHPk6
2Rk5dNq2FOCLAG2n/Ca0BAxZ+mB5Kx4GBL1RSFqrUeS5ORJoHkpEQekjti1Ek36aZrfeESM7bcTL
K//HGNj4gW0M2dGuqNZDUXAMat6KuQ4V95iLWjedIuUam0bkqvAqjIoEF+yGzWVMpCAQjDzBrPL6
vWAQKfcxpLqPLwFbe4VjmjbnANQSqMksEKFxAaxySQjEvV34A7zZMq93CNMBJofyN8dhK7daGoC9
j+IjprFms2CJgxcBT5EhF2PQkcRQAIVj7PdGaf3NvtTYyubmzqt9oFWelZCGWkUrvNPXqdRLMTmC
CYjq+uz7wwY+336RgCG2wUR9a+8+1IVipPYjXu0fvd7d5+bJyNZL43fjxHwJm1WO9QOJI9na2JuD
zjGn8MUItJZo/l69kqk72l6dCKTBo2ajelYyqoZ9ptf07WBQ/+cHwwSfjeaTt+LiOTGU9si280Bs
lAW3ry1M+cIlDtM6875wMOKmx0GkqVwkiFQHJ5qDatslfxZWvR26qOTm2L2Whw7TmyIQCuT5EXoW
uGWYvy51glwQ6oS2z7LKcxK3EfHjt51nI4SvSBkO+RqM0e5DtRGjGo6tiGNvRTuWnQ3FBEixNty/
sskwnVMuBKBK7EEKjD4xccZbZTs6LEEtCjBfUg8Se5DXxVAn6Bk3gf7arawVhRWCAy/XUYIApzLO
eBSbmJnBgtwY0tk8XBddDDjG2dPwLBbDorSIkK2gWnG+1pN7/yCjM+4XgADSgGtNFMbqIT22dHHS
e1tuP+oyOBTxX7fp4g4M0KmlzKCD5OjH8jI4xL75vBw9gi5K0hVStSDaX1rNsPdJqfnM3dyNf51O
za4qmDrHCzspFTQWaqhKbXIGpYyqn2n4RCkXTkwZCroWDq3uSO/nss7UtIbvjhTAfygjcA/xii06
RQt40sA0F/2ueoB7+JnuORnZvN2QZqJWSCehBjlqTQm1Imu7hko3eAYQaFuK74yhyZABjo/iN+Ge
y/g26hKCz7wJbPSHmQsLmxJm82omIZ1PrOGeIE3y+oDewqGnm7jM9EvQJ2ujWzy/5tV3BkemNm0y
rGr7LUL2ExcQJAuT4IZozlzwKHeI/ISZPSS//jiPma+vqcPuHWNWIB9APLBA0o/oKPeJDUwPlE0Q
ALtDpEa6piTFFlo4BEBQXlb8gtWmJkoO8d1rSFz/BhrZYrpxRzB3rvs0r/Jx3Jp6bY8aolX2oMq4
FWADMfhcwL9ZuyK7ZHnB3RBTGx4vFhIj8y84AE2uneaeSI6IFw0LHjlcbEeZa/PDUmBGmN4qErNL
mJBXuk2ZaF2cQr7MtfOxxzpwcIMP3+14WNkztyAbkxX70DAP/yyJmLE3on4bqRQ7Ls3n80BrCsxS
QvyNPOUka9HNSaMuIMA1ETwy1v19bGrAGsPY8gQyjJFHFevfVm3K53koAeklAgWBj/kSGrvyfu9k
shwWlduHI2QggCWogXlrIak1TsamxAP/1CYA2ELDHCoJeeVO9dFH+aBiUDf7eHUUxTy+wwMIjnAE
HJtyBCeR0p8OceqFv/oA6pHI6dC3OEHa5jZm5TYRP5vEkiTQ+Sr6dqyXYn2z8XOhSJuMiMpGZue/
HP0gEn6zeSo/IA8vRRRoAxbDavVC36Pqet2VRv8j5JNE/yu81pTYRU2mwYrUULQe30fuizycuKl4
SsluypfSsOdH1Yu+zrkfReedfiPBF4WawGKnwQGz2E1lsfiqASJgAg8nLxuwdiiavBamBz8AQQFu
JmpEhE6PmtIgbbtN/OvLLkQTps6GBTK+JLSUqQk7yffzbfT3bS8s4oUno+ITvE1BXIBrE69EBEI2
f/oNOnzgsI708J4OIl7r84aw02Q0TM/5B1s8YFkI4LBv1Au7bDC454k7IZZmxVeO2qmacQ1xddbM
QLvk2iAY6H9hni6gCn8CLWwOXQT8o0pqAjwlk76HW2j0cT0Gai6uvZeN5asiqNtMVOhSN8SMkl5s
JTFGXhgPQj+EB6KN8k3RhU+42wMtgTw71TQMZBfmQ1C5qIqrSQNh4q1MMN1kKxBFLE/WPAxdXIeN
nZNPqnEQRULD3NuZUmHrTWRjZjCcP1gxivAqazLTyJx/dX6Z3ap4OwyGZKqHGYm3cGe2xfG27f3J
2zgNsksXwM3ZLE0+KN/XQ4wdNAod4MjbEqynuxwsG+4RqanPqH4XmcEAcKNfMvXkL4nW2oFnWBTi
P17o/GaE9Vwqh2rWRBMulGj0MMEVckcwRRn6nuti8VkcCmOa1OCZlnDxqGgq/+6tHFcgRB2R1T3c
M+Z4rBqNB+6PEL2fKuCpse+0dz2u4mEvZ7w0ShKm9W3uoI15fxK9kHd9XrvJ14DK13DYMpt2bUqJ
/YCv3u4qY2fn9bURV+ZGMuV9UzLq8/o1qGIPH+0xZUCOWsrvUS6UqakJv0owF3IuUUEJwUGpLX3A
VfwTd1AzZae+Y2VWAE6rVcdsH2hph5fSjkQ8PoPnqn2Gmbh8jQu6YBrmg3QiZAudEVf54cenYkTq
nsBMovdnVy3A2EjYaKVnK6BH3XbSXZmAsLZV5VxJWlHvSYvWpFbpxNbOtXbXWbeiVux3AYJrPAj0
UWiQKmKjYGZqEbR5dWEpAefSyzapJGkaEf5OniKbKOT66g5a5wQn94zVUzu4XvWAxJA76dAztHos
ykrUoZzba6D1m7X2HNTAUzYXBJyviAhSEP4+elgHRlewMGIRysrHPq9jRc+jtjAqAQn6i7rEstU+
QkM3ZPbTmGpHVF8gWafyFLP/eU/WL6iVrarRSOVHDe50ZbfOY5qXxZyb+gFrqVRj2+17pUKYNhRv
SuF6dqC2PwT6SXMBqCPY/GcnUxyQtp9aXCXo58aLC/jQHfr8sQM5PHkEZiZP6T2AYnHkbiGwDNxm
cS/FQ6E5KLfGGnmE+Dm5UmVOySYxeiaKJ9t9xvgv0wjJq/hingW/vir9Y4AwAG0wUbvNcTrSTh0T
1qr7UrgrXKt9m4fVMFl5PxYH3MwaFg5P1jtv1zQAh38wPnsrxeMhMQBanNjeimokjCpdQQZkeDN/
jRBay3Hdk64o9/e0Patosf3YcxPdiKcFBFXR99Vg1JOPekrCxD3Ey60wOj4IscUBUcIJDJNy5HA1
Zl6AL5029oQOjQsOgoiOKdK2HQObDlNEMeHxsiZG5iUuW5zabjzM/aR6xj1smNFjrCck4LoWm5er
F8plHMD2cEczfvBF8OeUSNdrn9l4rm9FUaeZkyDGN+cG6KXne63rlRu8KlyK22/YCVsgSFgVTnJn
ywFhkVBAXDvqASwylSrAanZFu0TbH7SwMZHFET0glNxe19rM+2ImHCb90zTnp5gTEETQ4NKi9ndE
AlNvEQai0Vchic7aB+giJYsxlKy2qUqz4lAmh8+sR9AaIbmVjm32F7SjrxtKNsJvFKIdz4/MH1tS
DAT1YXHCbDJtzd8PQiEGUIf4wOyLWOnTUAb8KMAH3xjhCfzBUWXIxrCbext49NvcVmo2TwECXiDn
bZ74OhutkZllk8I3FcWiDEw1+j66IjP/G2sZ/s/+rZHg+UAvoxiZ35IbosV+/ZzzChATGs4CAWGg
/863t7HMnK2ju/uBIagbIsS+hADe5SmulhYwamT9p0q63A12b3aH4dVTZOurnXI/T0EFAlovmujH
7VTWXEcfaN+hcyDLdwuuwlIdGhr6qnf/lg2L5hO0C7cxw6wJxD2aZOr/jUjRsi+sfFKzbkswHNsz
pSEZ+d/Yd2iVBpBtn1FAnzpvDP5SOJHW4SfPuvBs27fMxgBk2GJ6aDsTWngIECnnN9PHsDNbVZdU
25r3VCQ2VQ3bHaO+g2ZVSm22/z4x1bMZ2WvnxzfZPP4+74DQWK9cOk6y9JCZE/Cb8jS8J60rsqjW
LjgwOccP+u1zga4dBbAQ9T38NIoEgFyuw1fw/ySsGIc86qU6Kxb4Xp8trYV1lgXuFlVuIT9LvoXR
Vf/aprQBPxwOY1hIz6lVC65DOFhj2Bm37rVSz4bK5QPezjxT/6u5aNNkf0shKGpVIiEHdAu9T7r8
4GzNoBMULvxfh2ibnhTd0UObAk2iHzHWb0GWpvoL5KPHb9hqRngXzoTEVr9AJp9CLozivdxNIrDC
V57Gw4wWA8RI1DZ1MqdeT3ikOk4BdMuRQppksHChiYlPcA2ML697Wk/cVxrlq4uF4FxEqs8m51/A
wlSs0uFWCilS0jt2CNHsS2lmyHb1Kjui9fMHOt0itzv0iOoSKuCCRBMbrud0CvO/REhoK8WLqfIN
N3NIh9Egv0G6QIg8uBcxHevGmMSadM+cMVOgTl/fzwUJnOIJnGaXictgl+3pRC99FsCg/pEwYsL4
VG1tZbJ99g7WcsX4K6eK65rQmYvvTkcuEPuUHJuLc7eq+UpGzcS4IJyRWWKXlALmugkIq/fI7DD3
JQdOQaQzjjh//zKL8eBrOeXBRytF3db7lc2373r6tGJT+oWr8WgPsIVMIcP7yTxL1oBrn4JC+anm
qLwOLwliFB/Aru/m+CgKBMu/AbfwERpEHvHa2meRF3LxoCX/FxHs1yasDN/TTnWNFnBcL14UAibW
IpTwQpfWMNjwhMPCXm1lgl5hP6hcFlcoWe40+XigH7gnpzMSOgyVxxclTMtP/ZJ0GBZikD2JHSVk
eBGFgUMcC6L44uBtFbxkKcXgXOKiOidBHDX9F0DgMFsbDKvhFCUgIZ5xzAlztyk/x61VCX30IyyA
PjsPQy4zvcwUjJ3ljiXi9bBsD/c/QpqAD61t+Rz+d8xxYVZ+eg8Iifyrl30fy0T3l0GJ4d8VdeLJ
t4GiUTok1RyrXezKou0D+Ni/OYMRASi/CQ8aDTp6EO7p6NCI5Ogvev1R9T52I8BeP3l6D8oMdKPh
A/s8j6EtA6P+3mzGxktxDx020mOZp/pJK+30apgOHJk95l1toP0M8s1uHnvfGkbiJ/Ht8NEOJYCy
o/PiU2ix1blTirp7jfVhHnCgoy8kfdDOKIBWsDrLc0pmibA6wHz8Ll06WqoOSRZHuXLF6kmeRP85
UkW83QxZpDpaAvtuhG3J4iRSHehJnn73KFue+o5ooQawCbE/8OZQefY8TQ090ujoCRLG+jZgZlqT
7fSvnGAY3PtX6Vocfyib/sYWtHulpI3CbBpJn9QlxnxXBJiQiT7Y+z3v2WvqpRc12ymN7waD8RyN
+E3O06haFpyeaZ3I38XgPtfrBqI3fD2pVcwEauYMwXVsN4UW7GuKnB7jBTT0fmvsWCyHoVhbSnr1
1FoDipxWaLbtSlSRiKxJpeu1aJyHD53WhojjvZWCJWi5p87TcTOdIyP8qWYA9pmG94cqIsTpdER+
Am0dkU2WIaR0wz6kY1RFjjdDlKldNR+3yvCKgvwthN9IJ2Hxl2gHTIjTdwFRLedHEqefiXB/c2KV
aHQZ8yGeK3xGXwB+09gqqJxKnuDk+fL3CB1XjvSMwfvipZYlHUdM3A7Qhc/bWGySUJDumYwSAJQn
s5PHt0gZ++e5az7VW0UhLt84SzlniOPv3mjxFQAcZK+2/I4PS2hckoFpazYSQHpzcDpd0xeJExUX
YDpBIZDmIBkdwn63NwaPYgdCynBiy49Y5CJQHlyn/sP7PGwJWXrJlIbUl5Vj9wmPtrBXGLqKgYjG
JAozP3tJysiAOtm65zfqb3d8aejd55dSKvLQE+RjdugLUnmcdzV+RjocQN7AN/yP6CBULLeb/Lc/
M/tCqZ8rRNLo7No1gjDV/t1eEQ8lY3c5HbvBZ6D7uMeWmPcfI83FDjrWh7CxpnlrqZI/ub00eb0O
zh2/7eSwW0ZPSmcKrhrCStSTFO4aRE/h36xyyGu6PY/hdlCnKNqFm2J5tl17jMe44JfwmsqS0dZf
8WCiUQ7ls4tI55xc3V3pjp8F1qc2Ej6CN0ZkUHi0y/Yui2jDmYtanWn1WQya0R/01jyz5FXohNry
1Ol9P8piN5JXaIsFCQu0q+UeHuOE/WETZj4c3eMgoBEITphpAPY5ZRBzQvzM22K+Pm78ZS7F2V5m
gf9mgxuPhYbRQrBOWFKw2clE8ywrwvQE8E3tK5SgjKdGU09mNeFasjfYnNbSQs3IHxfAQzeZa7fn
NZLCBB8U/mLVf3+WTypJJMYzMWzgPTEg5fIWNWYdcW/aTLG2Smcrowyl7pxrPKotSwcaErXK2/q6
/0IZRlRaEkUHvP1B6cVeMLf5QOJu0JDdS589J1CvyWVhlFZnFVFrrhnSYGLLSEw7tp9ciYvCJ+iD
CuIRHLE6nDXLiK44Hc/Oeh3eOLhBgUbvs/2waC8U19uRrtI95H1O+5D8Im1K27+Oc+FpITpv6KDt
wiLkE2TaVAv7mAL1kWVcgaxExo27L7ehHASq8NYbkQp7x/PW1qWcx7RxsU+Zw4i+k95dcey4LsVx
8v102bwiD139m179tp0HfFQzgCpK3Qc0FAlKfCCCgXCjGDnRn0oKFKmEfhfLg+droWogXsHsykSF
eQi9v7ZpivPlzPp12n3bHbSvO5zUHbL4rRP8bq2V82PTtS8Qp86po/afQk0qGRoeGLtjYXS38WJZ
2KEKn7WlA6uFqZOQfHt5hM+AUI1O+UYFQnmjSoEgPI2y6rmmqXebCO5oF0x3Taga3b/WhHtOsOJv
EpnmcqQKMXOixEPCuKrR/k+JSF8RdfqpiNgS1d8HOBAsi9TF8SV37QKMR8miZEVyXuvwKH7wjuMS
fTV8Dtg0R5tyFtLvSuEk0OJ5pH9p/k9LMFmGuKqsQmY3V1Ew6/NPYwcJKp4oWOqcROo0p3t/4Z8I
wFqjZC2l0+dVFuNktfZDfBKJazP5L3K3zE0FTB1E0CddQPHcbXtFfZgMUmnC06cwHnfCW0Him7iP
2/n/ZlLvN7SZE2n/WaL3KMrRYfLvl5BP/usyYN3C249I+8nBxqwqAonryEYqmh4AOTNrVj6fo7Ov
OnwwetrK1A+wXHxaax7fu1N8aNrxQ7IrH2WJYTKICefmbD5mEsljrmDp7xfLN2LL5Boui+BhxtdB
3dlm9Sp1BXaZY+6MBbbOcMxCtdUrFaQgOkS5nS+wfwiSPtuOGRk6tKAXMDKp8qbE/SSVqa33vNnG
zkglx90B4+RA1jW/8x4mi0lUk/WIfpRJ6hZHW8Nt6gbKTMNopLauxhLcP7gT8EmGb5LEBUTAIXer
dy++J/I/SI25XnXmnHTrHCUbI67Qt1QrmmLY9MBbuHIf0ocfoyKQeRN2c3BY3X2hE4COrF18ExgE
xR5w6CMgfbBk2ujfOo5njvdNDkcQ/yZDK8oQjopDudvrnGrgb2738+TnZ2rziBsvbm6/c5fHapFd
XPYCFNKAyYLGPuZ9a7PE6cWIDHB0wT/nhs3pGx+y7xQOcttsIUP7WUBVCUqZWKfZp/nauQqHjHEa
+8BizdaTo9bR6l2tYKzl5b88Fq3WahS04MWWE5cMMJVrWY6u6hvSuRz0IIPlJoLapm3bNJoL5gKB
THHfg68GQ56zcwkGaXo3/V5YMqulR9MwhoDJP51092/WMdwhzMdf1vmgv001wl4zJ/h1lFIjXalK
577nJsdDZjl9oqv1q3xi6N7T6jjN9MKedHA+mn7q/7MTMRAvnzkmgcYKzZqBMpmH3rjC0xKJEKe2
BO4uvlIvCyKLO9Z6v4E53z7Atnfs3+QDBHdpYtB7QwUlJD6d5P7iVismBG0dxJiQ4/a7TsorZQI3
tBNBvJBY7V3Bu7JwY1IKaYLSrKGhf21nsUaWmkCzIq7ipHCeR1sC/rxM/GffpYgTU+G2De3GTTaa
g3LsZHIjFcWJnHeMSJKSzygSFXI3o8N2XvIbnNNWxOoRRV5KEt7Q
`pragma protect end_protected
