`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37360)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCTcg9EscIq6lRv0lzTzbJavMUVh86XJUllIERmp7hUgdDKmDoiP4tLWT
vWHecVa+UCDOmOlYTpE3u9dfhToKLfZ7HGZd70AYv6iXF0wpaZg68nhtzSuhrqK01yWhaK3UUkU9
tYA4qB+mf4UG14CJAUX08JotBO5/1hX0PRBDj5WceDJs4BkHgBhK5UdoKj8Kx5RMZ8edmmuaxDFs
/sUq1uUMxhQ5kXwb9Kwf4f9Sz2RN9O3rbY87eHo/S/ktDWZrAWQJcxFD/lytgNPoZzUXlMFzVyCk
FEUQ0+OTjESH/djd5sQ/XUwKtydKj/386fsQWiu89cPRxQ3i+LU8sbiqcSJjC8QJAdVlqc+fAECX
dnzDDAohle2GJxlvguhqDpb5TqXKqy9z5Dg38WaOwnlTMZsDJ5m12NN2GhL7RdHMlADc8uAV8k5F
AeVOGW3TAfOKEq/Yo0ZOXujnFK4uwUTctclWh7jE6lWmadroNq2uj/iHm9ZX35FzVmQW1JMtI1uv
8tf8l+4JayiZa8cul0g8PYSOXl2zuzEZq59C9SPwW2EhDrqz4K9uQQiBT9GCARpGx/1tseACg8zg
ylfrGN1ak+irwOAKRXooyCwdKCBAxLqx0HAW6eiAmQJbXfXU1ykNu5p+DB2UN93h0flgciqS6LfT
6Y0qqiD/oaJPYVkgw4G9MrF95w1UEBprLfPP5U7uGIb4TWfGjKFNtT6ceJ/lt3uOM96CJ86rPHOc
Vb7EVXWIJ5KyVDt0wmCOrJ49PnmCq2xXOXJvdXAn3BcRM2Iy5XmxAXDiwDHfZUvK6+/Vp68DuHQB
VyIY/DqzMgGAi0EI2W7bmGDAqdLiWoN3kVI59mKOClMh+d+PlROB8TP51EaetCv+8SHzgjnot0yZ
hreSRM8IF7er99rOyemqGoYStuUXR8JR7IBcOiwT7iTj0yvqP5rhCOLm5LAamWGKtn3UtKPu+th1
5BeFq0+vqAiHpldxdKXH+4Zkk+PbnBetF392x71dB86lqqXGBZ39Rq6z06uE9UQKBvvfdYXdWo1h
QVE+33NK679TDvpH2Q3dQ5LPXYRV5dNrTD7iwyBBAM11ZBA9BzMugo0PM1EZkxFFmWMxm+Gp7Atx
QgkXKwaLXEsslH6cffHNVo55yr/uCZiLNlaY5uufg9MHo75FQ6a/WhPYMLQ+2pISGjeKaE28Gh0h
DLE/FElPp/dlinarRAL+s65YgYCFBdlKT7sLHX3F3Ae9Vyp3HsJErH9rXIfb/wATlRchsSPuKEeJ
OIsZZznxUlvDVa1n2agbBoLQghmf45NBJUkUGjnP4vSEX6xRnw3tVHFhJAGrD9R1PvQ8LeN0AquF
WLatpngTfNIkXflbooNYkHYelI+kXUGYDJ5lSrK0bHt4BoE992aIb4AFcqL0EVtW02gjxYQpQ033
+I0MO30hF2tA9n2hRKJMSuymWK94EUkW36QCBQ5FOtER1RIQH1tJKNZijk5WcpFNQngKE3Hxj5N1
dX5fSP37Uoy7yYZrUT3dKAUCmvHNGsIBEkKKBTCA6OaOf46SvIB3bH3HfQn3KdDUamuy62dRHq4a
Kv2jyzm0RzJyIIkpCrEm7vvN9U//lCkRTtM7aM4xeSzIzNFyczlxZhqYeD02MGdfRdMrOZBOzBbI
AGNWhKpTvtjH6xLEShfZRmuVXpvDLfn4FUfFFNr68ssVGSt61LB77y2DrVMgq9baGq5XvLpjSI5O
Fi4fKgAah9psSwyTP/CLNVGsQZj441n6sXP8HFbM0M8DzLcuesJ10GBsLug82KXUxRxlvxIqnIrk
++eDE3oMi8pHSxZlEDzd00Sigfh+aYK9CerK8KF3d/5tQyuBkARZ6CKHNhbh/kBS5pRdYUknyYaz
faGCg0p+isLm21GpViXKlsQZeIBx2RRMcMM16k1jXaZLPJToxfDA1PGoWilaNMTQtgRdKVNuNaSJ
yF1G7T+g56yBRg8uqhAOznib5kYLkcMMqiTHgAuFEHWduMPxa+2IcJQg/Bbb7oYYtdFcSoRfj7Sq
Ri9jH/JmA0RPftXy7nabLuUIAwn2G9mF91mNveti+yqG9bne0oXJCWiijQ52kgSbry0bTjwmmB/Y
oWyHTGolC4dSWWcZyNUcKS5c+uItdNYXh26zJaNa010XnjKFI/GV6Co+0a92iCBt1XtLVF2WKJEG
p3xfJY18TlO+ZK60mLetPlKvjEfCsnflio8epcgGtoqB99mUSDjoNixNTTH60GJnkSbFlkWWdv8T
Bf6UkKHfTR4uA3mtxvbYv+A+pYMdktlA6Z+AJGUt7nM1mE5NGnj6N8RXCkdhm2WokKswrgJVI6am
y/8Uyw0KnlJkr3pdJa/aP63agXg+nt6vZfP6V/dUYOYRMFkyyRYpgdR4aVDrHYyz8Jc517qUyZjU
aMTHpQV4hZ7FkVUMaiG7JKoLYnYciBOP5oY8Emn91s18i/KKSttG5qap+7jE7evrBbkzI3xqyVoV
OHLhjU7uYSmadHP426Kwnaeh/nnl4BAzujoYvjg92BH2yQY+uI7ih68YhZEvxpHZvHTSq6u6fo3/
IUgHUCcCvuR0Fv1s3NlXDVFqkX3m34KHaKW8F7HWaZ4HOY3H/ry9jioBoXXFAF6ZCWS2IAMvT4/e
pZpAt8ngiHF7Lhh9UrTrvXuH81PeiODHrlRS5UeEP+8aH1Wytxe1ceNboIB3CPHI0xiKAUalt7qW
dPNn3EctnzT47tHtyvapx+3E6HNLsgn+1If4WTrTC2/ZvgKPX2ivBZKkme50nIKwrWahMo6vfg3u
jMc8sd2yDwgEPuFiKqq29zJ57T9tbKqRz2AwcyYrH/7szCEBDpKZ8iG6yuiXwZBR3lCOe31d9MYt
k5EMvD1gSdTnO1qpPYhWDsg1fgZ+Cx3Ssga3qkKrvqKGNfhl9b7rHt5KDbSLqCgSXCc3yXHhuu+q
jGT5097MCC/xCT+kkQ/L3S6z8Gp3qTFxIV+9QZZhUsO9Mn7xZwpUAszCFwi2SrmnZ/7MZLTzgJ3M
bHXHFhOf0qRj7PfWrAk4/21hsGZsLA/FuqU3tKNY1S712jBemnI5+yMivv+7IeEi9cTWp3yISz+V
aJdHfjbf3QLKtlkRRSobcr3xyQglCfSaRsbidOt48K9wTtxQaM9AulQhKGYR8qqUh0qeS+6hHJpk
hYpMM5CgfjIpqMF/+fN5r68SeOj6JkLgx7kpuhB9M1lRdD9gAVwP8GguJD+ZFJ4MzjokbCMJ5ktk
2Qk1aS/45wKNvFBRP5snJELtX1KKeeKn+OmCJGnSufHVDAVlwcYIw9qMIM22hIE5cxcVsTwjAerg
49dNmann0aURucDHiF5XQE+7tp0+2gMJ301d/TzIFC8AG/ol1I5cZJTjaPgTkamklMFW6ZXxRJsU
OVkajPfOEvSi5XZM0kXCg8NVKcsugPR5qUzX2A7oQXD+2peXxwXwEnTvCZNiK6GPCZfi5VhLYqRs
PEKkVDGjeLA/kFsOwncx9t4BtLY2Fr16WO0x0lPnfm78phrz8M10cqIG16nvrlJio2rsWffa+52L
nYY5BRDVsLHOna7ZVOD+7SDUFWUHFBfWGcnetEvHIWtGIoLewnp9qVHU+6oTHrRyomvd+ymfw86r
9yaUhQVhe+yBk6icQCeTJ3xohzjicljucZ1BOebI8TMGbTvhogqowFlniiVBVD0CW08cd0YlVZx4
LmLDpIUIuLO7WZZPtYfWhzbQLsVbiqrILIRftSZcJGY8Esn2H9cY1MLwWkmfxgmC75h7Sq5Kcb0g
hL3KxAqMdei+N2zyqKUa+zGtBJXcJ3nSv2lYO6mbFrJMOVEAmN9B1m6Gp+DYRBaP+HoKv/Rg8R4Q
g9qVr0aVON77jpdYHGEAjPIlRAu7s4QXGLNYrLlQcNH94oRp3dFjI3MUzj9bo80wD2VmXn98wsuw
E0KAz4qnrPmMN385qyYcbCPX/0ZL0E0Jt0wpuUDz/nZY8DU7GBb1AY8EIolJumy4UXeCaWS6m10d
U6usxkfRH9N3Xb3O83sqDcsvTd19PhavFuvnyQ5rucx+13HdqZRLjCb0K6sHXau3sRsbK5rnKCA1
pVgZnR7F/N1U08JI4eJgLgIzHgfDIqSgPlQrCjPO2394okd6dJOw64+uouvG0QxTxgFux+o86G4Z
f4ejFdkfzVhl8RlMND0JHx6e+SYoWAOBL9cDDKUHYrZp/6g7+JZ1jfyeCiWzX9W9tC5C+IK7p1Vx
yqIM8n7UAPkKlcxAQBHT8FWy35By/Nnl0rSAvcNfGPJbsAvx69s2rkMx1amXKO7uSXe3YoD7Or6i
0ZEzUr9fMEOVwDyXwMLGuDztSnGtjJSC3kQiNoGyiE8Gc5utz3xYSKnLkG4ZRLTIkfj9XUBo5AyV
SeBzoD3WeYdXDvW36iPf9EtM8JF4TahX85Bi8rrWzkhvXiQN24hX8QnQyRIawV8LmaQTxqlX85ll
unWccz1LXmh+DEDsio7tTmDZOyuJaJ35rRnGzTmDVoI5ml8kH+7ou/fom6zbfxUY7FTMQx7DvD1r
qP31itlY3WZozwKKAntpTtT0tdBhHKV9l46p05zPvhNFV892uRMK213us4JP0q4J2kdoIAQrErGR
QJnvem7jz73NeZvJ2ShS+F6DB13bLYeHxnxyewjTClHqBrRrqcGlr9QiUbedXr5H/b4r94ThJjYV
PTYRT1/2wk4qms3LIRjnPLBXhppoqQTc/5P7Wuq4oVut2S3RC6qDaMPKnwl3KJGxhABvcY2I5PIp
AX7KSVg/C3JxpZEhraMP2aDosrP+iXPA0kgcaw2IS1FTbYZyvMZ+PBGhzwI4ZtR/sktlqJEwOGba
DYExCU4zsOm3DcJkUG6uu2AY7FxA1Pq7CJ26kC4/H036Bg0CXAl9k/aXu1NfpvoVevgZGSCdXROO
Z+RLp3uBrFlbgWGOJ4narnQPABj2d4xhzRw7ZVOepVh+vEk+/nzf9YvQOjczzXbB910Ettq7ONwC
GOc0yNK24+7urX5Mhm9x+itSBvqUK8MkyRY2ew02nh/SYk2Xy4PDufNT/RKQOO/gZj8DbEo69yzF
3iA5dXl0EE8Rpng8IbXw5JoLy3IKtcvyrY8OVVCg1FVQqSQ7roNS0M3cdLQLkz8UjjKVElxVI5I/
k/YaPqlOsuQpVkhKqZyoK6K+xDjJL0bzVmoLp2AQmMQx+MpAwWrYWjc382QMClX1eLFxxwnZ/xYh
XuoCdVzVyZW45a9O2NQ3fvSCr4UY8qeJKxk5kBD7dCMV2Twzi7RJIrVD1747/hRfglEPemjrCzV4
Bw1wdGVTwWww6DO2WdVvhEk/mfjxo7+UTbc/l74ZOHO4CLoBp4gZfCBLvgmD6UntC2PGFMx1WCEO
7EsDs5hkSX0TWrub/DPr+OKG0n/bJTK2OColzmF7vGl19SspPm+G2ugnqyeotz0wQnKcpjI5ylH3
qfT9z8agDInbuCE2QrIGh6OMdSneUpvDMEenURzcGabjhoKKKGd9nB+04hLQipcSopuTQxjBbFTz
f00DGrSYrHdj1iclqB+MK/Bbf222U/uOqndYcTei2ArkQ9o5vvuoku4T8Z2zvxZOja1CmQ8eXM25
zrrmdRFIDhFabSDcA4d5wj4F1giU8v554UBM7SqgN/rG9+VdUSw6SWgte/VBe/YwKKDMtuWK4ImM
EqAgk9yxBvl5397tydIl4mkqM8RHE/jsGQaCC+FBeEaAcVlQP617QhH87IUFBzYEDAfz3ySh0/bR
uaRRBn1XMd5S9ZK9kOxwmyfuBIcCjBls+H+xUOeOk6yjGhaBuN7q3AHP5v3jENH0EUxnjrQrNaX3
nH97tAeneWzo9ZSGuC1c6lviSWYXIdC9AF0yEDWYGqtoIuK21MJGrwn293CMZFzhtOvQhh3k4h98
Yvst/SFnDNN3dz8YgZgtVjbX8Fug6JibcMp6LdNQb2gVXY57mio9z/bwgTYMtY+fIanWMFQR/JA0
HhyV9MOkPcMGFWre63jg+25VMor13g36eOTSjTwLj2IA6IYIq+3Mr+SMlj24ACCQO6L06mXZ7Xnw
/kDgv05mUrru7xuQFnDpMzDvqm72JKFxwFcXa16dvNF0iwZUbXGgU1PcVSu7VlWGQEyvYVpBDiu1
yGbd6Ky06zdxNTLu78CiFrgNHrQQWZqohJ3Rkd5qkxsMOQLBXINUO9vPDKvL0vIatMJZxb1ywsOH
BeWQGPzjoODGxsWjk0eB/gy92Dc11G4Wu9CZaQNTH1jgwOS7kJIAYFIxJgZJx/TxPobY3mOuG+wo
/7ecpFEGdD8ZRYIVWDoEowRkdfvkvB+HZABn97z7dMLuNO7k9k5H9LbaPV08PtBz9sXS34spCBRI
nJtvUSqD8jMzi0R24djEG5X1lus8nJhT4ZExXwXZN1BY2hElHbx4n3WWBEMxpqxi90fLVsmmdvQw
kRxAyI5+J6KGE5RhDkLIfYYDFeQir0R457/QoVq8QIloeS4LtO/l8q7vNyAzuldxEiTAY6Obj23p
znaM1FECFDXkj772HZJuonzLDuGQhztDAOH8X07xZIvWEfPTqUnMPxCnk5BaduXk/V4ut7y94ilu
ghr60dkTa/IQH30S0L9je4plgfvLUmGaFUbSUD+P7poP839f/t1dGpn/ZUJi/h021llZJY2HAEnN
Ix7uNNYMFRrOK31ctOvDXlWAjl04EKtSGmVeU7P3Vpo3Pv03ssPzd1w7mOzWkkl6mpBl+/ZAgBbt
rtIVouFqSc+Tb1LaVz5+F6HH1jolDvduRpMigmqjCaC7PTu473dKKUTh2o5hhttdLaknY04dRUuK
vq+knaJBn4DhsqaupruRE93pXOrtIuomoOrlNapKMcHHxYMfQmRHclu0GkhZDviT233TVf7bn6cH
52fwyEEqF/aCaKmi61ihUA06EyOHXT/qEL4jzi/50nVNh0H+fgD7MMqIvdA/eeVAY4mW7CDaDAfa
LjffmX+96Vu9o6J1FRcs+cmyhw63z5kTag02FU1oMTuH2eiVZHNaHkg3huq4EolM2kY/1RRpndc5
dRiqTks8lyKkyYmIG0eMaPzGag7Fh268QbdGQNikstJNoQQW7wGemRrbrY/MI2lu0bGu8N6aMtiR
P2yiKW7EgMmmQDMhl3QymuNuXZ8VjWgV+nXR0o9QNwiZMDLxaAzoQVgcLN0e2ifxN/tDcW5oV2pH
5fcDNoPT9ngjFdpGS8Z6I3DhjcXWWFtI3tJ4qYQB+rU0i5awDEMBsLSmJ+GUWumY3QNaNgOV9LoM
ylZprrMLmHYkchxAKLYvKOcIryzx1KWzPWuQzjNyyU+fLtdRlU/fMxe9RGUQq2SQs/oFkzGDg7fg
1DGvI9jgxErhjG2uaFR9VzfeazRyzAHqW4BAXRhjKRwbS3nyRHDq6UoejOhulZFoIV4gNaMxtrl6
Ag0/X2uAFP2xoFn+xOIhtNn5LRUnpTm2kmImO5jLScbrleTZvHYSPB9txbftauHzyJnl70Sr1aEW
oV7Yrkq9rd/bQ9oBHbQ1PCFs/iBJkEcfWiMOSp6ZBOuilcjxkDvzUR6B9rej9D98q5FwAZ5C+HUB
1NyQsflJzq1J+goEPjXVuBcb1biRUoQ6StuEsZ6J6AMvn/b9wgu5ErxlezcU9AEf9YRLsRAEaaOt
gvSepA5EZXQIcU254n494VnX7af/jHbuILwxeuiYSUvxuEN6Q/Y4cvWNLf50xKmnQ4Ic981go4ee
a7fcsH96zii6gwnGzZaNZWpFiwrTG2EUT1+ssrxiHmI9AeKp/tuulCSWUWKSIHz3E6+13Y5RzuMU
JRaBSQCLlYqtQ/54vMjg84ir86jhE9TAx6A9tQi+8VBZBwlWKRV78ekL7HOQGEPkKdK5PfTYkCrD
m7Vg8uZcsnFLh21DklmrJRUGGBeVIo/pMN6/9nkbyS24Qfcu4tov/ZTXDW7xJQonHX7b8KliFa+N
1jbdJXMfCyM//Zb6/4Te/Vsu2JHeMT9qJFHfxPjq7J4h+J0TQuLNJgxSUB2NUr+xqQrE1ZdRm5CK
tCdnE0W2+Nxc4Sc6J7Z25mQ3Rd2wUiyEl7eSHRn70/JYM14HYp+ku9M6ulsWB97Xsl0dA9+HG2qZ
8dm+W3Zh0La+vphIYR4e3pESgrkFAQARY3iy+P4HYwYEml3/0cfC0wx2krAaVc716ImfXP/IMVJz
5wP25Dhg92tcS9NTQH/5/w6zm+Y9ZJGaQc8RXjJYgc4VR7YG+M/Ct3uLiTRJeAlM3MO4HnLxcxz7
sKLj1gaGZ/btDuS3r0T46A2UfnumBgVaQr17kONWsnwXOJHLduIJesArP4XMkpEjvEKvpbQwfFTE
Zw5xF24ASuLUMyPjOwChWB4Kyx2TgeGQn9Uc0L5tuzHY8Yg1OfMafAmRwY6ymD3HsgUvxHPnfXJR
RqV7Ldp2wJkN2mF8+QFR0o5aQJLzPtjd7VPUyzhYLS78UDbnQZ/9ik9TCvoo379NU58GRPJW8O+N
pcLHVcuQDU1jxg96kJhhAqRc3d70dHXbZYjXxlvrV+NITJkf4ST2eMEX5nO9Z5J9XmzKHp0OyzM0
ijgu5qYESMWfww9Poqa6Tu2sOz2T8HpXXfjHely+q3cramkABDNTRSkBgT3J3ApD3KV6bj25Nb0i
nXOEXH3Zya/kJXVKE2dYKQnZAagRBf74wcz2255PcrVQxL9oJSImBputn3dBCGIm27AK1ZszOP8w
xgrcPA6ppYDyT7xorABg/NQL5f+DJHEttr+Ckv4RAzMXkWyNeaePen1znPtoVPd+AS2l+RTojtx6
4XfO308o8hGew3cc9PkhSe/PIu9ke+5pGpktj4ioZgQK9fRqj359WLanpmZsIADxO/XyHE1pZ2MB
fOwH3LaCLoR4Yr8Zqia9AkAJv5+PYa5ZQZZzT68VAlJw01TnBuB+t8v0EiPpcB8GMOWDEt/tzWCM
PUV6PGAEwmjRyiKLfUzZT6P2EQ09IH4DiQYi4BEmDMOZFRyILouy/0TlmmftDSCPNgQCq/e2kVib
cOZ6PR5LgWmVy67IuTBz82zz6IJQ9huhKDkSsf38CaJ6SBkuE22AM9+HF47sHxJ4Kx/SUF6K3NXy
Ex/0jZLl03lJCYAwqhpbhs0OrPzIOl/P9RDLUsfQBI6BWviStahEbZA/0c15tsBK7C+Qfkt4Mitg
Z04RUk9RPYcsqUnjl800jpHFthg9/NNVjmHA1HOnLD9W3eVIuR4in9j8pk3XibdJ53yzT+wIGZQQ
J7JJNSSnPq3RY9CGSehXBalFTnFYna1OpY9ZkSwPiTqqHJ4sHRlB7SBSzg3/qBBIZfuwoAOP/PiV
Uqf543BAWEJsfDNjl3BemV2iiu+Z+kiI/D78Qre+ZdDPjAStSNEoLuJh/JABiy4SvAC9X4+9VHTK
C70ggKeANV29R4PbqfcrFpb1+fYZ+bfPKdOetmbUF4iejv3yAOQ1ZQaNX57Rmq1UD0vdFschOblY
2P/BPt2TEz8zeyDIQH1t4S4RI8rjuXSUv83Y4z0Fpzi6hhr2p2DA5eZ8O153rdeecrzotW0dKM0O
4nf1Ug0idaHrBtvfkPsMIhy2zU3kt1SSCfc6NbNUOEYtcvRDIpOkZi7KIS6lL6Xh0YE4RFU101fi
dIy+BA9NqXDuImFMZzhgBrJltNNCLDQ/oF6q6cpgX6GgAJ0DeL8Gzz6caPGDyI9Sb2fBe4n46cus
Di3Z+qdEIuSL9TnsAJUIm1TPtqW36kaUjBNXDmfMSJsDEJU8dr0R9fZVxkeO5uARf9V+xm8IVR52
Rk/aeaVTS1QC7/8mB7r/xKuIwx2kwhDasswUExiNU63iuQnBD6CIrD561OHSone/Q0FVo70mw7wH
XlSaCMJKeNU+pC1b+83S6OH5w32QHQW7MIwz1V/p3xrVKqw/w/rtN1w7Osvl2KP2TkBWltXs1BUQ
R0D4Ge7mzdclM2BYE9Tz+rCRr8Bz78Cq/C+imblEIt3fgokRZap2g0IryZ0kzAyXKmpWLzNSKPY8
HLvKryqCccAgm8u4y9RFGe1e8akSnzRp9vkRV9vHUVWiXugofmZZCU/osxM78//LCsg9yyZafQMz
UMhGc4wQlvmhEISt4bPXTzYwlT9Hp/AJd6rMvh/w6+vGmXAxHN9FgUsPW//cuMsit1ci1PiRVpzD
gVITUxEv5Q0LVW5yTxeC+HBYYodr+jZKi/+up2QSeq11vYtmXBnP5ESMxzn8+QXXpo6N+/YAZsKi
Tc+jjjoxn0gBjC58jMNb4kMbX5zSdOwOTkaLx5OolX88DXUlCsE3ykLNVNEmBkSl3SLk6sADBLjY
SRreeJqEnlDr3aenEZRMvQ+0zSdlDYjfbnJIXX8VmLEGemlegQPjb82ukFzmbXWjfUX35DM+vSYL
3ciG7i1rBGvJSW3kz/1dxOT88T0Vp1TU/kXU1VEIy5foSqJiMjQPkV+p4/YGw2FJ8RZGJN9JeILB
uKPkYzdtNjKcy+c4WFO6Ar7CJfxPTKOLNjgOKy1JjBgBHrLGQTcqVme/IQUiVSkEc/5Lhg5GVfGW
5Oezo+YWiR45WHBx7tCIYW/TXV7zl/sX6EJiVV+J7Qz9ujnxy/0ZQiRotNT2rqP8HhKHCxYE7L3o
HTzckx6xA2mFvKDgaexrrmbjWxOAkkDxvgjx/22LDFTZKnl0l7aNuhKNpb9TZZWpoVQgQ+aYGvEV
gJpEofz0W/gGXeYlJ2Kh1Tgg9/p/1i3uwQx26OI4RFa7IazBr2wlWPo0ukdouIlfuPjv+6Tu21WO
PgdZyyyt24T7ibNCUMGNnOR6umadtnOtMNxHptKFWet1QFSQwhFELC2qbNl0pQ9XEphMwJOtzWnb
U0Y/ls4szdQoQBwt4JhjLHk5JwS66fMzoU843/P0AWuXd/lqEM4SqB1eUUmsBm+01BmfB8Zqehvi
TsRH+QQ+zXbGWyvGY3/YPqLW3Nr4k9SHO6gd4aPmmUh88WqAv/oGuH+esvWob3E2yfH8NR+Np4g3
qjbT02IubMR/sZQjC9Lo9B8VgpoBbCxaumPrv6P0nRikGbwfIDvXQYwNNgekfnSVXo2BrQIWr6f7
EGXlj2fHgkMz1rht15Ljr/4SV+CZJOVOkgX5mlbHoBBcsczpJ0b9KLHNuY4oAjXnc/nVzRWa+n8S
g6VcYQnG4SbP7G19+bHPvTmLAfaFJZ1dwr9MM8J0y0TD83GxnwdCkK/fUMK1G34ZoVxSMck+DA4Y
xOh1pZuWqZQzNlLQCaD/BpaS7Meh17XPCJFRFfgNu0l7xPrBIgbV/Hb0SbY/BbyBUpgP0dXgIqYx
yhkr4ntx6RZFOSKcVtP7pX6JxLM34xl3pARTaqe4l6aJtgF46r+5OA8UYBB9vrY+jblct85DI+DR
sCEkwWxskpan6CQEt/P/EgIq+QDRQz+Z9ZJc0UCPeef4flM4h3Uksd+Last2G6BXZOCvBPAZXVsR
Qon+nuC1RkyTNBiPIwyXjTHEUg9EXHS+HGpXXx6c7ENc2EKDgJE0AR4tZbNU0bD7mjx4mFCm7+ur
zEawq/QWSwJ6ori/vTD3TCZ8sRQuDsILXql6lzJCJrmCvRMD8ymJguZvZlAKy6OgyBF25gbDxTnU
nZeLZVuTsaOxNaits8eGpy3+O6AZZHSR0O4RmJJ2C+zX5WqzhfM4Bm3WSveEgGTGhxTlaG+uP9Gg
EW9Ctp9qFs4FVBZw7a1vW353XtnVCB/ghcFAQeEsj+0gKCYBfZBq7nSQNSFOsYVjQmsE/BKrVakB
Oq4dlA5g86/xYGhVEaPnfJCBYi++Dgm8pLP8PsmEWkD4sU8ti+26w35W0TmEwv11mPmDF0rSf60K
E3t0oPg2rjyjlN+4j+pjAXVslaoXKu3J4lM1B4I7vZ39SydtbduPE+9CoiNl5QkC1NuYm2aJRoii
t2cq05e61hAqiXnEw9h+R8LgqWX62nd8ynjgbiR4rjBX/G/oCTpN7Na7vVi4LgBEVCQkdr8mCc2T
IGLIjJL5TX0B5E9P4EkIdSgB7+ejrgSA1OGKxy/yMvnzzynKCiBrxTrhnVU6ZQiwZbhzD5K71zWa
iFVYlXrYWA0RTk4694nNwLOygHlo8y+v/0UWBKsXKjX9U1UooAMxBP8Aa4UWIzWM4Q/+9BCMiNyV
EbbV0Nk4M0EP4nu+gesoGXip48+SPvLwvQBrRlvgNWsjPokP2r62iJgyChRrRdA08JR4D0sKo5na
gAvlTX5ZTa5peJHb16Cx2SWKEmf2HYYATvWU6X4YxsOGNCkiSegufoVbmqtUYVVCr7flWx8ADcUA
ihdWsnzjQj9xErTjMZomgoeI3oKRYAQE/rt5Ynrya4mtShcAysJFHsebjxCfbHvq0C3A//n721ak
xiIKOUvBKn7Ysm4aRlxSYZJkYwa3TQVTubLtdicvuoAxj4RiGbJHaa6NL6NXCrDARvrcphf0cYIB
GkinK5oG6+RRegYyzGIhdPe9f+l0zG11lFtAHZbwrv9hZ5BwDaUY2Ph4m9ef74YLPZL16BzMnfF6
EwOQvn8EJL10bzxRJ5ZLgObAtnXKJfnxRLEx1jXUGU2jwDJ42enUp6f4Gdf93UwwdDotDbMpnY4F
OIwSIIaiZjYSoaM6nvE4GjrDegcqV/zg/PRLX4ABOTOiIseZgalYNCYjwpfzV8U5PUyGlM1wsBcx
pMv/sw18uU37hoUO63aX/TZBa/xQPuWiSNgEcxkxhkj+lvfxxB+OC7113lpivcdMbr4bq43vMJZg
oBgTUHRAxrUf5rAhzvrDhNh0DYCvU3ntfO/pPT7MYrsXnMC/yXnlhYNnvp3x1VXInxffcuItX/Tk
0b4tyZkjb0NAdNTTiEFKI1gj9q8aHOFroGsLHwLVY9FsV5F3Tm2uPWmelxzZsUZI1QGjSn/0gpSV
NZ9nbHN7n2EdVksIIF5Gryaw/QDlFjk0cs9XEH7+DnGfZCMd0h6yXfKCr201sYc9vrxB9zpN+Mu1
0tJELvW54pBr8HT4MzAQdB1+A5dpPbWfpb9OpgvbsjB5ZmX1J6ldchNnFKxKZlDBdxm1yFs/Wmsk
rSXF+ZByDPgbyEfFF2xCkuMYNznD2k5zpwBAw7zxxfEMAA2Gp7YolEP+9TcVM+jQWA5ZA7APPWhX
XKbwnjQS7LZKOHsLIV76al9Gk5mmvy09Ea+8OkhHTmCsMGRIvk5ciRaZwSaG31XazFzp1fihWWb8
76s6F1nlUJPBJf/E1uXbC71Ze7cIultvjQh7V2v2ChGmrJCE5/D1/zYZKVBx61YYvFir6Q3Q5qm5
Ei/hNfuTWyH7xl8/7UfG0MPpEF5/WBEEOnaPgKUCjYOwCo99hVXFvE93aG9ohCP2RODCzwACWNZ+
JEXTwiaRCdo4rJe6jJMeXblSJo2ZZ2DDMouTI2SCzUyn6CgZye82eBmsfoXmYA198V/D0Z6QC8B+
fgQufgJml4fP0lp952PLOG1KQx899TA/dYDIsEx/Hw5eY5dmNdxNePAjHPQIkKQNWUKc3c2OeKBh
t8gXjk2vyFmPko29RlWV0mJtsYVMeLFD4MU0FsEMtYG+WNj9tgsiP9bGTWFC00NuE5DmUEmkf8Kc
MvxQ1G5xLJhgZlvXnA/0ShVj7wdqT1OJ5gA+aLlR5RBJjM6iEuCgu6O3pi2QyhJ6nWVxtwSt2OnE
JCz5unPx6jme0blXgaVsty05u9o6TQP0h2/x9teK/50bAgV9rMdenAo/GtecJUAe8AsUxXq52vZ4
avbTpAUZ2BhRql5fp1dZMIHlCJvkPmIPXelo0cQ5/NPcWTWAZ+WrBnksuyKE5eHbrYzAc4jwS4Q+
rtUahOi43aQIEt/uAlqCN3y5+JTmwnpo9kJ10HAorqlsVEWfEd/+tBfLVJ0s5kb/59UxR92alzsk
33WNclkmnbHZKOQoJ6JR9WEvQRvYQK3PqpEie3gvzkVJg1K9th8SCM5VgbG2oaz+b8+zsVpU5GVp
URqXaOJKYXRwYkCeuZSnGXfItMFFq4dZM40s5ieUdsB/w5oshetxOceJxtvnr+fQLRXqOW05O1nb
OSjpZMcsY5mQkLl2lz1Z0fK7iQLG/L3r6d/pBbwmM8jHlHazOVeUOcRgCE0I6G9Cu/gEpp3q6Jf6
ALR6+t4QG66rs/LZeN2J/gc8w50PhNzgVRq2Q9KdcIIF9vT1xdwan4o/CL5aDPHUIs8ne7JPNTZ7
t1t1R+B4I9RlczD4lBfcfytvGC0Vf2LSR1LZp9iFnv8mHRbcIncX8y6+Jauzuk8JNYlfJ8PEgw2s
kS4XZPvIYG4eeRLJPU/E/L/THfWYHO3/ZcknkT0mKjAg3hzh4e5iQStgPiHw/Y6iwNkjiI1+0+JE
8XvDhaf5t8Cq+KMUz9PD2SCj2Jbxatzn6pbrjoWld9zjp64DTnBoAcCwtcNAaUS9riNlYf44LPGe
kTl1DC6Aj7tImMgexcGH0qohozOvdyfH2ZVKf0cOxHvec38/P27zzhAK8BWI5LqKiaagXelSFxmB
fTYVACv2nTYsKdCiN5GwNaPPpTYYlWwualmla259W9cPa544djdsWU4nFssNX/IZhdJZBI71KHUn
WO8VwstfFLtpQqXRKI8tLIxK12mUvQhNLsMLHGDNAmXzn8OOwyiXaHB4a7zOCize9xN/rAYaJXiG
UHvhBSXM0AKR/flCeXAZc3r/hzhgZEUKJeg+5T0j2u46kJfc5i24tDf6yaxPMJNDLa/wT91wL6e/
SOeyfUDv3yAqgH2lwO6gfUqPoMx8co/i6urXQtnBa5Z458u8O14s24fRwjwRtCbCBXhsJx/ssHLd
RUcjrIyhaOrE26LogTzad2UOx9vvrpVp+VlVkghq7jViZZHacTwCn0NjivrU8jGVsSv7vYLNBd7Z
8sjU61Ci+N80bFBN73bcLOawGgpy7e33Z84KvTfT14KKU6BacWJzGHJToNjsW7GP2rTAiyuAWfgq
z+oalZ5nQYRZjWsIfrKK5QCFjH84r2Mv8NxaiwcGMDssXt4CDCCVmI0BQgyszY5NWxpJmOLTySzx
nWSQL4a2n0OVLx0r8549dt65j4LGTRYUlVNYHCbki6d910NiRO79lJIADpoU44QpmIaXGeFk5xhF
N6TRoT9z/DVEq7H4KRaSeTKgJAchCkTKDJYjBpGNg9EQJrO2phABa/grBKyb2e+VOxCujmyIHNvn
dSCvQQM+52az+ZT4mP02mGAxyN8FjVmBH+iO3F3d/f1aaLjFMIvaxHmXh/qCx8THUAE3Z7ZbocjF
afej6OD4PdF1+5o+Q2585ssI5pfOgVS2J9DYDVuc393A+XzzKaPtZ0o6rbCo1IQjDtoccMzaO8XY
imfQabWeb6aAnfp9+E0Jvi56O3nX3XIYgr33yzHE2rkeLNsXNheztxI+02ZPzWOcVGf0kiTPFcSH
JT7b2REiotdEFcW8zLmNZMBqbFFF+busNbGep+GXjkpHPQRFAdm8pIh5KXZYCrV3U6kpeyG7MMyU
o7de9FVk4AWnxG2nusE10jpXRedn/01ZbYNIFRF0mOFCA833Sjh971HnYBDil8Fd/V+ktCMTDQAM
SrqWATy/udxxaKtMsqKLcyg2cTNcj0hkpUOT1R3TeZOXJdwhzlqQHCYos76kqnjBY3Top7l0Etjg
5RVq9v4HndrgNPBCRwQ6FO85vAiLJmG0haGGqhSXvD79SzBkGRxxd8r767euFrUUP7hM08oi95F5
VKBD9w6dfVjOWFoTSlZ+mphbN2joT4tpiz3JvkYjGEa+NogyVTQZGrjcyDO4nPFnmdGYovmyoO9Y
4Tl6AU9Ee0SJKJhJwGHGS6lqBiYO/twZOUe+OaeZvuE5ZX1/9l6pSo9u95fY7ovMIw5IEgIfxuVB
cv8/N7WvLzqHqclJXrJtNR1cqPsI/UfbOyLll8x9avxcEJ7G4FZV6QhNMGlr2+4r+tDS8AKsk25p
G1IcPvCujSo/Wr7WpHsD+3+/Rz2XTosbVHlJVVm9YCEOH5Kg7ajVj5r3aE9ENLzWVZL/5Cou/3vZ
Ivn2wMMfddHsu5HULMFA37ECpb4Eb3y7CwPH1eZb6/hMV8TtKG77WLnfnqy8pJ8R3mXH9DX0M2fe
RxMaV/shlzu3kzqBH5MMvgAjEKXW83lS+p/4LbuH4X+hAURZ86uXqhsmam9bRLkMrJ/SGGfkpoaV
KM/kRVCDjzJ+x00Y4mvlXEj/60+dwWalPDHLLlt0aDEkRus/bxoiwmIJciHCroTNnyoFRLS4p4Za
3f1vM9mN1cyETSVMj+jEeUKZBxJh4GhPar4Yvf9K/Gvv14+JQsQvzwu6pKX/76fMvKR66pkRXhWR
ahVQfTQy7ZfgqGYjNcS13iRrgEmHJ4VGKs67xu95drG5UtAl1cgvc7/7DwwNyAVhJxzOa5ffeNvT
bsgIkk+/QlOwPruWhaFwhG6NLaRe1A60EVnT87DxIFpwpKrgh6SCtilbh1mUg3HzHGVbBNYXHRhm
cmPeD8peFYpjpouEJzHf2KtLPxcAVI2sU13OW0fHO1oUSIFoHYB9gcD9nGKCFtz6aFs3zFu19+Gw
Mp4l3pBtUMh5NIKTj6cRwwlRrHhAgAsyb2z2zE8BpbJ12ahpHwJV/ZoMAY4MVgH9bacZn7PmczgZ
zOsi5bFNHOcCNU5OaoxuPum4k2g7OwoTwwDX1gKSyrcGcR1V4Ep0sV2plU6MNG+bAIt1hK0a/dr7
Y+3SRqLpF0STEQNs8mWynVqHOjHI9hlMkV1JncU0GVTmMhgBDugY9LoTm/hrMuSASDJooPs06XxY
D4zCS5DfzlnDEpMw0kt9MfET/9AfweoBrbiJvZ1zf1ab1rVJnejxaSUX5gw9sWdJKP9+N8vW4FPr
tV2CmN+3M30FtE3dqnn76KplYBBWBT1l31m5yVCsZ2xI7yR4hg+0DIuFAod5xgVMR+p/uRUA+2GB
g+8z6k69d9vzmyQE+RJqjs4n+e70KPYHX/VSNjOppb2O9jPWYJ47uTnRzx5OHIpFDwQWBUZbDcqA
8rjJ0/125Dnm5AzK854BjpomjqtOx1pUjpE44w0VnIMhRcU5HDojVIxA5zctYiGzvn4pbWJ/+Tik
XXF6rWAYaLyrHkxYoCeTMV66KjVJFgfRPfXST+6utBGUn8UGXDbDaI9jonDviVsts1NBeHYQ/zGd
Zsw22dMP+vi9d9mbUT7H0nr4nfEwhVL4+nk63yDsz9hg2gBtxM4HHBbsoR+XVnB/ZODwgxKPA3eS
BAl9lkI/rff0lhdoBGjgHftdjXG70QnaRCQLJN4/SAyLSUq8ZxNiYKDw6ePvGNC085/jf0QG2yVB
HuJIsVF4lOrJLMLjY9s7OXLexOq+yYJMf6OCXlNQ/N69Nvkh3xA/kSriTS79SxXjtq+X+tJol7M7
J0CbyE/WukzR37qgMlKP++3nc5Hkybq9WG8s1cWjD/q/fdCmlwJ8w5jj0EovPL+8C1sjn5tI4abd
PwWq6fazMrPxBBAkbolVoWHYmpwzSd0eNDxp+b60+0Q3H1jmAkLzJyhSzKYRoFjRf5bt/sCNqC05
0QOGBfVGVvyFNySSefPMag5cpigc2q3tt11+2nuCmETUItQXjQVyKrcqedbdiPtsQtHohdxrt7hx
IJ/nshanD/0C7en6fEejveF/pyWf5iyo6VxE6I7TUPVLrt7ziMJ83REhoTrWN76yOgWz/5+3AGig
jfjBBRKGaHM4fhg7H1W0Swfo1IZRrIxbglE4j6aBgPWlX3AbZLJexfvDAlSlrazwQWbIv6L4cK+R
Vs80rOkSafHEhOwo5kAVEkiKaFa9K73NvNRe+/yJNpmoCd+l67b+xc/++ZXXhVtS1qIoCUpDQFZZ
ScFpZbI9T3sVBEbf/W9vtTCs3txKxHJSCL4SPxa1UP3h7O7p1t267/dxmt0qL+kGPh1n/ExOkj18
lDzGF/ucsTnGDjc2HH1ZUc4acW7gl8aP9QQLtF7n/+o8acmXuszvCJ8QUFGaicjMbXBPfhhV1yXL
4IjuiqfAuski2PIw7Gxxbnuu4DrOP/GtOVRqQnEwdj6R/tk4vRQURP++0urpcF6sGw8gpuQDixTC
4rgvhen8jrhHw54cq2KuKPEgUfvi9McXb1bBuL7q/KSN/aCl/tj6Qv7h1gU1cRDM/EXq9RnSs8SS
l2dlFAKIgUdvc2qpqN5A85lUVjAmxUe9JvTKhCZmTbG5p7pTUKSG8W43hv5vnt6c3IZo/in2wzAh
q4ivLYoBOz8Qjx9c7Zy9vPMYWAHNs/q1RBopysuBn7i6PpyKjbCF6TyXKZd/tH2yipkuk6ImP1eF
s/LP9AG5wAuJH9Tbz3USr55pmHZqyjMvlKMIKQyVeRBQuX2QA6d16Z5BxvNDE7n3lJ6HNkHM7YiI
UIyDZMZwn+gk3fyr0iWXVGOt+jeaG1++hTdn97UglsDZ9KqgQf+9+lwV9r2Zw9kSmU+raTEQAPzA
nOYqI4rhP+o1jh2vqp3pyOCnlRkhSghqqNIwuOt7upR94qHpvEtdqHpKM9lFvrDNUkuYdwP5vdk3
vr32XtGcF75l0lTH042uo4MMcOqeCy5K7FWKOQZwqQ+EdHUPmYcnyr8BhjS8Rgp8iQ2Wr5cBsyQ9
k72a+sZTkGaHUVeYfx3hwvtu/z3VOMcwW62/sh7Pb7q6etTYxtEP6HNsDtwPy6EJhNHO2Jp5qaz1
58ylVBtU948V61q3iTujg6CE0l/X4iCBouQKfRB5w8rQO3PR3nierviHohdjEPIINwPEe7/Ol52w
ltno/Uxo7bA8jxwmpDaWf2S4aqg+H9NQyefYB8yIMN5FxrS2h/4/NjsRIGxUd1wOSJxN1rBcyovo
TPUe8vIDrRUCWEp4gs3r3MN8Vhm2puyaqFEzCdVI9W7pPm/3OrlBXhuMst7cEsNC8MVJRRO9y1rc
TccR12gwvQY5EBa09mxacjniVrx8FBpCJmfvQZm25CzaPKoCRsiCfGFzuC+TJ2GY3fPb6HNVd8Eg
ivrj7qnBgd+EcZU1+v5J7iOV6nDb5JLW71jVAapiK/9p4mCWKPfy9KlBpJ3PkR72CmYoOUcrGHlt
qvL/PqliTA7oZ3di9wmVH1CIUXK06OwnXN+FHKNfHicmuD0XemqNF1CZPv4ZfxpgWkFhUockMbPz
dycgVD/ieVGY+MhJKJJblZpU33CrKHiCc2qJGnqmRsc4fehjToBKU7OW5GO0BHpXl9onRddRBRal
eIXOtya57tSK7pHgwNMQyR2XCPlEegnwCXqKM9yFrq5jtABg662wqSe/jexHHLIe+CUh9Eo6oU4S
j4JlCRZszN5aE9fAHxNKko58cwbejxmRNuyYfgMH7Q8HEWTy2/F8pWiPUu+MCZkYmQt8Aev3uTUT
gqR8S80/DcUcg805SnDfepDLaIQfYwTLTisL1FOOpjJ0kLM2LO7zlURHPU0cjY83oV787kQqKY75
Dg849o7y8dl6HNGuqWYmhIEuhcJa+Dv8Tzf71yRUg+cBMMznnS6J4DCKNMQVf1FX/gVoee/En5Ix
132sf46TkQk6j8QSSxrD33l0L6rbj5HjUL3qh7slfYUur/zQtTzydxxt7aCMoS63sK4YfKHz8eV7
9N2wSjQTbQu1StMrLnuX0yFrMv1Y5tnRv0Iedli4TRs5KBd5YXXSYdDlHm3mts9hP/7y67KbKRSg
ydSjX2CaiocwLAf0TGxzjJ8xsZ33h+RIdu9rw+ynA78z4Vz03pP8brrUry1ku8KOQQ049DSgk6fY
WSy88r2G3r/8NZfEUJoSR5okfOGUP52ufajwPtr6ZUR+PLNQWaSYov7sqTnXD/N6RduKL0Wabi58
yfMe3MdJrL+HmwHcQzW1RRMr8Y5oaNFLvh7ifJaeynUsLWXllAsA/EI222d1leEfwPeiIEsrlSm5
B6C+woTDtg30SyqQLU6UgFTFEr0HvJ4DmGORPVNgNAw3km5g/kg0B7m1hGzf9xfb65Ie8twRK9ZJ
H/5JNVjZo4nxWcen5ALSz6WxHcobemDK4m5F3855krUjY+WtZ4u5kzMP4SE1+G3OXuxJf4AIcAb7
cqpo+IX0rt/NUZqfJgUnkCgqU7p7BaLgSUprisePOoUjGPmCSZeL+zZgsrJY60CsgZjy9MkXvsu1
TTYQ3locPiBZXgQw10jlPRtoha25r31OmTAya5lhihNCb30PpzZAgYGL21rvuax90rKAgsXp5oyb
Sv2sUha2Vqkh5TTB/9zjkpi1mHNjJcXwzK1o7Mei4I3zqfTE7lOzXxxE9ruSc0EoVv0U1azMi/EV
RThdwBS7U6l3t24Jxe75y6w4pR7rksS2i5CR9HnhFECY/8C6HpOINeyg/hnTgeVr2lJoX0/LOpp1
YbgCFNcrK6ms8U8uaNxdelfawWQZGAPHFamg2aaHI7RSeIkylYxHiPjd6At13diqJK5kEEKfYenP
cYjnEYk01IWS+mfNyrnYOBAnhv1GtJc2pM+er3RTQ6p0ZctFAJy0ZKrfc3VgpGHnXjm8JNgf1pHo
AY/CZI0Y7ukstOCiVfJCu3gwk82ln6raHwpJLiQ5/0MRu14+lEV/3wM5ysffbjaknBI/LgSpBT5Q
P2CJGhhsI0H/633zG2TbDSjw9P+Y+y+lsEfe3Wmby74pcYyIllt2KXwWvPdeRPQBhryOonobe6Lw
rUo9EI/3jCxRXTHri8mHeor3w+9URRWJ7ikGSLsHvhxJaU8EEjXisc8wuKe/lf6gmJBAe6V8Qdti
f0rXZli6QSyQbNgkgS1GmZt4JPQajo6AJk5mnoAJus5L/Kt6moG1n2XhvY6dYnsLIazYIblv0zLd
/VroGbP1JZlK/yuVslYWfAJpGByFvzrxJXyK0F7mUIGENshsGgiz8IYcYEl3/V6a3hN1mw7IlFEn
fjjHCy3iezGAj2AzPxmzOKgkyZAoJbf9BnF6GJGSMkF0SbFsuiwj2BAnRRMZ5riIcIwqb/LAUYan
hvHgOSD9zFQFzltcpKhQoXlmWpWbGVtLPQWCYapzz+vuiUNC9cG1CMOoRd0chG5iHhb2YRGQXutA
lsXVqhn+6JIKpbBSGSh6nMWkupqaDzcFBIrIyaRQK+E/HvKP9DO08QlHbMULVtdqmXRxcAWYGM3p
fYDmiZArEXnSDLdAeDkfGBX/LG3Y5nZXsS3mV8K4svQWff+hz92cV26GA5C6aazaqndTJ/2qY3+N
EHEikIltWd9UojHwtFWHBZWWefHhLwbj2RyWJn7AnoTlYFDSEgDKsDTm5YvdzCb1AipT4DKZhSfQ
uDm9CT0CEUfkZ+nZQ+QfbT2pT21CEvHCWJJiTUQh+bICjZpR0AssJpPkhpuGoNP4WR78fiY9csgc
/VvTXP9eUnkUVfMuOv3pb3x3Z+dpc0SEtXFrtEm+eJM6dI8V8JAnMBT+xCda/HUxqmICoJHCqDEe
yWBXH+NhL2dQ9wLnYGC8IXbAqJuzAth3a5DeeznvNrcYgBIowWYB8PtpWfhedcF4BOd/6gZRlzIr
WDFTCHfCekevNJZr7HoGGQT8yStC7NMMH/zcS86KfLTaiUvyJZbz77tls23tRf+RVGAXGlMFpPPb
vt1Uk1IMAPXuvP8xiGTIoWI3WkLZvxdQj5puI8hLtng2+E3ctyWf7oE2DBi015f7TVY/GovV3nlS
5CQUU2nSG2/RkOqHiuZd0IVp27mF00KxZVnnQ1juyGX+eqIh32g6Gf4iBShQL4rHUwPcT5QlbVCD
TAnOVg2X67jGOAs68kzq4l+o7xG9faGJkgQIEf94qtmvB3rmO35Sqi277u8JMg5ejI1LUBbgZanJ
lRTkkJTzQJHJnAfT41IPF48rP+/tpWGYP9gD3I93W+wAy5eZ1ndouiozAJdwvjcnmCE2sMcbTfPk
Gt4yZ7uIxhqn4VbPD6Xg8HMLO7ZosdGKAo4iO/9F5pR9ojkSlrDO3eLd2nvrsrWn9t+gRX9bLnnU
ivVNsN5OENwgRR71hPKeARadYPMWOcnnuK33d74JKv1nyNk5F0pfuIvXSOqnp1AUCVyLYOCF9xy9
uX12l58acisp+CAxWAf5G32kVdsftz2myMLPzD9+Lx4yXLQkcbp6zVwDGJdVjoTd5rHs9vtRa/KH
G5eyOaLMqLwCjByVPosoWI10gRQHUDNx1IKEaRQwkrHHK+W7oe9MBR442OXlDNuYtFMlMrJAabZz
EmLiEC1igT5nHl/nwP3WwU/Ax8uLTcUWcB8BpQkAwx/Qjn0N1ZthSwK//soOo8gRQljHT9MX/w7P
eATUAnaG5FmhKAHj85/QiGYgqU2S+bQJONWZAp/5T2tAlCZsgyqdYXTBeedOSG2iR8fpUZ8KIDLL
Dg/eytAoGCzbga/zMVtv89SeHI1G1VmEMAHNIzusNF1V2ZvjY6Q48IrbbF6G9yddbf9jeDTVpFVl
Gol0DpO27ggq++vtgfR6PCRJaQr+4TjtXpPvaMl8GICvMT1spC1iQkzQbm66c9ULilEKAvCRBLCy
kpTxz1K0z2Q6lApP5UiXE3tiUKJV+nS0JRFxwaeCFsJEtMCChwEOT828Y7/svO5Pt8qV+zVQuU9P
EhPRHGG11CLn+3r4eqrzA9gl+wdeZAh/6MvWDrBVI5cgLn0fQ01bsWQCSEAgQM79mRHF80caaKI8
yUYvnKisCWvAJr4lordr3SlWRr5xr79fdGZhZkDkr0OyiZ/E2aZbERXWbdnC4ci5G2a9f97x7Mav
9QP9al1sLSU4IqKEBGeLCRftBRR2XTB3K0/g++nO520tTYm+VGeWQ+a0vRKoWbPTXxtHkhXvAF6J
iTfbqUefInf6GrQs1sfNd3mU/jGI8G+gzjZRjz4b7d0MRM42BP19IfQi1ceOWXMJti1yhfxPIf/P
6ulaEM+FfbLO05doXCjLnAho8G3A/ZxCRxuvrHdsoMQHlxCXFogLe9qNP3LD2ODuAqWGO2gJf0iT
eP9HQAqcA0B80f7TWR9YE4K6WJWf4M6nwJZuYvmD/HCG7FMqdOh8PYXpfUCm3ONwvkFwqOVSFIv0
INyGMUlf9YYBLZufZ+xDFdEJeg66ObwadijpU0aTCZmMdpq+AQz2Zr+tvLNgNcffvXYR5HvaWKwW
DWjZew9GE/fJSbvSM+CH7wCC7sECcOSQlOh5OlKUBOUrbOfP/A+fMcSc8iDxMVLaE+MuYApOq5RZ
EI319ACWkWCUzBMXWugDe69LJPxVIjMelHVykFFth/4IxDLzHlN1mvncbpxUUa2NMEnU1T7RSE/y
lytn+Zm5QbpT7lJ2fzJGAOGlWyAehEfBJBO+Cv6HbYR5be56fgDRcBI1d6aEDDcNOJvwwk842mJe
oAnSuIJTgPaXQGhtWywXlbejzphtjTZHo2KaQfBiyGMSZQVXe4gFIGIptniFxEkCywJFpeHSycvj
RDv5HZKgA0Yr66g0w0Y+D5akA8cEDosZsaJMFaMhTnGwcefab1YugiQU5BLDehyptGt+U1Vlrntr
uF2WNMwd9MJLRucbvNPEyjeMuCXkG/dzxDsP7JRYnbgd2XG745T3pnuh4IRp/9ceFUT3OpF7QD0s
i1mK25bNPwbXTYzNCzk/+ckvjimfhSWoDf/TxzsUii/3hs+pvE8zJ0mhvVESdgv2ERKpPqFPzftV
XuYWEiyrgMcpbInPg0jD0GMLXPM9QRQPgTsQgc9yE9hA7ugI9HNeFApcN825U7LhU5XBUasJr+1V
dzn/Nh4NmbpgVF6YghbcGT924rm37FDeuNiPvaGnhX/a2AYJ5h8C4A7EQ5wOWPh5RO2dAL7d8t1i
Qi1Rb3BdtJ50HGA3eAmDhcxETkKQdGW+9b15mYMqhaAeaA69B6qMrLh3xb8CazvntS43Pejo8nd4
mEd4wxX8Pud7/JeNCPvfyNdG6GbMRNRumv2hGE3MUk9mqljXWK8iE6nuORL+qEZUuU0Z8cIIN9yK
9xSj5NNQMZ9QK6XmOgi4gYNbjG8HRw9ajt8nId4E2Rhum+tt9O/UbtIhXGEggRwm6MoelrFkPbdy
r9/38lAXSkX3I8NVswKqCfjy4cokfzl6Wy+tU1wojFZ9qVON8kcxrNd/4oin099E3Lz2Kc5IychS
Y9hB5KdAS8N0IefSOjPVL/iXSckwvoOMZm3kSd+sCBFAenZsbOw9d81xxzbkDN6E1EBsMMaGEGR/
bpEU7/IIRqPPWZSIozsVHI7f1aJHeAdvufwayhxKK+3kE952FO8Cu30+u5NdpoyIFs7mvU9xbBJU
Tv8Eco5RwaubCMqC+32mM0zhcbAq3mI7I7FkfmyWbW2l4PCvRAI3BEKotOP1iuxHOVOfhU/7vzZa
FbjCXITZtUnkRzyk2YUFkrGxeymVxE8CaYPQPvdECz74gi7XVr/a/R9Q2TPz2B+N0WQ6sq4W0BNW
TsTijS0q/VblrVsLvYReKKsp6Iyf6CBeh02WcTWlXEMN56+o+vMcUAo798gQLIPv/NWtjOJLldiy
rpgR76yYDLIV0wXTXrcqQT337PaABX4K/2ARoTCOqg9ZRtmpz3snXUqTPf5mXEfBcuDG02Bc09Fx
glDflv7AXuv4Y8/fQwWiup84PMtU7/+S0Z2Argrrujw6qLgv0Muw8gXUlezN4JUCy1O/LknKnHzP
5lcAizW0gVyx05UfYcA/TOgXrLEFyg/KzOvCqg7wTL/s2lcC/CWxpJzRY0TVIEf1bbbiU3RvvP6r
i06dYthVVyeyFL3uoKFeA7b7za91QwHQ9waF8pTK9PfprEhbZ0k51Rs+27hpmATtznZTuDGo7MjP
nOO5UlMLUqxzkj1rovmxUXOcud/lTIrnnxCQD1Vl8plDMZrBTBmAgdaWYoAXkEgZG64rqRlEXirC
LRbZ4fXqyIjbFKyDiugDzSnurv01KqMBH3WAJ311s2XTGbrDYO5uP+b/r5O+IQFNS5y4+Y047cjr
4ELJlHYyd3MsWKzATS9nrCOwWLYyyz5PNfPQoJDfA4eGTEwQG7d+9nVuOtrc6sebEtmam0SaVvxr
kvrNC2HUdBmOqnoc0QXCvXRUb5sxL5EOtOVhYv9uUCdrGIW8V4pdAHzhaYgm5XZFFfBX7fZsXUGy
bHct+XCAgCSb+NJIK2Lv5HujKrBg6FZC0t89AchFjM2F/vdJGCh2Il0yZx545s8UMQq76NdDyTx7
e1jeyoKHQ3rg7nmy9kDs0tIv0bnXuitfhvwJYe8wTKGWbpp3CfWireYAUMpwsqiuhbuCJbeTtSXD
avGiU39TfRt4hb70AzINnRrbD0q1WH0gZV38DwikM4Vq0upasMSZzhrcF7TdOZDOx5yn0wSEc9P0
rnp/FOat4UrGQPDgdPDl09yf9yvY1PQp+JjxRoyoCqum1mjTT6iFGpgfU5xtvm0zCPZBS18QuITW
scUMsk5PxcHtFx+6CZ1CkSsH66QF69mB1BUCDMFJFgYh9CLd/gDPXAJsfWfgcvgujkKxuxbBlvsM
cXzUtDp9f/mJwa2tB9QoeI5JAzueZcKT+kJ5rD+GWrIEOI+ovGCz/bje4OW9QgWKzTye71fMopYi
FNHuw4/RozMyUFzqrBqKNSAIeqLK92c44XTARKb3TVxF9i77/9DrvA65+3m5dVPnV7wJ+A0qYiMg
vCiSBj3qbwf2/SnOajeoBKcAm/ElCjKZn8uIYBrpW67ts006HTUcQLkPJiKMFgXB6mVWGYRWRWMV
gi4V56Rj6fm4/LCzOvaKXuHFgFBtShcmdjFwyBbqw37gz4Wm8SibeLh+gNKKn3ou3aIammzRbDPY
7+uTNH8CmiPC4fCLDo0r+O9HjnC0hooJrBJt5eb8s9BkoazYeGhLfS5NT9IX1yT5l5G2RlyUtsfG
4E9odhm+ojoiw5GkU+xEfKtex/QL1OTIhP7mJd9hySdRPLHpgAC6ynRUjYzlhP85d2MH+29zkAeB
iEqatxofBBzvzf3Uq8XGlW7yj8WmaXCz5Q5Tn+EA7uRMqJ35ZzdnoG4Hzd8eOTdST30wBkfQaFPc
9l2ifQuda6hKyzV8jpEMO3z+pja/Z0lsvylXe4HAWkSA9E5oip/VY/erba538rPYcIv5EhYhd22b
5PXsbSBKpTyKtXWBoZChsrrZQZiMEpuT+B/qfbK93GWWX3XG0f/pCVc9HvgkvFInHkGiZk+OxBPD
cnkPnHnHf7tb7gfz5I66pCmV3jRoin5VomgfpF/MGzUx3dfOszRtuyqIXpOHeJHopLfYCtnhUNeT
5FO1HWhNAfga8yTxFve16pO1QE60zWBO0o3XN9Uk8zF6qkFl3AgPaK1bG24+L46s1i5sDx7L0WIG
Pfks5/NTQj1LzdymQWrdDRln6fcunBfO4RVJKWWHO72xPKqzZkp3riw1toSjnQ1MaxAmag6guDr3
VcvZo7bGF7LB7jVnW8LO2F8MrzlsUGaOTIrZGSmpPcjYxLgclg5JfmIEZME0nPf4nev6vJcaS3Si
sVji0/Ox897BgC4wTYfdAz+tDbNk+PT5W3qA1JXRyWPUUWZRkYKxLW3L6hsLXQ0ZZZCNL8rzKtQ8
vBXARuMEWlF6re7Z/IBH4Er8sHrGsLr7ZW4Iv9KWo6jE/qUST/l/zQKaPwGo7gOqHfz0/MrDfZQC
kDf0eb4ePtOpOZ15SK496mUN/nHD1C4pKjLntSapXbw/9L+SkAhCtOK2T+o2G8nBs0X2X+tgymPz
oPs7b5yXihS47eFKYL4u4hOegB+a2pc1c9nrDwr6vTNW8+/DB2P6cGT53B8EDfQbcHIWEpGpXn9T
aaH3N4UtM01pEeupLXqUcAImnmuv5neAWO85tNLl/YGQCuCq9CYUO+/s1t96HYkwECOA9hnFdaxz
MYkbiKkil/Z7u3KQq1b6oYY5htUHJ28XiHbyGvFpQfdqwL8TfM35ZTsyDnMHbEt9husQqY09+ZDB
SZUjudgb1pl90eOM1ZkKiJCrwrEMKEpfjMGpRnqdgZvenAAhhHw2HGR0Nzaoekdo+cU9VG9gbIml
3+d3kxudjZVcH64wT+eVhbj3qTEqiP0XM/J6iw03+s7u7R9+T5hJeURa1ZXl1SQs1v9ATv78879N
y0PAHukXkt8d5R88/GNPO/JYeEtkb5bwXvv//+6r6dr1MWu/fJVHIqxeMfIQprvzmb2/iHBdPXAd
K5O2srsWy50SV+Ka//SB+JQadXt6+/KjeDO/X/R0ptpfueu7DyIjdXM6cQ7S0ZYEOjbPeygx6xrO
QH+rwFgSPDoMtFFVyjAb3jLOJPqKlmMXj2lhFXrf/9e3f5UX9wEFh0jnZCRzzVz5Cx725LAV12Wc
iKh4IKxa+WbPZjOGA4LoSe6tXhyZssKNwkX4CeZzJPwRGuMlimAD9ggXfCKL7I1cUJEUYmb8IY5x
IDU2aUkYVXv5cCBEh1e0TEO1/4mfRLG7ZG1khyEWOmUZwSldq7rmguk1hE46tgVd00d2aO72kFgi
DVGYJ6G2ugu8X7X7BbIIZjJRqbNgha8bRRgClYSwVIfuLePeKG5xn9QczqsOr78GxZv0fVkw6mbR
RhCogdvTlnkPhzCbL4iNChelBwn8ZTHnOGdA8EUwwy4FhVvoJdWxw+er4kd1F2eAlg2GI4gnqpWm
csUonxjTZtOOAGoOXiEKpX+pFh+a8GI2GvmG7JshHLVNYenfF1kY36f0Rs+wYq4TG2N43w7Sq0B5
Rr+MLwotaUfdKDnhX11RGgl8Nvzxgj4rhdAj8LD3VwrgmRz+iNQiuGXcJJjPZottd5v1Gs+AVYkk
TpyX6DAPOry6Ozs557YCI266ZGNmScowNnDR8i1kxbDG8h9YY2j2n69FaEGwbqWbi03cgELALS7B
/L1d/Bk9O3lQ32Qp84aLs8/mdPZKHSOZa27UMPghGoI0XJe6noDZakvGN8yJIZ/e1LuYlUkB/1kI
olcmLTa9Yu1iWiI8vl2co+B/eHo5/6+lbqmSwm3EZ762vrCtTC0YxJwPFbGMaAxVQIIIwYNyuJnu
udbNvfzenAN1Z+n8jCo9CS9g9ORmkpHZKfCg1dux1oIzdzyxiQ8SMqWuJMI+kZJA40rErz0d1oYy
lu/2J9VdbtqtZt410Aq1Tj5rTyWj2++gSjKd/CS9LgTcxT2ApB06iDsNNCePR+n8BNsN1nOzB/jQ
pJO0DIAhRAGcIhIgKlYcCUVER9Qunstm+KqW2VXuyMWumc1wkXpbxkLEEwMO4vmHr4OeryQyPMSL
Pz+60WBZyyxBnVo2M93cenDHgwUosMktscgqrCTPerML2Wmaq+67STQKOZyB9cVkWD9g0jf+hJBc
Z9zz/QK1355vSv4J5hb+1t8YMWHoD8yaDiVQaKHp1H3yAH+HemBPxP5OXt2e/YSaHSl1rZ4kXUMi
zhylF8OfvT3RlXmVH7HvJ6QaX2SjoBuzcz9r2JEQNzMTF4dDnnXmQCCxus+gdDxVfpCC4CYmm+wN
qcstFNx9Ta0MWIAETIK6SEcPG9pCd94EtWxor2PWvC2QyPdj1wXLDLMMA344bxWtWzZbavdYXsB1
2KrOJTkM+cbspVi/TqC/TfpaBd1wRxplEhv/l6WCWgjYClc2+8ajgjWsKrPROssGJwrSGoFKLqGe
KBhnRattBGZEaFUhJhFYVbz71zDXkqJZsLPl3pW6cAs7GBlbE9jL8zbTiUWNsQU9hhP8cXN0lIEu
+2fNo3FxBtFZo4mFxUPyEgwZnDRtOXF0VB+MGPgTTAkEPzX1+m5pCiMrxlwonOrsf35RYIod3ud/
GdE/DjFFPsTwgTEZJmVZ7uEgJFxOPTyjL/9Tfo4HkE550FXWYwnYSFaMUNHoPxIR923tax6uOG5f
pd2TGh43ZofbVxNouDIDFVbpTVoH6D2fx+HKmJAlf4UbCL6ps5Ue9KG2DYl8RjdqJV8u+vArSDX5
pE6hcFfWpKuapOubaMT5ISyprWgLrOG8EI5iUVshQrK4H4asOQ+a6vd3Ctzjrqxrz2Fm1R0GIdKv
ZOJJ/vsniYSjyrjthGpju17JIdRwYZPujJJElgXSUnPHj4OfLxpsHjW1anc8wnH3pIqmafhgM4gA
L36bQ2ZedfcikRdh7Pqb1+2EA1wa0xMdKsD69W4NxSTTek1SJQHYdi65PVc0wh05UP5rge0m6lha
R6rJjbBNSe/zMXpAKJM6a9hWtSVEPof5CQ3BQEYdhcLwrvfilr06ez82EFT8zdUlA1beuFPK2pcq
uWBialfTqSKd7+qOMlqOK2L2FlX+cW5Zrffn8CHq/QRjvScO2TNG5YW6W1Ud/lNdoH7/retRZBYv
zo6baFmtB+rHyVjQIsy/baYhD8CkuwsQjx6WSNu3UB7nlLRu4+U9f5xKtmp4BcL7gEscPw9FcmEw
ANxA5Aod1aeNfYqCqQjeoW7v6k6UsI1EVK4+SR/5QF5W/nGwtDXk2Obixb5Hh15Xv2RPYxT2V2Dw
sbv33THxI3oLE9kmPE0TzVPgXZtoycayoFNAkxBgN+sP1e9qC0X/TAnNxxHnpselovWRLpHT8qEz
Gni01zS0b472PpMnkM6CoyzmFR/eQoBmPiUVA88k3U2Z2A2OZMm5CxxVc4/qX/DN1PA5QkC0BvwG
OKcZwMDZAqHNWBRrTQiykB0SXwCatYAzdrNWpw0KzKVCRe6yy0qFzA4k0+WK3Dv0UqJ3YBJM53XR
1MlTr/V0OukpnHUPKIC8ae7+MXTIyVJrRkEubmidESKhlhuDXDCiwpo+uGK3/k5rlszl+KUu8iQJ
Gtqj752o+48aR5aa9Vi4DpEjFtIptYZLW+xkxGX2rwNgU9Pxu/rY92Xtx4dnVrmnoOBx2/SSj+xB
9QNcN9E9X1c4YIzmqPS1Ky4v3Mqj19iHN0W5DytitMrBikQgrME3RLRYZuMLiP5Xcffkl2YSGh5D
ra62g2K+A+kHzwhNgMpTOYoGltR/hA99zEc4LX4NormebDRjjx33eDvOgOACXizuTHB6+3zeY+4O
9dppXutc35LYnlHLlYCvpJqnAOIwhTbkp858VUBC+FjaWayKpsP6qkOx/3gvckj6sZ0biB8zvd8A
Am+FGENEILFZPCqHQ7fFxQZld7uKWJMUWaDHRBhI1+SH5pRAEMc3PJZ1eHVqOIpjWvb1Fuk/ITIg
o1C/0X1BqX56dtep9rZ8RBmWxWduXxsAtjyMdEKCSGag3XJfr55WO+zIh7GI22f4UN8+Uf1TCpH+
khzL/Fc5u1MKISinAhEJ/A+g9WB6j/qw2WtSVQXziY+dNeSB1G2mAuRHv3dHWV5NEwNJvo0gTubs
bWJlfv0PenJ82WAnMNkSkaFi0kmGKTeGIOxKb7fUMiDreIa7dy1Na5VgdfvJtjKcDrnZJ+OPBXsH
6UI/WvIl9CYpGpnMTrOhpcleDB4f9lRSvvaGwiYqZTsrwxiWDk88KAn0T2LXnADMU7q69Y+oRcdV
vIavBJMi5UXsacjT28iuDaM5CiR76Tb4ESGEJNpaZnMtOsmdZK0dcCpfLYcHWhXxJPvcShcq8pjR
nHgaC79TRHIIdWnEY3e8Zxh3BGoXYax7oYKIZaUa8Ovh2RvG9kU9oboN3JolLAOs8jUZIk4diG+J
zYjQ2p3FOdK7X/KGolAZ2WPb7yqaUX7BJmW+v6+ErDUVghkJO4QhX/oe+CrnhqsrQNODdIEOjpVk
49rHCAgSkZ97H6utWxrHiT8FYm5A+gTZTbJ4NtkJj05CkGOz7ytXHAWTwu0dKf8gGYU4XVVzkG87
zeAdWX4WVy26FDWON2/Wb9BxBt2cla2pWClEHkF9OWL8oOSMtguT/Cw3+n+OEnQK6qSXGRG+LvsE
m0eY4arV3j/0fAO1QhrByAaB2MYkj9JSzP89AogwDPoeNeP6iLzG94IBU6qTpmA5xWduSLUQir+/
LTDkwd5vhEK1cFYd/AgfT8V06ICJOsKzIXYA33uHjFkZlMFO60npVEyOgeMTHHEaXTJKtkl+eTvp
VJU0f6mcZp5R4rCNv8yUCbjKza83HwpaEQFY1ouRffEyeIbxWoGyGegU1esmNpUbqYXTlMPIqZkf
pwgWsUq4o4UeFJ8ykTXGVCcCr6rFHgHr03FbHRoUrx8cNWPd7+KdWcSpfc92evZGOHZxj2TGKXj/
PTEjaWspXlzjqL+VX3UbShmb0GyalOXt2cTFMolnpU8i6f+3kO8QhVLT8vJB9569tyJROkPJdqGI
Rmia8nepgVqM5wQYDl2C2T6KSCe1TAJbunSLnFOyjLRijjL8+w25XaS1XiRRb5byorwNjRbfa274
xRK0L2DFxG2uIDcQsHchviQyRqd2MLoNIyVr4x2riOYX+bzVFORK9AhAMYqi5l0dsBzygJXi1VfF
JtxHq5xerv5bBwKglPaQX7zh4QVs8FNs6jSHwOgILKdX+ZBh1Gd7dQ/RLT+Dv8FYRgRewuiqOurL
xzem+lRcLGUO4wK4RRHo4eZOCcPhoHdHHgTHhy5Rfsyuy6E1DvJ2eLxUh1xDSrdxFPumvZgKeA1G
sn5pIKL+xv+7fejXj4ga3BGeEK9YsQ0OoYF38EbWhi0HXf77PDVB0VQY++jYW/gNc8qmX627EDii
k6nU8z35oStV4wVFL0O/SugntdHRlClEiv95drRTmc4lNBdVtbticwdYPOeylT1qS/heX8yItQrK
R2QrR/KQNWxtBcBYDPOaWU7qG88Im/KkiOjNi8Rqh9lGAGwYS6hdFILULjZBnytPIjxDfOGarawf
n42HBYvoNA6p95nOo/S8ihYGXC79aca7mYdbbangkbHuj8vOkSl9mEI8Ahm3c2eZUeQDR0WXaB/8
xBGbM7bBFBb01gtd1lfdv2TRELx+0u7/+o1NBns8M+zvX4rKQ83ENEWKb+WvHzQNTWNYY/iW7ozF
CcDUMqQakJ58lPjceM2z4vX3Ln6gE+9PQS1MKVEmbvXjoZCnVjMM57vkki+Qfv+dsfmpTJVq4qij
0JV25r00P+dFAGz64PU1uVquqN5ABEU7B5S6VuU+dOqy1pWASd674/pWC2g5slZURpp0irgF0zOa
TP1KUkugdqgjElLQYSAD87icE0Xhyc8KcYGoOqaU2XlgIL4JhhQJc1hYTu8dabls6UUGl6syxoff
Fy2XxqxV/nFkfZtzwoIuBDXvFXoTn5eBKvfsx57TEgWZfmGhKuIZAFg/dYQhAKc3yeKoMgR3/wpQ
bxnfYIMTSupqxxa1TpkFIq0NxCCw6afotvnmMPQNTTq2PTRPaMgPL3lHXHuSRQfwQxQ5TaXclPS+
fV7KI64Tk9RDd1ofK0uxo9HwIW9ED5z/C5fMPXAyKq5oeNbynuo6EukEJ0Zjlb7z0Hp+PFurFz6h
4FFF0SZt4gH593XN0m7ULheXmH1tiA9fYzwvcuPrTxESBP44Q4CuVMcZc3dglGQZ10C4OficBJ0X
QzcScKkKl3+uwsvV1JmrrmOklYONSgQQlo3PmUWj/Iqi61UOGs3XSDyvJHZM8/KLHkLG7ityfEQC
m0VY/nbmc3PP3m2wtOKPkY1XMNuQsVp80DBktRsvYpFT5e0AFFe4i/3Jage1FwshLFlznrEVfFrJ
y7BRJUbN5Zyx0a4HUAoWK5hTpTWoHELEsO6oOBuMDQYIfDozt6Te7N1Lab4SG50k202Rg//0P9tq
JqFJvojjSiuXkRXu3dfKugbMuBF53NN2dDfHbJvxRI5vYr1NGmqI3hhEtaBSRqThDkgAX7x8ZHpe
cfzU98ZohbV1/K/AzpxFLI1Z7IzSyD8oW8NL8Z5ZBVjQeBb6VtB01m0r6l9JLGBaF73wF2KYbGIU
3iLC1D7fwuPtyDnlnQ3fWd9o9dRATO20G8OX3oJcQeY9HZRCgd23opgy8991MQAgKOIfCC/hKFxc
dZRhtctvEyhkAGePgGJ7qHqAkSANQQZ8QNWDv3eKnl1fZMhqSYBpHFUY6O83NTf4wIAKltqxCQJ3
Xev4I3XM5G5M94Tb27B1tVT5ZfYqbPkkiIhFQFJ2QUGAew/w1S1YIbUJphzbJK3a03tz276oDAdL
FBwv7fJD1S5cL+qFrRF86KP7syyjUtfMsCx1K5gVQz1jp5kAF9hJcn0IbDX3JfxHaIPnCKpBhgID
FcfEAeELU5BXEO2xZR6+rC8my3SMu8RXPwefpfM/7PLA6MIMQk70p5o/M29SL2Z2clp7CXGSRbKb
g3blpfg3vE8gaoVnrLzkZwqXlu606dT+/ahG6wNQoc8NuMJ5wN/fz+k5uNdlVx8BOTkNUo7O24D1
g2MvqFwj1w1kBgjOx7wXPLzHt4Pr2EAw9pEtle0l2TGX1JMOu21C9ldnk1MyKjA9rHKiVpXXQ4MN
OIfuLQxdSXkhSfLvKmMBynQ1xS88tqsdj8nBn065bndrgYMgSY/yLdlthnpgQEFJU8QoIfM1ggBY
LLXDeuPAeONkxGScIp6y1EymUrwg/nx9cdrcLv5WPocUT8G7XNdvR7toVX0A0J9cCwTo5iW9AM3J
Bg0V9NgzwJYaBqF/x0nGCBrwPQIPEe5rIc4Fo49joC/3ys5toDiw/YM/FnmVNKhs4RKLhwktEVgr
DVX3jr6gqrbm+NrUjcyw8UQIFs2Ep2jjxvOqYuZ+i0S6ZjxQbsqHaxUe3wI2tMhPhOQ+mCAER98r
oYLG3sGcp7LBqLdgR/VR202UztCd/4KGgRY+zcJgwDaEyi+bLlXf8ggW/MKU2j2Tq1FoU+M5AzT1
rGDI/TGbvzUX7BsdX2sgt4gvDIjuL0BIsvwDD3HupqLbF5jSopoV4EWSmse5cBtRvcmTkd3jtBq9
wRh97aswKMNEFuB7YDtkKNo5K50iBzaPCIPsJtAGV7ZhV9viEMEn4Mh141m4atsP1JknedL5uekB
gbxstN2cwM0ybA+fv56G37ADbBonquYKRHOrk8UQ1euxfCdh5r44qnqxd45fXxZm67ykFn/SIsBI
4tEw5LO265Jx8q5gWD9FoA4mS2wA5kvB2E/nDXQ8GtVw9jOQBqoMUSnA2vxKENASFxOufL6XdXX1
+qiuxA7zbqHKWvBnzhL2RVM5b+4otyKHeR92dU24fj7Cr5I9T7yB3PJ1Os8B9rNDKbA0GH1gSHRD
gCQcGd3q0DkTMizo8O70KmCGloodykKlR3AUkrMBSrn2tKnYrtuThT1uV32LJuiKC5QCwcUAqpcJ
uBu3CGEJHtTpLwAOdmGc4AapstG6Vs0Mfd3AU/QOHgtqni/dCkjVIDK4qwtHMTmXqj98F+P3ghtU
tPY9IhkG0jYcXAVp+ZGrQwIpMrbnylXsqzJUMsDkDRiO2SDX0m2ZAVdQNbdz6M3Ej/n+zjM6O/cJ
cZMwD2X+O6g4Y+ChH6ONFC+uEzFELzY9KGytbgJUAkyJHhMoBPVZsbUkInbxyPNrbOFp2uF9W5Ri
46tMfYF3IbUf1vbtNvgyH57s2ilt4H+AZGllkQ2dJ1aFy159idyPt7XOZaI5iXwZ5CLXVHbwzTks
sQ1JGdK//Ip3syqcbRjihEe6XXoSNTRHH1VJHWTiprBsAd/07/IpW+HRzbuEvIC0dAMl/sb9mrgf
0YMk1uGKpdO4rtVhpETVZk9TJxgeqxUbxLNpr+DGVO3WrKWxTaJ3NUCJZVLAIfM8c1IwpxAY4iZQ
sHZ0BMkl4CA6vElCGp9SQoRdc7qCmeN76AHch3+i3UtWiyhIbmUAfwWwE0zpPi9n9pVZ3XvYMWxx
av5BOOoRLSiseGKZBKiuH6ab7YDfZLIadP+u78nFhR+ZFnlH0XpLOSzw9dMGcDvrhSFavm5L9ItV
yige0rW2Pkyk+n/ZXA2KdXg9Dszyhh+CMPe7MrC22MFe9LtmYPHSIoQfBOfgrURg9+26AsBxpjkj
J4lxcHt8cA92ceIN/OWqOCEIGquCMAeqJ9HaHurlNhFfJ9gDGWcS6MsvX+zsWQ2h2xJMnFHkp8Xg
7DajQCaWGBB1W0zZsY/wm6HpriTuG0j/KwPbUBJsl8SJlbplfh6cGPFGssPulwS9KE70YdUncUaC
TgwJolz0YwmSXUPyERCjnfyjSMmj7d3RSh3NsrUKlZamQ5v1Z+AFXzkLLloAjulN2xE/+heGpXaK
LEviqftWqePPajl/YhgVslS5nyFWVLNgtt7MuxFdIjdozPWzjbHVxJ2DMB1xstca685xgAyWAQBZ
3NFRZnX6ekcf7RqG8yz67XIeZI347PFH+mm0r859e0fUrK5+zrUF9HqGP3Ip6QiG9ymUeZz/45mR
By/FvpTkrcqrQrOm4wQVQXCJMpgzawFA/1RQDSJIOi0EuGpkqIjzo5Rus1C5R2mWg3JvU5lH8rab
OLDOFs/aNRNx3zq1JjWo5leSrlDFYivfYG919GOJ+HsLvceMfe+syuxmt829OwfujOO50nvaFF5e
dc7K+0yYwfpnexPOni3s+nORH6DYY9WnJkby+dy4ZmHWeipEtfjVVMr16p8iRJSzUpDPVa6n7VhV
7mG9T7hNNK27IfXFGye2Y+iXVizMK4T0IlNu1Cf83wZq2X3LjxJJIz5qjDFN1RoYZy6YVtmG97vb
lO9Zu0lW6Jpnum391Ixxx+Sh9uh3uaBF+AGDwIlpWn1BG6j0kZobMEoETf+3JBW/J1fgYRkCmzkM
BVUoiYklJNaVQByCXN6GOeYRUkBd518Q8P0XblhcBzz5lvLRfp15O17A1us+GlgQP+o2htG1y+oP
sffkky0evpszgNDoRvWT2pcxDAFQX5gVAb+h82pfEOSNCeO0lphxJGL5MNnlK90A5preFtW2Ul+V
od8sP7XGX2TgN7blSXDfEp2ev4PM7NtWw2uTqg51XaLUAPwQM2Kp0jqcQjxzM9KhdnfGsexNwjk0
i4lH7+yw/tCRwozgxAWqzj14/PAAbVbgrCtBAMyfW/IJ5PGfldVguqkdMFfnPw3FNq3kaa/fmGwL
QqXglLvK9hvtt1++np9MWMrjZW4db7If3N5jlyPlKcoVCBjjQ8Tm6ssdKrk+Osx/t8nRu+om/5Ya
LiRgZzfDQBHuy/6i08P6ApTOCtjfJTcbJXB5gYVcu1Ll/EOFGjonPqD4iB5wcPTcPSXbCDJQYw/9
kBkkSR/MIpo83XOTTzE53fvYuuX+zAYsDsiYmZLGIpERtLG+sSNbxbZF7bkG22oe8oxRVk6Sbmux
euic6jpy3bZCcewA18jq8uhO9V+sgxdqiOm3v4ecB9hvxz/Ws/p0MvWesu7ARKjRMcSD9Q4TCErX
7njK+D/CeVwONbDxQWV6bgquY9OVo/J+1/3aWgE419nVBoy6ZhhSa1lIvv9fY6e3JA7xODg0br2d
4Qjcwmt+1UW/7AcqkdLaJcfn0MSJf6hKtADEpvs9xp43xiHTZQsx2pTeT9IKNayDrlzQdqWALq6+
dMIXQ6z3Y9SXp4ecEpEB5KdGcPOF6uyQqxvgO5asVE2qbfEoGclElU4w6JgQM00K7tf33Hwm5aQ6
JFXbnOtY4wIriZ9+XJsZMKc+C6SJrCBVd+kq+n2ZqwVXr5HTUrjb4VKu6PovefpMdsL48P13lyhP
ZNRxvq03rxj+epz7GNvZaPLUn6Lf6n+P1Czdn392l53VH7tHgosKEC0WLGe9LEbHLFH7wtVpdd0p
rn7DD4VMyAjg/jrcGnSlLuJeL9DV32SMW5j0QaGVOHYRpEsNPSeIgLlxC9O8U0Wt/Es5ctK10qQH
T6nMnRLwmZFJcK3mpgYGrsJ6qgy1tZJEgjnp59nLeYYG3VDasqfDbtrvladSIA7GgSb6N1Z67F0x
cmFUrmh9iC9tivN5aiWA/pRJ7O/npxrcDZkE5+s5OEc/nczNEeUEI7SDNkVQOZTs5WlLIwgBqHFt
RJliOcb7Dzsi/k+P9v08h6G7juRAF6CXRZhOv2s5D22lip9jIlPXSYZ/OUfGwTUvnT4sIrYKK9Zd
9e2SbhmIXZOdsau7JYJt5eTrM8OkqQxB178hrCXiiiync0iRzG/T/BoYjPvdNDmgTVXbuB02RUs/
ykjPA1LQI8w32uKF13VlCPPufwUQGzFZ20M7bcBNEy5DuAlGGR0JKI2ELbkFYBysodZqvyrdVIdK
A5KtMNkuzUGLztlVwXNLvkDjcj3iX7+iZLu7TmKBLmKWpVj6QPiF0+qx6bH3rfRQsajJAfHduE9N
JdyVObr0wDxZVfoYf4+T32Hb7ZHs/PCRnA7w73Qgll42YRRx71fqvEAmFVFd0n1OwOunFKWwv1ZL
lgU/jy/I+0EFbtwAtr/8DUJENnqYnXdu8puzhDX1CUBqTletMdOlxZflbOIh4Lmt9fWmbIluLYFB
K+F7tlt7T0+//MkcuD6QEONB5MsS/+hDiBGW0AQVVgc/ABOlJwNVNcGNFTJ3i8mPdAjr5M/eGK/b
IpGy3jKZV3tXlgxv5Br4XWhy4jo/khbavhrjnRquXrVf6sjWRE7VlhsrMJ1EGgPlkm6JJvSOZCeK
JkEQTCuW+E/vaHU4MKA/2iUoyQoKnr2MDpp92LUeqPw1AutA38nMUBT3lrdZcj6qWMBsDcHE6s4Y
EeVYLyS9WEzJNLMheRR2ErCnTiIUFgJcvWdPAS0bGX9ixFSlwlcmRcsvTiKiI2nwa508Cj2RhtK9
DEZBfSNXFhcnWZhgArhElTxcGzbbWspb/mRjPo6HetC65dkuLlDjFdFkc63bdBQXGi9qoZmsAXQl
Nc3I5mnUs2Aq764xCZDWisCtkVb0illELLaOB91u+ZdVQg3AvWkbMNayZIbJ5lsIsrOwcO2dti63
wIiQkfI2OpztE/HqDUpd5fepVsQUqlW10sAHin0Jm7H3tYyw3jNKZvlzXpZcJyQ0gmhSU1YaHMTJ
MX2mDNIq8gGbpueJ2UU1HuZlFd5orzeGxyTFDAeWCfXpL+Loo1n5csxlO2nK5oDTTMJEooIjedJn
ITtfTO3mxBpFzCxQVGob0ls5pm776Q+fAlehN7xpFgJz9ApIGvdR4j5DOVaEUkF/Hijak/SARP19
90Kjh4B7RHhV3FNQ++QJTnvfasSS2CqCGENVVE4+byN/wxRdLQBBVPhiWba6ZxBX1EqXCnEZnASD
uIi+ZbasfTjv/kGJL+Z+sewMGjCAkGNcNCg+r7bjAJb5vUozBHH6+unjV4zYTlzzHnXmAWCayl66
YPg68uQ45ufAm3pw2UFCun8bLy4jFgMwjuciT5om6qv4WjhFgmRI4JIvlLDzD7tZGzuf26+xqPbM
ydGoqRiOC2+9xhWzFf+701shwM+WOXSnDSnSLwhx6/g1pIUtb7NGDGxUNjJFI9FEm+DthtX0mTCO
ij7Sv7FWA64lrwul4j8MYXtLA9qLABRpDPMk8jSRIfeHfaERp2bmhnlLy/h5w3LV444/1//iwveR
UQlUUvdEAiQquwiMq8IyuBy37ukkGRR8mSLQbirwIDn10l17kUwKOtg76bubjYtULAaZAepCNWW5
wS937dwKEy+DpKbK+sm8pDRxWSdO+ixzCsc/Mc95ou+lAVS4u2gQ2K0UZM23/Lr8zd4B+9zY2ZIr
QoUn8l4cDpGdFaZ0XQvRwBj2bkQTXcFP7gwCAz8EKAt6YSb1RrVgk5CqzO7HU/AP8J0Fpf+hPoiy
1ZnZzXcJTc99HX/3/yxAyWYJRh32wkt4TfWcXPAjRu5sovQCALLRfbfKSSWSaqF48V0j+V5K4B/R
A22ESBNZuK2+p5ym5ZmGRYlqXxssksKlDEsrLDouyTZb4/hoWzy22N1KFjoGo7aPunMbjgcm0tTN
R9qR4ArlubH17s7gvxG+l2WJF/L4lYNSNQGeOA6c6sLRNsqB9VS6HaGe8GNhcMPzQpNV7nIdlgIL
j/ZbHT+Tbq5bcTnQuRTybTwIm7fAkVfn8iz7Tjq3vmD3YhliAEZmZXC6yId3PgyoFoteM/og9ngT
PxDtOu/aPDWTUQjT470E/xAdxN8Ez+YNOrIjfb0lrDyho13PU151vte+qN6l91ao1sXduQwHBsF+
oo4XqSS4PM3Dm6RafqFkFYhiS8OIWNeyzwRmWhjff+soA1E5REv9Yvky9oiZEk0KjwoueTkrG6w7
Tp5ZtKArIRfJ8qx/tx8GNvF9xOghQ6QrpwdY0liLlE2yIlJfUkvnmQ3uz7QJQ0tKMDXlX9E2lqlv
3IOV4lXrhoF//su3IJ0EadqpQ0iBXVDdotTPH/bqZIjEzysP7KlRJa2VUyqnWJy+QuQq7qAx5kn/
2qZ68ykIDZBD20vqPw4tTcK0Ay4JksilEEIJySYHCe/d1SgviECZstOW8wp1loiNYWfOU2SRl78w
S7nMnPWDQBjaQQjd0tRXSx+VIIT9AG4VGUk31MSsr/pA1iPjYEYThQ3l/qJg0JRJ4PLTHtJNR8xM
pSRGUXj1rdGFFLwo90DuyrG4735aKrWvxTVXTY8ia7sc+btF1q9Jzy2pSCtjmUDHNa0hW6vPEXON
LwB5m56vNrvDnz2uSHI1wclhfvWodSxSImsmjhezu6mndgnLg0ozHI8C9YHH1mAW5vo+o8Zc9nDL
wb0zpz+np0gOvBSkhxWNAZ2frKp8fJsWbZOVCnWXJvDlXCoMSBFYd6rR5eDA5cAEAyiwMag2946O
O7T8Moy1sHDBNv4a50IzvRZ+qpQrhYtej7xYzWX5fF5w03VvtZpUkloyuq51reFsgjQmlAINv9rY
kXad0yNE5BJDQT9PJoImX3rD2CTZF6Zb+Y2cO/9wY+I1Lo95twOPMTZp3UQVNYPbCneaK8FokQI2
iDhPKSmYruV3moY/38XFvGNys1yJ+k9+Vyn65cJgXxzi/YCBAF/+8FYIfGRgLgeIJIqTXEjToVxf
XTJyj5RJqGwcuk+sEqN5b96zB4SkQv8LauomJ5pjuc6cSVYIvic1REZMTXIz/jMoXvs5nDmpJh7J
udWE8epquqg2uEPlhlcoMXthglFdSQmtdOeE4aLf6SXBeFgK92fkSzLnmdJqnh2ehPb5iHDUpmPZ
xc19GCln74fAhERJ2S/HNBKS/E73qedf5O/zfhJoKPvtjr/wxaNMjC+rNhGJUyS/sSZPuMV8NdJk
rrm6HbxsRd3nY+l8JpVcHloSLyCSHmqA3lK42MgXAb5Y6UZXVawlvAYgWJISJEy824uUpRC1sv7Y
gSzbHBkWKJ6fwqAvO0LTsCGZ2165Omrn9NRpNzATTHnNAD85LEJCzBej4TLBqJCDgS28tlnJnBY3
UNoV16rCv3SQD9N4ByTKYgDM+JKn0+pMUsFDFbbXvZsxOKO0l1TyLahN/EcwVha8fDTUtESLK7It
+cMERCkvRmtmmw6fyN+WlsVykBgStYq7+9dOhW7vHN28/O8l9rXgcmasuNQUkJYCylSlkdOTJXEI
MTT/qG6dNQ8Szv/0kg3fist3cma/dY5pu4PMKULVJyo9iMDLB/F2uap6RWNG73ck7NYDbwmH8/hb
rT8apXE+K8hU/TqIV7FRBZe8oXwz6xXllhhPB2HhIQi54QxvdQ7o6oOh8jBs1GYWuA5Xgv570jQ3
5F0WbvvAQeYwTbXVbgPOofG+cz1O9M9UYDjIXshtianKWI19+09tltazwo/iENGEqaxYYXwNKOMO
ofC0KaOiRA+965qqRnVcnj8LXBJKZiK0dk1wJlPqnP6idMzwsa6TVyr73RZq4nKi9q8JgTbOUnMj
CBuCAt+mTbqMTF9MzHbMaKwxPuC1jO+4cUkGpV3x49vSk6t3SdpOS4CPtzGU7qCNq9gQKjtDq+Nu
9deJ1FyQvNIIl4clawo5R2mgZV1pvLRA7IjZR3+6cCli8MuXg8RG3qyfs/uDu37tKeL9UA/raTb6
S9/J8nOaGPd025aWwqsVjjqGfhDKhHmNnBRr32N0AaqvrEfmxPqnuWNYrlzyuXjPxaVMvbxwN/Yu
D1BI0mWiyUYG/qEyc1bBeF/SR5NP/KH75mvlURIDK0hQ6fJgISFawD1AHENyivVhX5VgEbfUkJ+J
QKe6bwjtFsrJevYIWAkGbKcXKz6QmdtfMbkGTNbrdp61nz21+N//u/tfUbJFn2aMVSRBb0aiPkQ6
bzy37Xw9GAj0rmb9DSTcV4Fgx5Sjm3TwEqKuElMVn6jQiw7mHG5QgbZgAj6ahhbgbFmczeam+aK5
6jlMD5byvZ3Gi7h9GWaaECZRL9aAjcnZKFZnpk8p9yfwzBTSfFLC7jCgs+lsoCPCky7+O2A7wOzC
z8/CA6ufNpIejyeLLmaj3bVQAfXiJDbP7tTioin/4YvjjuLpb9d6d99ASKkhwtqyFyW16f8Q7oL2
Ji2csiWH+aBqqi7gKXoAbiUz5sJGWtS888lCQpUoU7EsUoTqAdniu1gKQ8AtUODRzbn9i0qiuLCJ
hXCe11m4TiN64lAjy31fiLP2D1N6PaId3j6z09moBxGE9vs0HnCcAhXqxPKrExv7rF0XY7Fdz0LO
s2LwGvmz7Z7TkFoZ5v/ehJb2fzd0zrMl1AcLLlEGffzcLmLWp3Ahq3MAOGagUSnHR1kMEXTpNPnA
RKt6q9CNzp4LQXcnz2YBr6Ro+g5sqKzp7sym/qx72GRfPStSgNr9hPirXMMJtMJ1PJd2vhXcMdKX
S4Zld+q+KX7p2875qmqegwkrdDFbA8xuuKZ1CTP+2Z+AsP3CCd55lulMC8OMXnkTA+Y5XRzkLfLB
BV9rpuFE2rJXOcYTKW3vYYuKNNPeZNC/XjjIjzJBihe9y+YdCWpdxGfZ3ZBYbS/m8YQzX4KZ8k8a
oVqkyNBH79+vlIzm4ArXVl0wc3653+lo1q7RDRugCLA+Y8xWG0yci3Nb9xDwrllEuFqlrP3v3xpG
yMO6sxlIR3Mpy53miXThOzFqGEXo/U6RK2KLEZxSBtTb5Ywb4cJCaG2zMPzoGDHysNcJv79AH52Q
/4xGQzN6L1BanHDRZ8Ee9lKCmkdsyS1bLd9NjW6Wdh0+xVh4En4aMh16XQgm99YoAOL3F/Gll9Dx
jQur0DG8rTYnBo6h/0oTZ2ZoKLYbCt1a6FF7SFXvGeH/7QOyDYCXm0E36t1sKMQAIP5ISxfepSB3
CGxX8av2q6Y+q09g3OvG9vKshZBP1vUAE1yL/sE3tdyKzY2NmVH4TY92RAmzJ5v+mOrH7FN4C+Fu
FlzqVQiEm+HNtjtyP9oKtCrYAEc7oi3a89z+xQf1Fk/Ms/kbaC7UdJtamtQH83sKBDvv8f7fFhsn
4P0mNjKTePaG5r/61oOMVI5JlomzPd6cBhcf2PqDKYIl5WVLESC8Q4o6Wl5pjvUBzKb/JgvZFWnR
ZcE2DKT/j+O+OWRABYxT4/BMH12mQOFWl/4DAZxhYeJ4TQZ+GxM8TVsnqlTBmVqCLoy7sDSpHK2h
YXunNJTezjtOeq7RG6ylCxPyrzRKkRGCtmpGHxF0MeziV20iO6EOrFv7ThyILb4KHRIKn1IXFaLA
idNXzACDidYxC3B5Q7bnF7bHET6B8JAUfaCSAQfuCzpfS+c38jwhjYdPD9Sq1cA2DPzivjS3lnEr
ZjlNSBc7BIuFPYgDzP47zpF+1sxjbSVb7SayG2gQt66XuBtOk3lWK/wsA47b5o96RPJRey2GgcHE
aAUzrKQ5L4uH+YbXbFjM+xNwTx/HF+CDhDynKlbt67g3tvH6cET4S5Z1S3HfZ1+C7d/Xg/gxrP51
4icGE5jT2NZaE5a57JMVe1UUKXUIMegw7C94PHr7zfuPLZL+skfl7/YShM+XcfPaxIIdTh2nXF+3
9wngczXq+H2GXLBdpsfS3/Gvz20MO+YTedcSEjyTuRhvEVyXnB0spHzLr/1IGBwicVr4h2AycTsH
VUsQzZnuDXiVRRNo74gxkXStQ0sQm3NiJQLbyOWeaojdSlS4+KlUjzGn6ATwKt/NLW5BgyzMQn1O
Z8eFLGkx3/BJWEHxBPphOeJ1VkMQWcLc18AhXADhsHBzwRX5M0XTWv0RuHVXJz5iI/7rnajc4JQ/
AdwLcTQhyQF3JU+gnU5XNx5AstPY6FCHSb3+gE2U1IOFr4kk/MHIavt7+qu2x8jbo0LVcZR19V2K
mmHICYwWwj48FoMSlmch2KgKO3aLpNxvqw6PaLUqoyurYWXLa+ZYZxP4W3T2e2XnWAjJb/Q0q91k
EWrEkbAFh+3L0avg9PeMEN8LDNn/Tdr4w4MWwNk6s2xh6DNelb2ReoP/TBTXNi/ZrpGJDJUX16ZY
FwT46COQuPtHPx5StYfaJxc5EY2mC2lterTbdugiCpZuz8EVYOS98SgI+duXD8Bj7HG/TmY2JEZK
LJDd+iaag/Njd8derzPBSzs2EURQkOU1h5po/SxD20Q5rR1lE4X3DMz7TVxjgNl3FFphYJCZTj1p
jrtxHxRZhKZ8zWgvk4SOYCD4PDRkqZ87oy+EmQcyrngPtHrCc6o//rGbb1p3iu/9Nl49jLyLFbyg
Z2BSdEe9I/dsykfH0KUaQGfywgTdzj9lHIyftY5x0/gWO9AfjKTcyScHNnG5vcruyLyANnCiTFo2
2zgCr+SrX7cuj6KUcmJhENEHDoRtTHBn7ZUX9K6F2htHF//y9EkolKHdvnW4O/Zxh7sk7GUtUJfG
Jo7vxBH2g/O9dnIdcbMTQuIp6UpDtlCTYslkqwkKAjLlLUPXpqz6Uos5thkGyQ14IuGInesVrdNf
ahMMd9X2/2znaYXPdOAkLI0YoHR6QnG9rmGLfkFtEMGXGwOESBpX9RwVGbqSmRqNpMOFkAr+F0Ul
DexWpSRe2XsEF6MK0eveDaT/2tZnSZSVwRfIAT+RfociFG42eiKUfRMDnUzEIe9Z8FCY1Dv1Nq59
3jQMyfJGkxiVgkc8BccJmkCQjqXYAtupiRCuvthNxx75j3EmXQxg/d89myE7ji+hk3s/S0a48GrA
/PRlLuCKuL8t5Ru3coZ35cE8hTg9lmmcMCXOOU77ahKtIRHhqBL5h4NftVWfkZcTIWbZsznhaZVZ
8cBa+RiuotZpBEFdZGgLvF+8ZBWJ1s8MJOqvq5Ax5QaA1tdbny8nP1gI9TLxwTJvVSglmfberiCm
h0x6waVH/KHWuaJab+sfh5FPUclEJgWYB+QpLPf+AXjt1eQm82g8SUPpVGAPv5LowCy/E0O0wmS3
/FNFMSnYjhpQj9gWrlFqtTDreg2ysG1NvX2HDPBXFAiX6zrh81yjaEAFVpuwI6ncwPO7GYzQyKFN
Vj2lP5tTuSm+FQ3U6OC5iVc2LpMOvQKRpX65YbSwyxPkY4ER2eAqq0fB7PxdCUYSN/uu4xjEkAxR
H0tsd59NpZZ0i5jzoxDOBTLl6mTDu4D/6a8PNjWOXXW6xjcvTWBJ7hCpVhfUhHV+z4PJr8+QaqMB
voM1MfBgC+hvR1F+7hIJuRmuO0uS+GmpT3P4KfE1ARyHWKTwuVSFdZyTH3oZXdz411D16JTO30ul
Y7gdsAZS29lIGW7BYLSGXmWT/iFWN0HmkaHNF1oz/BFxS2Tit00sod0gQaOdKuKu3z49oswphrQO
JejsT4AylfBfevKQpF/E0ScPmvmxR4c9HnwY7Ls69TEHbhA1RIB0oOC8WP7AvJKivoLh2dZ/0EI4
50SA/FTxx4IL/C4rCppf/eRzUritbd6K6ww3iiLAj3dt0Nlu8sIpCCPf/g6GVM43lN+enQ5nhGHF
2C6CQV0BGS46Q88DfHt8YvGaNS6DsTt4VMU5Vy5LdjGTHe6BctrMxAK7cwfU7iruvSIcoXskp8PD
gqQuX5RS1sgAtcJaAvExtb92DdkT5skgEJkZJrPyYPPUD2UUG1sahfXisQbfLvVza9nZ6mVThuf2
Ug5WhRVsJzYYgqwIauqDN2hjXAwyXfsz1z47Qk/rGHgdeLrSIFJ+FIndWATrXBVQi2iKnuK51ErD
O8c91Hh7Z1TBf149HpYWarzQA90d+TmmgtqqAEw9Dk5yDWAvg1YXMgokutGMjUF8pOhHEfOtHRVZ
F/f6cUwxDwB99UQ5R1rCzGctz/IAn9xYMFuFrrQLRkh+lNWPuYYbGi1ajbMkmxTCkS9oKlBz05lT
GEigT5iHsJ/wkZdXoQGd/VoABrmvxQyenj00m8tq9cdR7LzKiRQPQBMPAgT9wQD8r7vKH8cRNGhx
4X1ZtiXFpfNPXK9QL/3Pt956qzyOBeSc/0q99I0/hQ8QNXgWVbbhwufZ9aFcG1kqGw6aBipOslvf
qnAmgimPX7cwAg3xOkHq1tosLpZbKTXt0OL1ZuA7pLjw541C64j8xtYkhQREbaCQlVfryCvqVvQN
i3AMLKmGlE7Uqx6+Z+3x8SPiZZdHDu8lflOj/FIE0pGTGSbx44nQvXXM//d6xFm5R+TC0lgek3Kx
W7dL5aboK+4WU8sqV+0iR7ivcnTwYlnaWCd0N/4RJ7Hk7ylLpv2//PRDmiP4Bk9nw8N981ZU7cXo
aR+NAs7newQAtsrWBUuDjpvoRK9PzxehIkUCr3J8oVdsSb7eFbGJe69OJU4gbK+ZvaNF1JzUIW2f
0YegfplP2hdu/t/14JX6N7fh8LkYysENmodF0RmD34cwreuzTClkYu5xN5ren8ZfHzJJB+3Hu5uT
H0CGsRfyVjaaUFif/Oo/CbzSKeXTrzLHujw7yKb25qmzBA2tRwYnA+z5aU66fm5eKpssJQ29G2HG
52WIgzSrVbJXuSAWferKSmOMI4tAg+u+g2niVc4eHBuS/xGXRdm5BVFAchuS9b+njgX/4ouFW8y5
JrPr9L4ExzOVu8VxiczdJjXJXimuoiERRmKAUHXNPwmyY0Tx7icJ7t6p+IsIS1R8XhvqJokNBbOt
f6vTyeDxpnnpFvEy3vFvGaVaED7oLX2v/1UHb4T/laUbko1vb5YNpJJsrYpofGIvGX9IRfddKXS/
jjxHD23dHgv2FQyvJBoWhzLDPEhBPY1CMsQCedryxTY+OcPlCv4vdr8ZZ77MeSg3+SV8rXZHHhKO
yH8J+c4P1vFR4k8CNegxo3Y1w1mKJxDiz4qfcUhPPI4wiI7VPsQJn6WzDzbc1oeiY93c8U08NNEU
3S5jhzqEpvMKmRkq2i7QH71nJ9RowQdjU4Z8DhFankU2k7dYBmKlGEPd7y4H3Ni1gQMMpEEAq/yv
erdsnNAq5WpFK0hXedviW7kA/0m+c17HLTkK2DLDfGUUC6rysCroZLO1RZ1In7buj5VwAfc90cNg
4GD8eXNHmUdUCX+zroZ1ul3hHSPql124+PsEBlS0fi2nRdpSKMu4EuW6HdB8pMs5SWeJwRDpC6zY
eL6CMOFXkNg+M1I64dsoyLDobY/Qx+paMcKd1PBfGbUj048kvkBI3IFwzmw3tj5pa6Fa5u2JBzIK
V7PhPOBn3VTbuGKBbC1dZxCxvAm8ODRwFvjAvp+3ZGCmDudk2z3Za97wdCH5+P3HfzPPEt2S273E
5evjO94GupYBzbBWo0k3fAJ/c1Vb3yWa4ymTGPAwPmMtTIpCO6Qxhx3DOg06VP2nFv/lZdC5U17w
8gD95rDhxY0TFteEmnrT3E58UPy4MaDyr0938bNSbl0il7K6XsUHCypExSgD3gwSzVv5NTR/gdgy
5rWi7jnzIXRqyYXuKkddZCldT0VDrURZxQOGpCCCSZuBZewLq2fGHtcZwM4XHV8T6BF5y55fR8iJ
aWr7LMLYIziaPwadJ+wrKj7k8jFT7sYmkVDW7o0ZcjAwRr9kcJT4LOp7k9F5vk8iJMw7kue6DU4e
PMRud29YT/b5fecMUfwuq5yjZBMj+KuHb66bStWh4zxwAPtpQt9SEtK0qsteT/175CwRmc1FSF/7
clMNPA10fL28YmumBTCzGG/v/eDwmykiqtYBXnAG56aOubGgwl6O4DGg5tnozrI3CRtPiU6lW18Y
jGDJ0md/7xY/7UZ6frq8mOxuw/sIwB74f+sY+6kYlXiCgt7vZxrv+6m8UTtD+EkwA1NjD+Ug3Kug
YfolJGM2SJgGbVQKy31aPfsoiMyjGbIc+47h9u8r14Liw+X1BiTsvSbOL2Zr6imMnaNoGnNt4eCc
76v0rtrKMzZu59Et4VUl9o4zszjExHdlH5ETDDgDdBmtgDdVQuoBoke+7IbSxeyJsCZx/SbZXIu1
mPkhaPNGArfYVIr3oNwd8TOwGI0AR6bKkpFAhfyI2cKMf8uJEUDOJhmj/6Z/3FJFonLP1n9qylPX
a1zXe9m8DBPUFE0jwkAGbMFxpTzDWpGCOGNGXkZaygjSh8ua8hW4KgB3MVQaCMzovpIbz7KKELk0
kuyHsU+X0m39fJuh2K4scG81tYOki/ldXg++JGfPVDXcx0nf7i7BkaP5Wz09VEAV6xPd2v+cfhgY
/wB8/Ui7/Uv7+KDIT2Z3gfJudXTJrkqtWQJraANg7XzZqQF5C1QUgkSDwUq63MsWYpl+oN25fEpH
Foa2L+b/OjSdGFKyQCb7/iSCeEJBr9UtvGh7UKKBVzifiknWB6z/oCpek91tpSChnhdVwYLeGvm+
xxS3C9n0M62jvQbjuCz9S22FF9iHZEAfaYORxojhfsozb9uIeSJZNgiNpC0ROfvEpe5AlxJbJfSV
EMFTuLsECz3Oqg0UlrBUaVEsxNeUYYbKzuK6mKke/eZWZAmAAQQ+j3jhHRMqEHxVIp5uhPkFONNZ
sOf7CNQFRFNCWFNcyyjDdeK7rFWg97doAWhGemn78hn/H2qFfEaLVULEbLum82i28cWhhQABgAT4
br3wjZM+Rc4HXQ/lVAma/vYTJ1y2agBgsnLRkoNc6j0iaM/OwgwtR86CcsCHbyyHa5YZ40HWMPmt
vl8C9j6fslD/jOZIggcKXt8XOlmK7t2AbeZB9KQO5aZkNsnJxcIpApWAeprlIjYsiQfYOcT5P0OL
d45Tfz6V5jqRoJFNgvLuvjQivhw8Sx9KmeYP0Moq4+E1dPH5OBxHySiec+1E71VEwocLeOnv283C
s5vqlUKMDxz0viAwL5f9n6+0eGi/oRW0pYpPONVBFJmKNXMvabnKCrJ6+UFJx+6ZLC9AbQySBs3G
hM6KJ1k8fv/SOmUfJKT2CY8ShSOFR3eMR7aVNsOgYTrvsnRr0C57bC/T2X1oG1D9cfVTGgyb586C
0TvPs7u7uhrtK7DJU2cuS0lAB/kNj2rGbmiASa/HwN/9CNDIZiBC5orj1QKMOp8M4szpFQGs+YFm
oYAIQcpgZtcRK5/9GolLBmmo7+8toUBSoZHkY/Ig0NZUWyCNOZ0ZciOwdBt//rLxriD1gkr/TWxn
coBBdPaLjjIj0ydvvnZoEIxcqirI+9HKlzXVGJwrobxRA1mZeHhoNtR8Q90KrRV3ScdnKjfbvSzp
L4yEf1hw+aP+hWOUeIVjaxh8n0gjBOshhrMp02hT2NM3L/3RCt++ae5obEAEKGPI0LQSkGV8n0c4
zButMFeCYw5FQBjpKcaImE8t4NBft0gAbgTOxwLcXa8PxN15zT89bZcJVU38pOrb06XkbHTq6I80
pxoBIBWZFytklq77espVVuRk+V6W05RrXmuWB0voKu/gnqdBf0852ssn6n3yVJ4sNxkIXUl2XElU
jctoMi3GsGOjHqOjFyLeW7tkblpF+hKtr3U+y2jZPwbg7HqrgyAqZRHtxGvZoMixUO4Y/MMrB+/c
eGh1NMZH4YT3adt70xaxoULQ3w84TuvQCqB9wX7X+0ZVyuli0rO07DOl/UyOXXwOEbIxkdDK5TXA
eKPRON9zAmKSH44D/hkTGm8u20lwEd8+8DBCx/U/Y8uvzJ4CeASaEBOaxbXrkkiEJo8U0ql4e7/Q
rLt07wU3EURiaRfcjcjOheeElRTRTsfcvXemwr/MRatrGYtSrPFfkzSRU8Xzgle1t9ZhQ8umNhk8
tY42QCxiwEzMNuozSRktGGtZs13fRHCmI892287vLCuHVCHcW0vtbjVzlad7QodFZPnv6ci1sPz6
WMmxdI9hlpld+yzZncgCcnRD5mfqCg5ExMIqyHt7tfZyt4gKd2EEeA0lc0MCgre53B/uQLyVUq3a
cjUpb2YC7ykBLbnmWzuQJWptOnVZvrhCcvlq5kqpCGI+2hEck3MoeqjH2pVYm2UPs2s1BD0aMduu
LgG0OQSUfn9FecwTI1vGbVcUHMZpX9UAymieDGJHsTQlVwcfaVUEjgbJXXdIEAZrptLjbEnEUrix
IryFyFuzxFhNSfwGSeRF80OXvpYUlDFAyA4jrc5HcrSVkUDhnzys1t1ETTEhDzVkSAjypiFjBQrd
FspseTZNJAXAaueVocV25uHniOqw96DSl3ZYL/36mkHbpDo/m8gWzPNvW7edCJ6QmAMMi9VEK46f
ULDKfNMCcrlWdAAABo1kMgDSWgM9tuP5l3F5iRaC0zHMg0H+WNYh+uGUK37yBXrB/Dw/g9L3tYO8
cV8NzpzXP6QZLY57BT5TYF+cL7LOG+wtOm11+9VxCOe2Osj+XekoBSRN7TRv1Nytt4W0EgSWoiF2
G/4SNM69rasg9zbZnNodxSayViwND6OPiQBJVZekgML0hWWL3ayNFO7ne+lcrrJZnZmqCjzhmmoI
BSnL7KQm9koPgVhctv0z4qQyDhPqEkyCgJdk6syuXFjIsWn4rpLYzCMmW7fdViGZ6LnKjD3aElXw
s8qBKWw2wyneKYtovpH03lciYajtoKiEMNWoZkryUL5VquotCdEfxh/u2YOUFQclv9SP7/jr6iMV
b9RoLTHNEQL+L1VmkAoeMqfOubvegHf8o4phL3iuVfYWCwcS6EdB5YZWJCst5Mpr9Apkj2uj0bVs
n+j3TU4OmVadsFOR+eyCSvteEmLecUtAGJ4MjrVT3Lqzbacue2mD7XoGFgvQB2bg1JbyAXpis7bt
e9VmGWS+DTKpkI8q5G5W8LJJOuPcUSQsF8qSnTANSBESe9HrAuaUr8GOJ5hU+RcuQVfDCYEe/wzg
HdhBUAY9lK1mjK8javMvZZ8jqWA42Tl7Xg==
`pragma protect end_protected
