`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
EOo+OV15qPDCNbtm5oSy57JVGmqEcsDIZYhpqQAEnnEZdtZNjeJbDKGI5ExMT+MomRwakuHoOzuj
nl3B07w6ag==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IVyvSBy8s5ePNcOsTboCjC6nA4htNoBygSYxgJwPBrFrBtdZzZFNR0x55LAtJ4Bv7gih05dhU7BD
sKQq+MIA54XtRKk0UFPOBTL+WRqE9AQ5XfthENit20ovG/Dd9XC/FOpmsqqTLHVkQzwMBplqDwzC
f+GNBTL5+swMUtZphT8=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
uusZIhvdY43/hVpa3nJS8HYRDFDDyrct69SIa6rD9DyKAHDTJj908z+6yJVrg30FYqu0NyJkzG0t
e5pmKS34UqFTJYpMHIVmubUQbkCQGgJZ/gRxEOyXUtcJfEhpWWHIdfsGIIvyvVo4PCtiq0iL7iRg
XNcHhDAi6NiCTEmdYWrRPNCTNBq24B+l0zRySkxc43V05s0LzXMoqw3OgSlWWQrtuLdvPKCCxEWK
HdbB/8kdFZXzuNnezEapTeeVYb31qpZ8WdST5OOfSiIjDOvZAREgvrFGtXqwhyKvYKTGY7np/7Bd
JSWR9FftD3IgkkXQhuPT0itGRU3mIrJLKgPVEw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
S5Zl80jcHElasaEZbOhSe8t4Pc1ge1rFqBX8dE/GiHBsqZCFIp2f6KBxOfSmeP2z32ERKc95de2B
ArU+VMfFkI3In65T7d6dE0zgEY5xFvjUekZRhoJBB+c8VXFopg6rn0Kb2gWxFeUB5eOMXHGoCu3T
pfdaRy3fHtWupkbVQzaICbAY9GkqlWRdtYYwENFa67M6DOYvsdFlnlowpu6WotlOBJWNb7s/A5NC
nlawnUMlpopehiukxgpv9mVUyFpqeY3G3CJjQhRWF7skQmoK0c3FbWwExWJjww59kC3F1vtfG/O/
+vbU5o8i9k+myT96+Eol89a8bfGRMRCI8+vKEQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KpZr1Q/1Ci2aNd5h6/UbX/cNRPTq0i67JrJUlfhcoClVqm8Z4TS8EgDvO7jYiJvbaBJmmWNMLxV5
cZAAO+44ouXFA/uUK5aN3oA9LmmH0wfDpnvubICiCFTFfZmP/X7fMgqPgyZn0WGaeIThIHJKJ4ya
Qray78YicX+UEwZj9rg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HaBLux0ndD4Nz9rgtXwh2LRdlzuWRm/gnVVuiI1G4VPpL29oCgAGdp1JZgIJ0StwP+5kPsihvlPp
N9iwO1a+zFeIm0spM+uRn7YhCn+Uu262FfrVkIOx3EChVBk+v/i7/ycjSvPWSahLpJ6QX37hIqRp
8U2d4PrjUkZ3Q6AjRX83ITX1C8zX0gmP1jQwNmbMnQU8EPzAZSxVC5D6VC76yd3SbKJ/HFaPW6RB
/tTB/EOy2eEwtOV73MC18qa7v0iZTtZYvmiVdpFX61uLxxJPbig6LZg5MIsZCK/23zSuMxt2LGUC
xvFdoOg61T58rIMXr3iK8iu/uopflJ4EtCtzqQ==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
q0ZeP+16wqkVpWynebloQ00OdqCbOxlWC/uwIPMFnd+5Rkz7smohiVvzLdfQvDy6QUtckDSdDMx/
MuigsrTACEs9O+LrPFNINiKvF93U43im7VNa8ZcruDGR8vODQq4ldmNZ+LZBBaW6NEXaB7ngiY6g
P545lyMT+MiNiFZz+RNvVhA1su25M96zzrwYMuZPLnbF2Y288eoYTGgqH34suISLMW+2a0uwA0d5
2BM4J7gHau2mppX1B46czp+VliUoGrXaOWalLMoj6OPUXXkDkKUZgubbFb0WIaVHR/1lr5R0e1aQ
60o1AMBW0ySOsDQ9Qull81JwiMDovICmUA1xCQ==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RvpW0zvS8QTll7PgbpJAkF2QgOJGQNG4c6m77E4XkF3uAk4vlcMxPkHVXfVsBA7yqhhIZkUg7/x3
Mhh/NjGHoYxjpB2d4Utacjf1Seunr6UE+bbXM5QhG0iYUuQfJq1P47HA9h/eYB57YknHsW4Uh35n
VKCGR6ZAxSfYTfdjnwUTaeG9ntyXOFjpZFXiOrKKOcnJFW7gtMvLEXULc9ezP7oIWpIK07ZhUl6f
m+K2t6KAoo2ziAXRHMJv4EK1H5NWvGMImLFDSME0dfaSd1peg1LBKSHnGR66jB0jTSk7cjpbzcS7
fSUU8p5dFT/pini/3bFtHj0szA7+m6rL+C3rNw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TRrl1CpzejkAq5QsR2lusda1NqatL7vENjpF500mzaz2/zkBy8hBCkLlG++yN2oaFAj08Gp8sZ1j
LCHAQVZ4FZ1TgbPiEaMYEtUxyeCKkpUEPb7IsbbxEiXdJ0V81pi4idIbxVkfS4uhaglon+8121Bk
y8DSIENlehWPt1e2BaWLjCo1nPxFKOwebaWulMO4oZrRXlYjwCZao4WUofPV2sABjYwRR3WOczcg
/7N5FWHT+RNr++OxJjIpiUWHz5hmgZYVIoyi53lo3qRtLyFF8sCtKdYVB4bKvNqCIv0BX303v2G0
ey7yFVQ1jJ9YdyAysOhjklN11oxcqKd1fzxMPg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432)
`pragma protect data_block
d6hhPoOQiqhOkVpEZZzn1NjeK6BZtnfWoSEj7NfEYQJJPQQorQbCwFDe1edvvd+FLyQ2MXDkU/YP
SY1ogvoqEtUtpIsZISYT/paxlgx3qqNPukhPwnzzTA/0lBPwr9cKlz67sxd29wGMg37zqjuS57Py
IDiL/J1l8imCdoGreUK2w1QcbzoReZXJOVMa8NQkgyls/M9F6JRzHEdQzBMg7eM/F6f1A/XzvNVT
f6nYArjTrKfjDtFhq4abpZxeZu4AXeCok3mI9vQQxbqYbb9zBACT1kZHAfdIo2fKZZ2mOgGSTAYY
96Q0AfUL+wAgb/WHSVkavgIeMXqsGsr3exzyLe3p+0K3N2pzFiIuq9eDUOrWcihNsnzXOx6v9MmP
UV6z1z2E5sfoHv8Dtq/dwsKWuHVW8Hta5GMFgujqdPXXbHjxmmy0wv1n9QW9v7xGzarGUU+b4KAs
XKlt9YXcq0hkgfRTBj14IKEY1r8CUxJopHiVYDAWqI8FIGQA115CUAOg0QAoL6hDwwMHuLYW0U//
dHvVkedKdwVuBiBZU5x+J4HIjiP8AalVZrg6D3cGOOrR
`pragma protect end_protected
