`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 78688)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCWkq9Q7sGKUfekyOUZQK4PRcosgQmmcCzsxuTnFB3d7s6toQeIIuciug
Q0f+emK30TdB91wsQZSjuTAIoNWYKRzulmWs/bNsWh72Usw34oZuM18r/NXqk/zyOpOYqDbkKl+d
JK7fcaF2pPPBhs4212VhL/lYQPvWX4HAzOgKKEY499gTTkeUYoqXvDWK3UD4QOPk0ehmPUjD0tn3
Sob3GTzCPy6690TRlsERv265vgqCMPNrXSdlhP7G7V4VjF9U6pFpSM9NjV77F1yaUskIk+Jl0BqQ
DNeLfxnpF6OaTpN1JAPqtkKvHvgzjOQlCvr03Bd1Tdkf4wZirfn/qDXkUTJif2prfzfT9eGtsIyq
WM2FGMtpLPycBXi6H2MjOTZKL3ohr3j4855brMkHIiWWhn0cyWHSfCS3LeuCFCrfRWO22df37B8m
kxgeHYAPYxHcOflG7ot5Z48yCjpRnVeJ4y8bO20URqyph5+9vNrJdbUY2XFfm8EDYkpl88MzBNGw
Q2I/L4hn8sCU3jX36ZSjzNl/MCMUrSzRutzRFMbn1YbqSACIQVETa10K3Zb6vw6yzBAvfY5vVIwi
5CVTV85F3S6hUK9Cv7juxqppiM4sr5CQAsP/b8rWwiRcXIVf35oT039UqoOmj3j3ybepui1xrDhz
Z8PrrhUkou0Gpb/MiIIzJYHKRWacodBLAVzD/UaaLlWFpqmCGlK2V6Jka+iFCXAAbyPpZSdcOj6l
43jwjVAu/bRrnj29w3sHYqlmtCb7uhlTIE92kUHXUhHHPcxrA+giqpht2zrno7Mx7Z86vS05aPZJ
vRQjTBULq5AwWZWKLPZQk0Lx3XFzvLX36L9HxacUddpr6UATiyffXBL/m4ksa08I9yxbzqSShjO3
ibTONn6Or6oha10lZ00wRUtze4Z0lLPMlXk/AmRgVYoIXcQDAy4qT0hcW6iQ8we2cM1CTIQyXCVZ
DVZhDSSRtw/4mJArDSa5ehsFGcL6biKQlZD2bGqjXHmWdtsHPU0Mo2xQDos7cdAk17iBLZ9wkuOC
aJ7UWe8nVUFwYXGFO3EiMQUJzx1j+hVeUWRZWR7XGfTCle1sUh+9pTMmfuRnBcd1hlgWNm+vzgOx
bH1u5gNVbzT3W0W3/KmUHl68rJyRZW0QlR+eaMv+mohMMjW5ik5zuDZa92SofPt4yzyJrRRn0bZ3
zrEJrwXUY2d41+EDCZ+X67GvV7QQlUaL3bRe6Mx1XW270vU/IY1hDE5llPoam6IEoypbEGtavVau
175hVtIaDotZY5Cl1SQ4ZCtACs57jrK/r5bf3bGinhkD0RarGtizLm2/hzojHf0b5gnu3F8XikUT
dKsukQLN8c6P3lKj9arodvx09L/2an/UhAIkoJW7zBdAE458z0FCzxJbhtK9FiapbZmvORmX0xRj
WAkTvezlJy94BoJs+vYD75VTw8YfGFOO4JKP2/T2TM5PwdtRyrNSLKPVtIbwrXMBdYyqU+1vB72r
ua+zXIurXnA4jOYQ5PQ+XG83NVQIniXhHj6QuZEhlxuaCixfPc2TMrqq3zi4Rg/bkXiC6ttqaO7j
4DDK3uKiqFYELF/u6aMQWhd6FyFMuk//050DkXh4Pt6CyISfK3T/KqgQPRD29WWPFaZ/8egnu7pe
3UruRWn+wAH1bF4N6C5lYg+7e/YsMQu1HSeXcbap4OjOwD0GW4LfVrWzzwtdYuvId+rnFBG4MqMz
sOWK3APk9p/GfUKnvDFUIw2mO5nWRcqse6Egwk29ZMXKVUoO8KmyjYDPTsNwBDqHZsR1m1p0jzOV
SFmJpn/+MiUQZKjy32kinY8EwNxxWfKcafUn/08eGmWOpwSkx2wyXmm6kE61/3nCVb2IKFBa4o8f
mE5cMJWOY0EnAuc48xcyCqXW0aup4EGGTHrzq11RGXy7+JYCwSGEnl9IkmOOCuFxVc3G4x3A7o4t
+NbDgkCKmxdi9G+g4yeD9CRy608xCbHO0VSrKAxKBCIQZtdOy9m9P4r/G3L0gCKv/j25lhZhFTsp
6sfttQe3sYRSdCWU0HA3y0lbsSqdfsUu2enMvQuEEltgJSq2OnxMzjXTyZCXst2TcG4L6rmXyOZn
9o2DlKYvV6GRDKrRsixtz/JlmOS2WourJe01XUQBZ6uGFFFIE7JmjxjmfRj0BIlTW6ucZk2qk84B
Rid6xpQzmjYpJRiwDZmq9K6u6O3CGK8acAzTEGzd/kIXT+NxMcl7zguCoCyRCzulj35hi5g2atK+
M6mfyUuV0YAM+ceyxU2L8RJNU1emhx6pw9nTprEJWTZwKWc75VMpvTxD4Pn07ZVOxBErmn/fo+cY
FFJiRgcF66TjW2Q5VZdwQtsov9G+FP1deUumFBX3byzQ7KPNnDcPzjExRUvRmnlsk9F7ChILAfaq
Zo5F5qGhnjzlOZZX/6rZUDV+ETJPRFnKGzPzF7DjRh9Wu+iBEsOeWYyKNOjZ7npSjIwAWUY5C9S7
kmzti2LMrnuhMDy8zEhzkJacI9ejn9X6lQnLeSH/NiHERjG0l/56OPDC7q46Gvdhpymvm9wodfrt
RMNddqLRl0X28fJ7d2h3LXcglWyJuJqPWQB+taq8la4rmbqSBljf/cMxaXVsg8B12pN8EQXOdFWb
+j8JxTLEppEXRlUiwX9MHSz6LZCQ9Av5vsSwIzwVGAF56eTZeKLnWC4dhvvon17qfUBzD9U+DLMc
cYfh7r0i61bQPmlX+8Hmw034QQeGaZagb9qhcyRnrXwnSBwAmj+wTULRdCshqLbGJ8VgfYR99fDN
VIzD1+4ARkzTFvS3DRkD333R3bhujh3Mx478t5wRF1Rgf6h/yQPc0ociRHBU1mPvPqGUQ5ktGwmQ
WCFCbu7+Fo7r+20icpaRMzesv9aNoXJiPi75g2LOFeY0bZUxGDhwBqMUzUAMj45OLs6+o0eTgUgU
iKBZBFpoXNN7GW+vUCVBbCfVjknU9hq0qYAnbDCAxfClLI3QdCWxn4tw7eeRLy+dOo48H1kEWK7Z
Z/c3Iby2uzTiZp1qYo5Y5Jp5oKIfOPMMOyKwaG3vyqLxiX2q/UcDny24+44Z/h+dhHgdy7RA+m2Z
KtE6EzueG+IJJRp1frJC2EAmxhHSv75sHq2xzMyYh5Udlt6M4tFvwpspMxmMIr+nzo6wLjHTmPkx
iQmWO1Zu0hw5otLSP+4PVak4hXj0va3P2TQ60VpIa9L792br32Q2boXZFiTxT2VFioXUblW1ANf5
/3tpPfj5EKSY4y0221ausq2gtckeqpFOzTXKZOwKzAIDW9AUqrJjtVgxwdmlgp2vHo94TJbR9L+v
JTK95p8cZQhR5wBft62mrB76dSermsfhuP3iymlk2vulxdIOiePJt+XeAYG1HHcWMY1pxmAzk5KP
qUpULF7QHZXQGg4Mbhe7BoSZn7STgM4AUthsbqc2WMxaImqHxfqXLnZEWGbJURqQSXJxSA0F9oQ+
IoC9Xgay9eH2C7szwP8gtTx9ZZ5WhEyvNvxsfUEB79+9KGxeTMZ9aN/TDDQfrTLu+qh9NehDehU0
zKnti4/MjoNuKZNnyEXY7PoiQS0GLK5TJcIfDNuKNcvAunoaUkXO+Gc5f+OO1qdi7X/wGs91zLgo
11GnVJ9T3hgKXX3f2GQqbz1eyTsnFCma9aM/oickA//8Qzg54nRR1s752RgBQGhkxv5LSZSPtrwc
Zn3SLHxtcXa7e45wr1LyfETIYZOqrlF2+onQozayy1/k1QKaoPokjYxyWDIC9rVqsm1Nkaw2UbpB
Exp6oEUdjxvHZuyiIkhUb+t3pAg4uuvop4qz83aqzS+nWip37uVrUwUX3NQI/G6vuvqLRMUhWWDq
xwQNS2F264bquObYNiQi8R/no47/ktj5QGqLudotS1pcujoB/ewPkB77Vlptv6Oy5BSPgaRjDKsJ
cYHqNvXx684Os0SvszvSPfzpyHo2kslnsMLMdfxE8Zkuw2DmNdv0bDTXkW5M8Wx6DNk5VO9efLOV
v+GeYDGmw51bJqpJBVSrETBKdwhIQBl12ff9bjS+N0eXMkBq8ZuVFeewK6H0cZuG5zALQZ3tjmvc
Nb6SsEeGrt/eenv6wjv2/8btsSkau8G4Y1CpwASK+d+o4LypnFrDpSeTDm6AFj3DojsTM0LOvC0b
4uX1PFvm2B/D2KrpmYy2fad9uM8jKpWxqt1yZp6n4bpU5KylRHLnnN6AIsECjTWKCbrvcY5uibQt
gQCuxcfDn8fofPbLG37g5QVvwn4gIJf99O5sBlpJZIuc2jW+ZuvykOwAXxmzjTmhtxyyXrT7vWpd
9thTR5eoFN+l8p/GNV5KFJcJiu1/b+ZtTA0Vamziuz4SsvwnADFuozyayoupU26pjKCuDXxTJoQj
XFOU0gC+bnHgLD046KfaX8p/zRtvKBDGebm3f4O96Za4nzn0T7BmouRBVY19H0fKDX4rTJI7sXLp
sRcH/4PT64hNGSxtEp78WNUWLmcp7js/95uVOOjZfKA0J/vV4XV7AgTD73GSnO4eFHw0MI1O4boN
YolxB0OGsvReBZwHj2gfMO2hja4n6/7pm/1j6Vvd3nPvFsIsSkxrERK+OCpaJl8kuyJYtx3KqJMX
rqZWtik6arwn6eXgUvsm63nMT4iuE4R2wdsVD+v45VijCeYLglsrkkVKvayBXau0BUiNXPlErQoa
Cu4WvZ7l7mbAsk4ltmeI84BiiY3cVcE7cNuO4OtH5qMnejgY7i+E2pzMj4znUMzBlFMHDk1GC3gK
x6ereMk0ukVWoTB80B0sPvCnauEbk8tlRoZvRVUcphOnwLDLo1SCwikvpTRf6i8vS4gzul6mrvor
YprIBcXYiPSBrnDLMsl/sPJgvSsOMyoC5la/lSmStQZwf9f7v0GsgwKr3Q7HpRnU+s9uKb4Zw/zS
gFsTeeYDFUhvu8oQk/HQzkCV3HsRnHEMFiSGff4Xpv6FXFi0y45r1Y/+3Trk/CtGkGUubF+uYTvY
prYMJCqFncvXQEZmwJO+2u+Mdf3M8JlHJZbltL3NtI27zp4/BSSlYJY17p6naCabiat9Gm7nsYUV
2P2qwKzCuSDZ8xLYPq1qtU1rqJx1HY9QUu+jiyZ09vAM+Cvv8fEvg0Amt254NDqa1cl7Jhln/Jzv
KW68aLCmIktQR6HGQhChCgt2NGon0bKJi4uii9ZNCyGYgleO2BaIUBVCTLILOkXXF7ZDd+F/fcKS
pRGB1qfk+9hxx5GySgcY0aSjUjWDpaccEmHz9MSAv5aNn5aQ3aTixXXDPBFGcGr//ry3S5ekQC3r
j6nNPIaD4jTxxVhg+O/tcqmcZouSRGRcOHMUXm+ryIDSa42+/jt4YlEjRh33upE9Nx48cRejOuOH
Q4/dYQupgK4G598vT+5EsBpY7ALLQ9XD4hIGmvNUXYKmrYYjbR0JRNtS55mxcjqK9eTHOlS5dMrS
9+g6o0EuFIagL6IPvTU4DmFLbo1cdYJUoj8EzQyEIZcOQW8gTUgbbXFmNqNlgfkdOEjqR9BOG/NC
+yILOYOCSeP9lgZLPjvI2hNk6csn1Y8YdzeJpSdQpqiJ1q1Wvv9gK/BaZiWruxQhwwgMcIpGe62d
LOYwgbuPdDF+X7sgLEu6+gbmgxp8OJtZtAJqFLSLnGnaUou+Azcs6xgmxb2tiOu9L9sUnASfXJPc
Z05a1fp1XFizSXmKnuCjZVlb7yUqAnxOiJEicIXBJQpmrfJIG8bUW0Boh7TARpK4c6F6oWF7zPZ7
B2VubR6cRdYKnjFNvc2C03CAlgMvDa0iOqRQhhsvayzylRnOQBEvd6Pod+FcEyaSxIlSgEt9gDRy
Zd1ahyXcELaAOtcea3XF4SdSo95QvaUXtuRusEIQvqGx0psDx7cIOptBb5JfzNeZDxcp3sFK/3Aw
liD0ddcqp/d4L1jA1bqB2XI1VtYZuAZmdL36SdR6UD1JgYl2CLROok9cGD73yRCpIqcCagfvHp99
B+egtBKvhJYH5ffSfX5GlwIsxfGHNk1/awB0yRShoHutDMC4DDXugo1tFEiGyrO/yVoPPDPPnsvE
5ten/TZwYdzy2YeqNrO/SJ4Z7Xf/ltfEJ9yKixuuidfrSLOAC9UNezDyXUnOxy+G98b7V0qLLCUo
qRcHyJ8Adefkljnk/3axD6tGs0scD5VsVuOFD+LOYKvRJKuVG/YeKvoj0cAqWXmFky4zPGNrxXm4
4xVHWGK9rs00WxcVj/O7seC8G5Wo3uiEQADC4X/K3s9Ai0PMNLNM7GkO0jXNZLFz3ekFi1eLn9rT
a9uln0vaWd1ZxtbFzRN5HLoljffCazzPnsbf1HiVo5O2saaajU3hjNzGYsnkut6vu1bdQIbOAGiG
0ArWwdt3u33fm/vHr/dow7u3gotmnEZi4AGuGem+wlS09YfrYk5e0G63WdyGz2B+MsjhGhDRKk0z
naO1o7eCzuVO3FaC0rHBIEHx91ol9Mwgkh+uUqCYzFQURj9CppOj7gwMEQSUX9qLd9AUeUUHGMV8
9l+hAGSlzSg+HLXr367/Z7q3dAtnrlXOgaIdyTsziQmQDkhVpZnKm2gbX6EdYBGRYpOiXsIfzotm
bRBXsos0rMrnKh8XdWn53dtV40yaD3Cj67uICfk4P9EpUizu37aP5TsSaOmvGDJTi0NXxJiIcDW5
wB7NKuVX2K3l2z//OYNbb0+42pzsC2+jy7acgoUiJPC3luMZzqinFio+0LYDPRN8ALzl5aIG+IzF
AvgBNlF4rkgJoS8pbiWReg3WDFkEvi3EDdNCJks0ORr4NViCUof9piGSNXwO3HpzNzRCECGlVYAt
UMxBEF8ugeytuAtU+X5zFLRnn9QJjpve6LCytqmqANebXDw9aSgrmatyNYo2Q1ehpiSXuucOArBw
wsDGpQiwXejIlmmpRZrxhGaRyZo4IkU5fkGfbfCJ2jq/HyIq6N/lTiaq87p3/5NS3szjy1a3r5t2
4UGdD1e4cH8/FLVPmtr4JjUnH7QnC/aoZibKf0h8hI7lNYix+qXMzRTxVpqrNCKHYk+FjH9C96ot
juZMEVtDfabs8ovXqJbPYuudgDHhEkdPMotLpxccAP3UT1RPSE28vpP4mnfWTFDSQGSnjm/+pJZU
TtMYT6thiZ8o7Evhl+UfTepXFfLDSshYzeG0u/ONAD5YyXTNXaaRF9rSzVxEbKQAa5D+LzMcIpGO
neXFB90i9xgvbdqxPvXhjef1KHKPHy+hqHfcBBN04ZQrUCjXlRDb2ssJRGEfP4VnHyE5dU2ARvTQ
riZhRuOSphfScefHRTK5wulPCoavaOk4mHvSy5WDcns/CgKe1N1ni5UdCvEGQgK+NGvUc2tBMewu
7FqtROJ47KM0ZzcCo49AT+TVItsiBXnoQcf5iD9jL33kqQzxcl1554bXIddCCvR+fprLi0oE1cmc
NmJz4gOu7bhGQuVpXeWzJOx3NB/3TPuv3IIYc/yBtN6mOX83Nequ5LicdhZNSZIWatJUOxI9VtSE
CPGsr2Xt4tD7BZtS1UyBslIOvHEjFtMZJCKObjc/2wWhPI/F5Xcyx511KDanIJgjK6W9U3bJBGeZ
tJhcdEu+2TVoFE82q91eQpOn9cuSBIO+G3Z5y1SICQQq1KXCAXhcm7C57/85t7UgS73PLeysQo2A
TwxGaFvVTUh5eG43joOaN5lVJ6TSpYH3r0asAS+7jdPRSksHY/CIjIT+5EHk9LWho9q72gDDKfDE
Tyw9XPe71fdimeWTekxMN9D90ZQ7NmFHG3mfg0nvnUld0oVzbHWGG3WzWkAHa4pACbvin1ePRNDK
tEos/TNsscms7BcIfq7qQmdShePqddseUaPEidiqjXvSY6qgruiTOz4B3I6nQsC/RqkgQQpU5VpR
mHdsX7W4fFyatvzCSQ2Bhs50TgPHJimKRaxTbUZF/ibD7t3H7UbXHx5UMhK+RVlzhHuRo+6KsGbC
T0msyKHkgvbjSPN7R+tbiAGbJ1eO1CU65cAQWGdTZUKWSfpmDwWln1iG5VT8YUVaDpODL1QVHsgH
IVn6awgPZikDkeJ+N4e091B1IqEuoHxt4l/0XdTv4BV61y8Xtu9ZrOmOKp0hhGLlXcMXQeA9KLaM
YMywQfPOR/FT260coh+UcIYB9MjS1V274AgCINmCooGtPjrJQElSFRbbFlVMAiORhgOcZBYvy9UQ
jbEQZzQqw9UkCWJr/3qGg5nN/81dKnjpE7Entarvxw5MQa3/5Qxf8tHOeZfwFii/x1csx/KqmGJ3
8I5aVz7MWoUAvowzKCdbyrcTCtvsIY0SOfCrd1BLG8FoBhiAIo3spnzyN08JuWkH8KP5x66t4NnH
20qDXHD+6THaacnpoQ5WlxPGBGEYnMQ0bwk0FFKHKC/m6ZdfAl2OcmMhskbWJMIcxeIBb/FHWNfD
z5NWqO6E169Z4i9xtBLfrpmUhRm0e0vAKAxFMW2gjEx8mrp2RaLNFB+nNynqiyX/IIr229Jt8EYz
5rLFgWAsbW2SXM1SNxaqRqngKeNRL4akyfpfkYzSWLJAYRzfio18Y2wPcKmKdwM/OjfnzQDdRkWc
AWaxPdrg05KXw1BitE2yxebXoAtp6m54NFLMwHBt/Keyc+ALmmsYl5rhcaTVQltehbtsN2dnfO88
KGM1ZTfWjhKoq8HfPNE29ms9UiTds3zdhVyrhBS9MMK5/DHCH+D9uVx1ysTq1GarKX5BswG+pAx8
X/e3JZYsJumarYUrV13mJhxloMbPIL7W1NkaT0uWbvOBx451chdQXjH8OSzyVEVNo1SIfasMIwFP
uFSjHpJkj9mR4WG7bCC8SeQdQLMjB0TcTih+sNkEyGp/x+5QxAJdWAPrLx8NVF5IAqwiPjaoeE6s
g1/1zary4QH7PpFMG+p5jZtvU3tVIJVxK3tbvKQL56vtSnpROOIGMyQcizYNx4KKcM1IpKB1P3Q6
0KcMSDoTUZU9aKp79V7L1Ro0Y0ilVr1PGForwz5NYltjM6qmfJoHyF+S59zBIhLzVO59o/yAgO8I
UoVNhFBRsyswI9RfKTtYVqJmy4Hs0lhOS1uybZYyYopa7X2Ism0KWbINU7JgfbXp+hrRkUwacrZZ
yvFhBBwPSxA/8RrVjsHMiCUUb7tr8LRmQtWhyqLycNdLej+xWmh6YihZqkHLv7HA/IbHYbEraiVx
Z8G/JpdZ0+zJIa+PiVf0yBdG5aopkVulSxoMytkkHks34sdGN/Mib3cq0/yPKkrJyvnEb7qURj+J
439rVD9x9Gx+8VQwBuZwz4lVMW33wdN0nJ4jTWb4UfVH8/cazTZP+Y6nnVvbokZoRf//JMoCxf2B
btvopc264Aq5n7F+DXUSOPiPbTiVsiKo8pzCsp4ILCz/sq2HN9tAvKdFaruB4zTDsdfZs0Ipy5/L
k9Gbj5hqr3MY9gcJhU/1VjheVHRg9IjLoeZgi2Hcp52+y5Iitvyv/8ITt7+cLtbjaS4nsbjG2928
DmssLOGRILl8qAdvBbFQTjVybm9AhfRmzhkFYH7Ju/uQkDoJJul2bZ1J2Bs+RF7RHerg2DAKKPs4
42yarqBQ/gCpm8/ohvDtiCqiPFJiPgv01Fcy44TErHo7b8/EUwb/Q/V+xaKurW05aui7UEmfV0i4
fOP2iLbVjLZMCLLzygMOBr12fLII+R3PaXnNKn2cpQwPp92DfFlj6Sb7fA/Rk/quaw36X+gW8rrk
uZNhmIOMEnbdLNPvwKBun4r/aWHsko5jZzKg+5cCiKAVYCR99pKcnrPNNOongr0lQFzFPtQSb3J+
9Hif3BrRtp69DRlmyEZgqDig0Lr4HVgzz5/FreckFzoNXhM7ViBS52JzOyCccW3Z4ByHAUgQjh37
3pn99O+KqXxZan2rVJpKAxbM/a7kGttK9/79Ej3LNX6cimevlfeedjyRPW8aKLpDZUUPqJhZKQ74
mwH4Hkq5cD0z5KYhJFK56GuuM4GzeLTNKPuqisZVPbDmBQHjIqMpwMiNqLOsXqATv0Y1/e85EK0c
sH5ijMGABkPixgPFC+CigNPobZqCYPUj5CeYge/MZ8vHwHzW3ZUUBwSOaqfwR2Jd0b9fE4MfMBID
hiSzLrP3Ek75KBRxxs80j8EyqtQmPQmXhImFzyZDlr/uz9qpPcVlazjUFVVNimnhmMRpmo5TDIFb
S4EJwF4TLdE9LIl4cq4otowSdMIZIMUj+ReuhWFyGzJ+iKe/3ZlcRlesq05L7PTHm1Iqp0E4EaXe
Pqjhjs1e5rF0nz/yOzv+PnL7ZVyhmSRynvqemv9E4rFze8gI0ZTmyBO4UQ2oHia0uS97oAIj4Dou
Ae22aOxzNmKt9XVmVm+ED2P2syhJAufRrB6ci+0/KyCmjTaVaz/9M9Z3Vp47S6DpAW+Bz6z1APU5
qtAiDYYXznMX+bVvE1dD2OMsjdH8DXtOca1UMhvjBS3XdgNTTlLFy07VjqFoPf1kbXojWJWPS2rh
X23OH1OjOOILtC0r5tqC1DKt50fdkloABMVcMqVDkxIXeuNey0+A1DjCKn6WB7rz+8eS5e4JoLCD
xCxGAj1oovKNlGk+zpnSPxvm+jofDF1p8087Q6mjp+fDg4wwYvwgRhm2TXf6PUrJg5jHSYhctrJ5
6s5TU64qASHhrJ7+GEkHabwshI7LI3kYFgtge09E2OXl3nuoZjvmPSpIW/aq+W0XbLe4a2zVrchz
6FOhvMD2/VOi8f+OHVs9M7EKE8ajVQHrHxgSDbG2/Kp8xAjFm1/rg14WqPdNEYctc7dL9y4Lcvpk
I5IwaoD9if9Xj3/JDOye+3DkVUZ3N7q471geNkcnbapXS4MOFx+Q7jRZ0F7mvzpYaAPQAdavFOsK
BJEpRXi08GEihypUYZf2NR7HtOeEk6ooCIpm+hjO2Mvbwcg/FV8VTEN6aj7aqggSSTEVUvXNFe/D
CKKFbChcF+qYrX7p3YSBy6aNQw8K7xP7pv2bjxiCazMqYk4QX4Ur4Vfhj/kzdSE2GGXuq79ur/iN
SwM35+SyLstSYS5weTgv9dKN4PG1ezDWSn56YW/gzWv3c4QGrX0GUc6GIFRqLArz6vpc4PjeFvUH
T+8SuSyHaBM+OUww2LleyaBp4ph7uBA6R7sy36z6XwNE8M7MMsUf9BVxn2oJYEEuEHcJKDxXju2n
Tb9TW320+ziRSdCTqptbqT3uFp0xgpLQIuly2Kz08P1U8l2XtsIuco1tAHu3Q8AMxnuv6C8r+Mq4
VUe0O5/91zUabJFZtcwuUVgBvkNGW5l93RqOu7ZnPiY6cpu3BYtPBtV6lXxqIxCDDqDVYBDtcUjz
ODUKPHlUxcQ+SPRr9e5ZeIL5sEPa1g2eW3k0ZC2zc0Osy4lKovQe1uP5Jsr4KieOb81V0p7ZW2k1
YwDRkdmjr3BsEgn9NXKkT1U9gV2B+18+BOXNZeDenjsPnQC7AOUXE8M5odtYUybl6+bFOgJ6F26d
PBTDygs9D+iLmAjfpiYYef2Kpx3Vqo8gUzQAPSE1PKCb1K+TJhed43M9yfatXnf3IvWb651LYQl+
LBFJnbdSXo4awFQ/3tH8+qlgUzJ/DNi/RuJmZqjqd2+5NSm8rnI1qU49EF2CX5TfTxl2T2AWSjic
yvFS333PHP74ptxXmCqoKoKPMRtABIeasFyZDPOPv0Fhhad/Mf+As3jymjbJcW8Wn3s7Xygs1H9F
0k1LS+RpoLrmgBdEohvTuXlUD6BPdzePYnFrfW3pCPqSvQnFtXj2InWni5oUCW3IflrF1XPLnpcK
OifeSNYITy31dXC3Uj915A+lCaTpz36OJImKjLlXkoMwe5EsOJxv+0bthshSkm73ouCkX6hBj2oE
PZw2wutzhoQAmWVnvxaQMNzZSoiHZEuwxflPrElxfv+5bMPI1sCM0zQwqI6vcx+K8iyl8FV0c4Xx
Sm0I+NlwCa+vXkU1FjzT9dpnn4yNCqfLZIG2K6Kxs9UBiAHWYYI/MfdAb+raCjulmMhFnx8rjh9a
smNsc/srzWWyuSizQpTK8RrpvCnnwoL6q1kuq5jTGYPq3qFNVTaEwb4TYTJzjEDZCY9qUP91O2Mv
UtLhlUFNF//bYtUHNlMRFyuCO72uBeQDN+vGGB+WkSDBfiYD7O3Ws5rOPu3ceNrmmsdhRMojpFso
Hnsp5ROvVPXdiL8IrUXF0iw3X+5HhkgJ0GMTSMTmx1qbzm6V4kc4uA+ByzwbRm+2FPBRKpaLWcc/
w1KwVtKcG1/3ELVYTnnULXohBER/gSm6gQqLE8A/Tsg7TWwdSunQYo08EJ9KAgdiZKkT95WvpoOq
LGKuD3eJJ0hZmIdVEVFpOuq3+CPv1V3HEfc7wRcPrAswe/QNp2f4qRy10AESkEjXbjnar4r6bBJx
bSoXQidTIbIakjXIdqLuhT7do78zrmly8jMCuD0XbP5+gcGM1kgW38g+M1BgrmD3LeXDHOIqQdbz
dJVa1524s1isb3hE8Jbp+ZCsL2ic2AdZJ8Zsxtfs7D7HaV75gGfoxG8Goy2AMwiy928/GF0Olpt7
OBaHv39xrTYjkbjo1zm0linAEL2IkJIxv4hSaGRPZwcIbSI6gr93fxCvKKWcKh0DHn5gwCWOZhbD
V4Cnh1WNQD8/f6mF8/e3USehTu8zI6UDd0AnoS2ya7+BTUWGP8x++whUdIjKzHXfMYK7wHp8cthj
o6xsjb6lS5VbApK2KjyDK8U5Bq41gRKSd1O7qhGyBiIeC0oLM+HdnXCrx7g1vIIoK6S2ZWF2ewp+
kVvco7afgUd7Nd+m6cxKYZ7z8sMPFM9XranUtRaAbsHd2IRcDdhTjx4ZGSrTXmiKXvd8ldn+YY7/
HQ+OL3OIsDXWsQlATSToP8tEPHf3d6wlPthgqUyQma0biaCvOEPIdXB8ZRSpIvOt/nmCWQfTo+/0
GPXiT0PU+TcBPXOEnJH67Vf+dGkkyGvv2rUe7TWOV4Zpjva+BGspjY1Jketz1fyKIQUKeYRBQTfo
4gLJu6gAmiwIqb0bRrNaFx9utHS3H+w8RCMnhO3FbdNzSWcwUADscdffyIbkK+nbYZYjkbbnrZgL
0OgS0/huwLCloQYwyGg7lQs8ZeQLujwFxJlhS4IAWQx8/bRmD7Pe9OEIUoCqY8zJ8F6UOs8kbgYU
Lp+Ehe1qUdSQBJ5daPq/2oQxx0vSyiaAizhX/2NIOQxi6JyiJkjlWoQLwnMWnCW/A2Sb3NppL3G1
Mxo9APEnA4+rRUbg4pJ8/5DZAvEF0TGQoTUGR4gfD5t+/8xdu/Fg7he8kgD0VK2D2lPjpTJMjKq4
IT+rLVyvRpYz4d+C5MUdPxUsyzD5J1QgLt/tn7gSvVnYb1IR4Mrbg+wD/5HLpd3XFtEFKaQq3yju
a2+Heh2X6V3oEe7UXZrfS/itXH+3TVm2p9zoywOSZvLc5PrOQQuFKnKT6LxK/Efz/SvakGkcpoS4
UjnGU1x41rPM2CFGSmiooBV4YBI45FjHAopMnN6m1GEi4uBISkr4KXtlBv7fmsHRtgw2yFu0gQPE
Oyt3eZEAUChZeG3+PGv1eCPFIyA5UfClPPRN7iR2fJfqMCc5p1Hu/sT0nndANohtSpYTXQZmgSZw
ezfhv+oJu8GqiH9/iEmawaJO/JGwelSCyQBqFB+Oerhjcw72CLro5+mLSY3vg6k/8H2aljlcU3Qz
DeSVEP3DFaDunRLWQt/FzhDvrxuqS6Mms2x6a1UjYxknxZSLyUSKx3xDinfjfo0rH+B9V/Yiy+5k
yRaSGHw90e8C50t+EfXX2ldUIdgiVFpZS4FaVU9y9PYA0TchMs7c/QJDvOkuQ0DzxbGFgZZ/jpSK
/ZyPnu6IsWpxPjZR9cEz/aQQW5nkPUvjztENBtAoiezGpemklX/hWcc1Js0NPCXjM1bH4pZ+48Ye
7LkcfrVxF9kyQbi+6QO1Pq3VdjNKgorl4LkCm5m8IYHm5dN7VsmH8WOovDODr/AXdb4gNWkss2jC
2hDmvFnXM94A+79gxSwwHzYznFyXzV8GgpBW3Arqf+aC/G8kSUMuZtC3lmpvk05F60qu4TRuoj4j
WAdCswkPmGtNsgWmB82TI7nEgToRPEVr7p4+igBgB+Ia6kXfC5r/QzEMzwK43JTRDTHJGePIqzAb
ckET3LtTnZqhtbkYgyLhBQreQe7Mb75HVdQaysjDRKkJgAJcyMreODIFgobXO1NPcexKKSbboKVc
+g29bjd8dFAskEaGyZLTqBmWQlDMIGCXmM6P3XJx+NV2O1ZNVi/09p7TgtTSDRYbgk6Ahw2Q67zB
SkgzEog2iXX2O26I21w51yd8sghVbn82yHb6DKLcOIf95N+Fs77+TcdMb4MQdGIXP2eSbbO7J9Nr
oNT3cmsoz0YNh2yKRZXHddUNgUmb+n9hFLMHloZ01rQ/Qs5EPozlYjU3C4D/al1FRith1hQi6Pip
DrKsjnZ7CpgqqqcJAcCSzvgby2AtWYQENCd+pMCPNSlaJd0e9uh0YN5/uAyiqtkVMzRL70YeMOzr
gD3z3O0t1jTFRHBi/YltlT6C+UFZ5rYurwbgAXGTYpQItJwyt4JL+SzdYnewnkUfgkXzhcd/wMgx
h5Dm9y2jQ8Vja8cw3Pz/FFIjOktECaVt7SCrIrqVi7tUfdKHV096SGbD8FNEmenjM4S1I+/5y3Fz
jmch/CIyAsmAxjw4+dLaTTeAtpnp9ZTShrVM3wMVtG4t0UDne3YlWr1qY1ZpNYGadhuz9TYsHd9x
J/KmIKRI7/RSCsW3qX6XfZA/DS+rG4abDrEZ743WfHTgWzutZg3KqS2SkiNvJF0yoJdkzPkYBuvg
a9bCMNK8QettTTa9W5G0PBRhlphk42Ezy61Qtq2fZKtEv8TLdgXskxZ3wdYsIv3b2Md20C30XUZI
7cGcLqXKGqQEh3VJIIflMO0OIsv659m5ZN1JCzi2Mt4jM9Qgq+ioE7Ad5EOuDuL+v7tMzg5ZVQV1
WCN2z+Vh+6j6nd8exRplv7cVINlEqIWBjcqN7lgal/qYnjIbh0i6fX2c+oXT+qrEWDiqQ+SE1KKv
eMr3tNL8JFv6M7LFb5u6OLHpzVRrwnLxtbu6faN6ttksIwJL50nPk7fYU9nH5+naim+MSL4XWqDY
tnA6v4GUvI+3G3D45RaUziGG0Pl6UFqx6amYp5wZKTSeoN4/Hq1tLu6ou1RpkfSmvXAdWIQWX98+
vbDp/gyOemzdYAgfZcQ37dzp51vV+vCVmY7mREmWLY96crt4hEU/z5G4/+uEqteEAyEtmCyRCgr/
0OuhI4NX6rhPhX/0t3kOgZsra2wZwfO1enB65leeRTdmB4KXWZMvtMDF39pIM09rTA5kDjnls+PY
6+SlR2WmTc1rijDBoa7vGaZwgd2GXxoWPx0O3pGyQdAq0S1qGSEyshBJ7ZWYIeP2XORKX5ldt2cq
WxJ9gfVbkj+WTZEwxhhQu68UUnUVORAv8ib5mM/j27UKqKncIPayBPGo9bVEaOyfFDYJ91LaI10r
f/D1Nt0lz0CzQKmFc2+0e3RUyhpGVFFoG2Y5qAz0IVZEh0hRAd8DHp9O3a+yI2epjHJX8kSPOEa/
0RHV319zNIhlc3H02IXpA5PwdZ8kp0jdndIzXpBLkQUbHEKa5iMV+fcrBpeczK0hKk0p5Joi/dMl
yT1cGgjVn4tfl6l8XvKMmiYX5B4cQ1JZrtv1RlGUiR+lUA/LVcEIJPZHRv9lm/m0rg7aEVOMhPMQ
SiFphiqbMU56zQoH4wVz5WoiWEgfHjH2xBC2VIPlNaimMHDgteeWzADV7Egbqdak0sPDZrWo6MT1
adS9bYZVvIIYkpaEleoZEOIS/yTTmEyWj0sSRupQ0JOHS/jyt/fRE4olBO3CTQPmIoYr92OXCb/t
2YkgDmU0JWukqzFK/y7ejRaYfNON4TjgEqltAMnrcR6LyOxn+gxosDsG3QeOCatX3QmVGZ0HdaXH
VSWqVrA9ZMLXhNT3jjXCPY3uDzwD/adr59MdXlZu3THUpVo2D2C4mqco4Maj/cibzkRpKBHukpoQ
6ELVaUi3TLq6iqkPvN4Ocan+FtN4BC4SRn1rATawvAWk+SL4BzdNFhwpUKxsyL6frJ8qayLbx3mv
POq6ltge+MNWYsHS4KpLU7pmrKcba2ajqNJA4s0FxuG6aJr3Npb+W/T/Q//+G1bWSFHb6EepXxer
+uTdvFZ3pMOEyhJAdPXPnjkqHyWzS8tQ7ou5S9Ra+HKX71XBXs/URCRW0eHjXSKJs1qnRXYCYclM
/muRPThzxRD1ZhIhFID9Tm4mCSQoQZG5w/rXLZzxYQVrNu2nhrJK/0Qo2g+cQcc7QgmR8ZnjELFH
GSrA4/nd2v9iENiTysl3qdzPG7l9mTNIXyRRFnUSGBju8UBJmHyDxz5RqYznYfcm4cTlvdTLwZu1
GbXkSbOfCnPJgZDc4dmnSWEnS3EKlVXL9MXfVQiVISXre6sV7p4hFyZvC581C7cLBNnwT+P2sJTV
qBaK7VPIBQOp5j8+xjwS6ugm0kK04lVzt7peeXG3keRnXU/kNSEyhLwb2OApWagG+LgfywF4IWUW
5+WP+MNi3lNZSBs0OK6Jwx0DS00TQmjXy8ZdYbX+gIofeAAUkaWmKOILApA38vyrnnqHclJJ1Ign
Dqus2ci6jpr77RXlCxClyi81EPBF5DV+IrKSQyS4YS3t7ZPka2h1/g0OlhFzc5ymGaJpavLdDbX+
GQgcW4dSE1EYWRdvgtyl9z2CZvHgry8z1sQQ/VJDOZZzVvkwvhlz8ifkKFnz6weMoYey9hW6X8ci
lv9JFpklX4q+DgM4Va3fVqSsFlw2nOCyAa8epqW3pM7z1pSY5MvOKt16yKwyrcxdcQsP4TMuSE7O
l9noxdYSL7wmqYmh1Em+fYD+IgfUXVRunxvQpmLHgkHjDBOy6bt+N6GgET32xYi+teKBJLQdvAnP
rzvjOnQBUArtrAREps9lMkLFzufLPjecyxsPsFczDh1acxZYPZx5IulsF32I95Up7c5+M7wLcZnF
FR2tzBoi1i9lsWImDWAJMxN86O8lenJbv0xc1dsNbI+rdcm399g63va8b2CVdVZZSB3NLDAmbbQB
Q5boSXe2MUcEzMo/YayAljUnTCNaT3LZd5TvuMvSmg+MOqMQGtYKDQijtR0nnw2ThZQ5AoQl3yN5
apBhM6xKiVT/c/9sp4LqucLV5g+/UMgZP/fLGgHXIPJD34z8oAGrGPFjfmpyfbfvoopHk0RmSfX4
eBZG9FJ+LP4vfSMELiKQNYc6YJ+CmhqUP5QQxMTSBUCHFm3dqcXfhdkvuwiTRBqzbJSKOBVnz1KX
2YT/gA20WZj6FlQs/C0hih5DV550bPl9Er9DZvSBhTK9sZ5fyM45cHW1eX4IMomRTahzZ1Y6R89/
07PUVnzH4a2ti7G6W0gkC8F/7rX9A5T5pmZo8Hs3umNcAoZop+5Zu2dulowrEwYecHfgH3N6u5KW
X7ht++Hi6DbTsuu5ciOOnkB/6f+Q0M9LL/1mXpOFUxtDVVUDckXuMCcKXVqiwcm2Vd4LpmnrhHrE
UD/Bzop+XouqVk5MZYW81mK5CspYkuFBiZz0DDuj5BnsLtLhae3HQRGXnqVvYH3bhNKp3f8RR9K/
COA9siNWk+0iLGkRN9pE5mJl0Nepriwt7TJSlJZAOXg2JzuSTDaGg94WvCEr2EMslEaRq0VttPm2
svJ7WfJJrKLhDbAQ822JnVtCzNXna2sJGj1uxssCIrumXV8INr4Ck6W3VXttl3w+3Imy4GFmVzM8
k3SUaf15zYLyKHDSDONJoYnQP1sqImoaNOtW+tSq4DGiFC/k7qB2TQ9g3rck1Sn1k8K8RTtK6hOx
qjO8ZalM8cOV9H7xd8AuKuP3qlVOlQgkgt7cgJBjAtrruWUtbM6XxM4smLL/ZiB9OyGzL31WxpbF
uVmAzx1weXMARVcPyYVe+WAZ+KR60cUS4Dc/orEAgnXLXgC0UC1vardhgrSy9c1hZBa2bEyi6e9+
4dozTxH1BJGNyGRbsZqNiK1dALWbkxm49hbgJlSnpQgge475v7n3gvvODyPsC1itfxLfiWH0CGOE
ZrcLHU0/r7MPkBtlNNPkqkZ4dm1rN0/GXlr2MpwhXzS+RUHHeM/0RNunon2txuyradFJdThba5x/
VHPVZWGHErwLgaMH4CyH4y/gi28WUo7dt744owP+Rtypk7DAsWtXXcJ6yXu66XbnzBF/ryWVBOgf
FoDPPtooecIQQTI6MtEoejGQTskJOEsfqe8YHy0imL0nYO9SwlGAKAVDvswot/M+uFqmsODm0IoJ
+Z1tfzsPmtQExLC/ggEljE4+zrEB95JoSsn+dLcQOSwvzq5qYM4YucvXrhKOVp1fF5t6bw3tBUjy
NSwW63gR2tcRPC4KndwRWmWEzx9VGKtDpb0kQCStrq3NQgbnru6sgd/oXMoL2i6TrBpNz46/aRF3
dWpm+w8QGgovJ9wrU40btETOxEcw8y39uGEOuB//j2INNXpKnDGOc7zF9TmNUvhobYn+4sL3L7Rz
ESC6Cth1SoERvrmBMXyQZV+lpZdUhejuXKjBRkxMLCtAOftAMIcMymCpB7fezUmRCj0M9vG3uzq+
Uzzs03Nqw6oIMVBrYw/wLldaKQGqm+9AqUr6zM6GAReQ/slVuGgFOy/qyu16SiQG95LU2xcJs/pz
Pqq+wsx2+QCoQ1L/9iGtkprEOyj5tE1VGg3DrW7a8tfEyRezmjSH0o/ncOXCzUog17+o4cv6L1BF
eLf1cHXeyt4rqa+LeofGu8l0GNK+Ws7H9JDDHuagDKV0Zw4MjjCDB7R+FLu+zDhux8X0b3w6yfux
q+gKqIvTedP9mCp5Z0Zlm7SGgf6ZiydCpy9ihRrezpbbU6qcwvulQAa7RcEAkrItpv69kHYF1dVu
HCnWmAMnaVY9e+1qZl/1HCDj1i8f+Ov1Grmn13d3NbVSGQ10UZEupIMvWZkuIK3xch31Dwfr3Vv9
wXAij7j8G4gIEbI0/39iuQPg7OYHp1ndng4ieCe9MlOZCMeBdGDrphrMQls0usmXeXuxHldrJ79c
7IywGRcUNmz/QCcHjynWI67+Ilxpo+KUCSalQEfQARUr08IrUnXYlZyk7tl143WSnAoocsyXRCZP
l+fL4FG0K9rgaPymcwcDKOAPnrYAUZSRg6/ndMxenjBjjzAVWl5O8cybRWqkAtCxV2THuJ+qiUGt
W1nS+g05cve1Fc5tFIoEWV3W+OxrmfItB2lStkdusSamyc9zdN0V5gD4mqNc33zymWRbk2drA/V+
hLi8ollTouwxnatSnGlbETroiYM8xFHaUCX2qbBWPKH9WXlXbphNTnOL2p6drq5mxPu6UqA3J5ux
ACiHDxYRhPe7od+STqscxk/u/bdpyWFi3E09F51rvVjXqgQSuqTNxIAtjZq35qQVemPlq68qo6I7
if+5ELBsM4mTsxkFEUiSKqWljoW8H7NW2SyO8mUkdF2zKyQxvdQ22IyY/FaB8bZh4SaCNkOmWoMv
OhUZknsuZJd9/lfNV0p+Z5XatYyqJyxQNXrzB9Ayqt1TXXlO0e8V6oVCNibEyHJbJGggtaHMR0Wf
3aKDC68IMbgWbOiZNkX7ktJmUrvGm78Az7CpXhmvJS3dWF8AiG2EaA8i1fJYfTH7JYqq88/95fPW
70jeDdgWSGQDLp+TIINw7xwMhUcprJmvjXNlWk2ULAGLPjOPj/kn+XHLDy75BUzn3SOW9dlf07st
JLOLGAhbwOwgUyQKs9g19D2SV0qNpC41oeovQB9x44yF9Tkdng9HkJemapJpVOxZv1CPKGkff8hp
VAo79sHhmlGD0XGvxau7jLGgw1q/Gqb3XDKI7WjHxsnBhmq8OYbjNM8giwMdpQaFUqNiz2fJI5jN
mAeuS3XffNaS2RO+INKP/pvBibToGPindQiRC5YlaTA2uvQ7JaH51YgNK0avYuy7GGXkR1d5TMfQ
NnfHpJUfiy8BQChCzuQMk/chGYebPZeikVX4MdOEz3zWbPfU3ZgPcN4nv7jK/NdaSOVOvwdtT2PW
zddDw8wFj+FLkZoGHGmacQiHknKO5fXiJQt8FY99HnWQLYc91YD2cBcVEmEZuD0Mb/Qd1uGT22ZL
Z3LJOSRIATxR7F9S+GguphX0ElUmf+fxXa6GjB/fbFQ1SxAG3OCHeyYoj6wZPomdGGIj1Y/AFOmH
HQYq26Lj6syoCiueFNEw1j+x8RDWCXnOD3tebqpYMjrK3f5pWiNBRJSlJciUmOsLNk6enEYu9pMi
KvlfjWm1BjDoKg0PYb28yeVdW1hcFoggZvOXD2OZo+creZZVSGtnKZ2vjCXfS20GwwoMePz+8rgR
UqBdLDSiqCaAW2plkaXFJjSIOmm6MLRqYP4HtHd60Bv9QMCTHurbST35IhBOj9aj/Gmc4sy0vNxn
W8+Ect88jD68rqhrD7qWLmVTkATiou43wfog9V4PxEGXU4qY9LtgASaULBAUtRVu6BFXidnFUGnK
iNqDXE8MgP0lR92GjTigFeKoHAIOm4pIMwTsCWXMok0zHXfov+eDMO2sb1Ehk5fFTwggDSXXvIMF
gaq6Z9qw1m2WOJWVQY0fMB04UNhODEwNvshxbFbv9qpibpw0mnEYEK9Hl0DMurt2B9ZiHC+1jVUv
HZohNwnpwtvkHCTJyzy+NYlWt3+fHiBDsNygixSKJVhRY//8w3nFoHZaGikHKj6ucLc0M9daYTyg
5CtQiFhozNpvwNPWF0vUnO8eDRZ3lW2d26NRtcjlMZAM9k/Rl9P/9pqlJkqXoxQddQDl2km+8G+c
v5LAeIwXbDrsUOMH0J8uCe8Tgon7PZEjzFYwlKhHDz14/+0MJttYu8a/8X9rH7i7YGHWmPzzZMWT
vs7Udv4oPlw3vf9QspBA9/lr5lx9uHJjoeoqdGnYqV78RW02HkYjtkdsFes75xq8vsVKJBEot1U1
jHEZolp+Zh3gAQy+ENXbA3Y7gA7gXITkGiVisvTFmCXMjqMvo6BciSuFceGTCU5v4NOtM8aUfto8
BDRVsinydgVrFhK8kakzYCUonvduHbXaWvauCh1I7PvEiYqhU/wB+Txe87cdI0fr7P+Kpw2S4nbw
78bfXHu72O3Bq3ylMas2PluiRPjeJysDCgRmtHHYMYf2vCOT3G4lyIAmQqerZmPmletruLpmnGt+
I0lN4WDXpUNhsa+iiOOnSpzBzUKzxvu80yKI3mdp9QCzi0lmo6GtGfURaeaaCzxUJytclp6i4Dnn
k88r1Hevt3+LK0scB2BMOrFhB8TekUDavKqwcGFjZNocd22SzDN6ETAaDOOtnjxLd/vL5tis7sAP
4yQ6tL7p4CtkK/9UvWMdhd4SM35xPTfJpL1eo9r1n501/fM5ipscnQKpGVDoz4oU7JV/dq8VtW36
jfp96COvT+slH6+O+5KRPp+D49wy8k5fazk6aZvZNrIDmqPJQ+aF93VqnFvACxrAjjSAcUP0HBR3
2/Jos9uwkKIvZOnw/2xOdhbk0+A8VscuBhawS7oG9QRfKXIiRPywbaiv0uKVcefWVs3V22Wf7fil
Su8OOapPHdEFNE90uH5MfHOf4rgYt0PHXJVvVqRBHFa2Qn0gJMK4oLUuPSjjQJmF66VH5bT8m0Wq
Nwb+aXt9wvOofGQQsNpm0CIV7MB3/nmAtfGKbmjtAQBYyLoo8Dcs3xztPfM750jcxt2CwrrkrJ96
f9IGonAw1Irxr679fpibnlf2rhtnoTzs0Jm6VJTIgAjTrr4lzjulqOARlqd9CTO0qsq9OIy1z0kC
nWvosuG42LItUpiHzIW8VQ2M4BZp22d0S4va721r+8hxG2OgszQVm4NpdwKCiA8iqbl7HfkZV5FF
SbIUgO80gNnyNDNKVW73+VtOBKzTsk49y2223o53599qEcnxo/EmuG1b203D+lwSebcxw52J/Vn5
xkFLcSuinnlmS/2c4RF6H8Tuc8VbuliDzDYeJJD6ysrEV1TfvkSV9neZsDl9b+gBVEn4EW8gv8Li
uJoKVerKyfYx7vRH9/8Rct4eHN2zQHceBMunA7FjcbgAu2SNS83VxLTe/t9yrVNN6+K4BscQ9pnE
qiCJOFG4Go8SZLIeTdtHG+QFB8Z4tbzjL3nFVVrNudTCyUAHgpiGOP0VGRAejRG9y3UKllROwhTj
gPt4v6UyPvLCMCyZFv7tP1gjVhxikDRq//uAkPTuKB3TJMgG7j5z40716opvSeVh5w+yQcD1fRgT
LKBxP3RJngRirat5PlGbtt7RFsRJRl3Qt35DAmpJjnx9K8v5Y70e7cSIHgaTlssUMe4YYKlhffcS
olBhUVTONUf0VcYxeo3OJWk0BBUJu1IkUCMjNUBWHbvOsnsv1sq6uaDWeMX5srThVz6ca2g43LEh
AU5G3R/U1DMo+BuOok3efwLHYjuKbvHoNSK6htGm+gymy2FMxYjV3UC9ci3t2B2OwAIzdQ8+pNtI
NWv9+nLQ6CsdgFocMSda+4EWLlvZdykg9jc1aD2op551t0IbGvwTN4xYHvdkxUJ3TdqFATfO01HA
GucBlUUGljS4mF4us/DAJAzJZXTeOBVc+N8ZQZyBtNgM7GKS46xF2Q1hGcXeRhQWwLuoXsN0Ubx6
NdJsxpIdjXNXrcolvxS0vGqI8fkvJEc4tIeLp1E2Xfj0G6gqGogTRimfqbMEksvy2t3EQEW6t5+Q
msEvUoLlQIHu9seI9ykdKmH4XAARbVEPdIUpUXsf6owMqj2MF3+F3yuXMhJ/scmmLBKGU/ijTAnP
eREFwnKd/XquZGM4/ylf21bpQ5Ywgm6TNb0CqVMyJbcFKUMQnV9hM5bFD0nn4WPPfxiu+qnJAH3b
7+9n4vGrh9En0CEb88Syq65qgc8Nu0bY0RNruMedW4sgNPAC2Og2VdtsfKKU3k6JiuerhwvPkzlR
AZTM2bvUNcXKHGnhKO820mVywo7jfTT6jWMBhtu0kSee3k/kdkCMQx5rvdzAVXRm1kH9EZk7RvrE
G46Q4h7JLxX0rg5wBZxzruvT837R0Cv7b5fgla/b+qbxt1FSbYtyLc1QIZlf/pyXWTU+umregeOX
VW+NiyPCjTsufYi7w3dUvZs/IspuKsKeKBGnwZ3aNBMGDygHx877AA3wKThrUOgEH2UgiLh58sam
G5wtW5ypr5SaWVQCpv0yWOXlf2NmdgJchkXsBe4wpT31Ew4n5XGTIqcVRkDy5NTPfr6r0kHf37dP
r8ufnDzVW+nnHgghwQ2Ev11KmYSP0gkMd58NA/5jwdhCfTtqaxE9T1lj8tQj7mgJ8DuSXh9YCJJ5
W/4qJVpYU76YiGQKamfcWoxO/S9GewwXH8+z/T+ef0BLx7TTO3qfVRTho0lAItrXR0khji5pLgkt
HpHrvmfE6mKI6sFtpz32KEunEoboO7qVcfKx9W8QZANjwsrDP1BgSfgVU3lKLczOnLyTKsnTDPwS
3bpGHMiZ7FHbUhVeo+Li8KfpnertVdSXTjrPH1NREyAMjM5EjGh253Rdw926G08lybtLB2XHPvmp
efMns8VC7HAWO22Z6l3mWA44oCki2CiJixyPnxCaPo6EXADKH/k+MssUTqWyEszeW295HEUILsM4
exWvYsyzx7SwYQQahKdNBjiKSHFG0ZXHEdvFYQiyKqhtYzmAS0AZA1vh8ixMzUpg4UXv+eYFqz67
mPwp9i0DndOINRKiu+DVcyDtmswnl9aWuNFaUQbfI304tLVt0BtcklzCYgpQq0J4QgjagsNPflio
kNDRSJfgLVWHqd/VIx5lWEhLkM+y5fcFjrNj2+btjw6jzRPZ7lz7a5fzwxhr6PNcDfJaeEyAz4QT
vcNcFzP28o8RKSLksmx1C5xWCXqw5PVnMA6zaEyEDWFCBodts4NaSjIc5BtnfO9I8UjqBcY8s4Uk
8QHmdLvgfmqO+N/eW+z89FY279I6b7z4kQwLDTEpMewXHco3RH818VjTRpntwYRsu7piClSY6vXs
gYlME1iRsXVpOjQfp63Gj5TjXx4iaFFmh8EmHH9iGZRv5hMPRV/9e2EROFfRfo/ujxDT9/lUlWmx
ugI6vEYczrKraiIHTS0MM3GAmNduPduucNwpbEZkiQt7Ra+kEFe1QjInFGfgSN/HStLPHc0JnZip
6f0Bp9mqV23yIGvHjAwyuyCkViPQ5Fmj8LwFBLMTqcBGjcomlnwoH6WChlNFdsF1cKg/aj+kSgPz
NVdQYZX4Q3X47/2qP53670g0XhPR/Q7Wj+WjhLEeV86Gn19vhN0ILN1dlOvL9vWa6c19+ztULIZx
rgE8qo56+f72UNTUlxwL9RT0286kRQ6ikfT3jMy1U5Z6ykKfUpwZDInK8ypftyZetOOHCvyXvJwZ
HsxK6pq8rWLZZ4O6GH1tVF03t4Q7lIIXDWh1gy7nfXuthIMFfEWrwRTfBGKorh7so5V1zqXzgOTl
qk9/jWV4v4ptuhb/lB8tJXw873bp2+awiHTjg3vh4BPo535HNp5V7AULTQA/rjiI3dHqiY4B+u4Q
gWVT38KBZzaOqkUeK8ZXpBgOzAQWB7SCvL5OaiRVBiUHV5uLSPQltARLuh58ZqJXfyPky5PM1Ut/
LsU/YqX/Lw00N5tgO+uctSWXaG+2jwueUrG3StFSTc0Jd6Yr91i0XmcrivH2mFZjvKZKENegJi0F
A2fMuvMuy3AvDYJn9P6n31lJNuob8m9c9j86U2WJq/bB6bmrqGhYV6CfME71aJIIApZUGjusMlBL
V/ikRXcHJpQLY/TPBZSkwe2cIWysAP/4f7tPjWCJ9c83bD1mREbTdEZt+W5g8gUo0bVaxCfkjUJZ
REJwqH2f5wu+wjwUSYOfchIsdCbQQ/rIm1XtNF30YV74CpuuJbUiTkISsDArEfMxqCfeGZ01tykr
EUwUFAKi30lVKzCvLwk2mlpZQrH5tuUn4xctVFyyEmfyTYzG494JfMsYcET69p2Snhas42+wg19o
iCAG7rCDL8h5hikEvRWjFPPbTeosxufRcFIdc5CPruGT6AIkEY+2+/VrzKRh+xg3nzr/sQ2q7LMf
o8rt6hLCzkHYqesglAOUYkdUKQeogeMoJ1vWzqLs5XF+bbD/EBAAylrg0814yxo6zhicEYNvyEl5
K0KVlZczL+ilrcqrDFDqNs6Elg2mLAEsqhfciwGYX7sABcKvmWrZDNqw6P27bt0cePxlUIvDPUrk
XRsNO2WqsQBQW97eRAKMWeoNYA7wQoVwuVSZiwaXJEO2fQUKyAM8iKslf1OvK7AsiKEBJtmdTR4r
kzHT87Ssi86Or9OAfa5V8wQyK4GAiqi2wgi6nJNHazI3uFgCYtPgoSIRpjalVfHnF3iCzbXxgBST
qdWmjCHhDJEA95nf9uFVUljWI9wfKa5Hb8fdyf1/UicINPPxBtFoHexk3za6m3cduwHZ1dOM9oGK
DaOdNz3Em5jTZ91k3aRXOEguT16RqqZ6DPpm5f6UPYNuT6pEXgXFghTNdz7yo3NlW9pqQ1sbZuth
2rIUDO8BJMI9+dQU7PMlLxHGPO4oaj9mrszTpmXBJ9yQVdqYgLm3gKf6JzHSitG/ENyRoMDlmzIo
X8naQ4J3aZrIu7QTsJZ/U3nWsG5oMF4D60QmUFi6Bg0RLhnZR6utHTRxAPcgRMFwo3hrPY6opnKh
fnZTt/G9rWSjozkIjLuCSb4Y7hCPVS9s6XPtTAB5tKHUbkJ9Bwo8w74MtoAomYiKlzOk+GqsgUxH
CvXhhFWDgtFA0gZU3FuOO2LP0nxU0ilwhfi+aNUACu1KDCg8C+bN5Q3+FiwzNRyljd3kdKgDaKIA
I62+jHTOZH3Ubb+daOSZL6poMZ7OAqk14dPXEGJUDrGH4lRfO6c8y46XhRPfEo44S6rSacKeL2ta
i5zumBy+aa2voCnNy6DbH7suEy1Bf6eKzFE5pQBUoRH/XXbwqqk6C5iC5SiIfiF7WCyFXidiaGCi
NGVHuv1NBxZlhWnh4/Hv92uRbuN6AJqW9dhnTN980DwJCBUa5IM6inXEWhfA45girqw5OuwMOPBl
r/Z0lV0Wt3C/Z/cEyuAm+WqNiglHU30J0YozQunrnpa9S9ifPH1Ay/PuddikPox9TPIRaG4DkR8g
91fVRY4bA/9ooe7hGQGI3jtDSIh46ZTEugjKPRF9faQ3e8SQncM+3On1cj+Hf9p6g5HJceTnwhdI
+la2hvyPrHhaQ12CNtFHudunD+A/DiXT3XTIeb0AVD6aUXyJ7YIcY7T5bNsFbUolZY/+bOJu8G+k
CXxX0iWNpJxIgoZduG8zpXPgu94+We/cWv2zSdwFsq2ITT+SCdW22eH/Tj4Lzb+O5OvTg1v1v0P5
YMyvyugJllBmrzXOvD6IyM2Q9Ye7ooOZtQABcyNYUUKqSozgg7/9TrsgOJrjt2DIqyugGim8PueD
i+9PwFR8sSjrl1Bs1VY5rEdcm67JO+5zp0e02F+jSqIMrXRUsNJLrzVbZjBkjNzr3lV+ZpzvwVS9
LJhkE39CQoAcU8tp41p6dONaqubtYvEapYjuWYBGVaytNA0aXKkJiZwJyJUVeFc6XP9TneSeFt9V
y0wzcfksqXIwKm2H8C3S8QIquREhGEWtNwc2F1n0CubSXglFiot69tb55SXJxw1Xbx0akAVqy7Rx
Ioy5fhFmx9EPz8YfiIxMvA5LAcvqJ1Q9MUcMgtR7QC/gN1sRiX7KHol2m24sdnAjpOtjURxYWnEg
f9qCGzGgNccCjxvvcAgaO0gi8kNGq4qg3h6u7gppbDG9GH3uH9LW2P6WDZVMEHa90+NZ0xZj67H5
JMQtkScVk/DjW7C1QNoMqbPHyssw91HxYoSY1WewUrC1Yofp+HN9PvtjIrw5arli1t+XNfpQbs0W
s+NPYG0uVmByt2fC0U4QQ75aQ9FRXYmK5pqPvWkVqAy9eh7bmfhuIKT/VIoqwCL0FYNJX8/5z9sl
dvy4PxS00lgcx6mRVELf+E6pxFa0cLTYxVd1NVsZBdMZUacRlhCtd1K/zMb03lIxzylSzv4ZdaZT
l2578GsVhyeCLe4O/v97siQ1uS0tFqxIli1dAKPivfzXyqMrDSksrsUpsEBgYBI+aUJACr+vR8/P
nQe+mGBnwAuDmmsfRB3Fan+wKHZzfpSeeGQh3ly8ScsKqslXoXfZpn0O8Kw7eavWgosPnCJc82Xl
q5djjKOzjX+vPxsQkJpZtXU9SVw/OA/UbwKubKswW8hhzHSDR3oVq8ALxYzUMoDVCAtfFWFqKot6
5p4cGmUStO/BL/j/zCwMdxjMPsIyvdzd3ETwcZlC1tVDKlkhF3Z51Yk+/hHUOnZEB9aQtCzU7pBf
XWOlw5NBRvs+ywhChvCskvbGat9JYZQS8PoxbdWh33WfRRl9/ElSIcf6Z+wnMYKHLVAKrgbHdnsW
o0nVyH58z56wBKDNEVd8/ERICNYrkrxnxWnJsZNqm7vuyKLU6mT+kVz3CWsojckBIpr152kqoBFl
laCx2zm1qkMLzkirNYMBWSvZbmex29i7u7EAb72mQagVf6uflgvxS7Iomjx6QTXnqi5/fOmNXxzr
hqVKV946hU7Sa5FSiABSkeNZZ/BrUp75Qr+KKN7btHTO715/UEiQI2olbCAFkg9+l5ArAIFen0N/
EL1QHjG5U6/p9n1s800Ozb5IMZdcOboucy6kRzZB0vsGrt1stxp3yVicO+2VVe9bzwiVrfzgrGfB
gdG5+7AagqLJgD1m0qQC7xh8bKpunhJuKze4bIWXk58s7BA8sNURxLyx6crfbmFJ15CZUQaEzw+0
Y6q8baL0dwDGyf8M+83u+13hsbeHKPVyWR5QqWmYr9xdMNiRX5UeWY6NHmMKaz8bBKaSUrBWPggJ
O01pICEuaKgCqvZehyhYcwvX5ZiZ/MCJIzCs1NSMfnrvNKmYmMFhqVMrPoZD5DQUk5qHLjhIgeRm
BVam1tJYwCfeMsZ0XpwJ3LXa38RIdNHJRkNi4nhRBWz8us1YoEC/ATb3WMCrIiIc2eoTQFw421Cm
rrbDrAo2Tnpxe66cvmlhZSOPfHbhe8m1ADKwLssSkJKEEKsRW2EvuO5nxOdOFfZ+/isojDioQpJB
gTJpLAIyfiP3IcezSoA7jwxpdYVMcHMYGt9CXYh3vVrnXXYZONMivILsqN3zehuQJuHXfbF5xcm9
/vjmiQdiaZ/bm3ecuiX1xkBJmD+hJtEDriMQianZru3RYz0I13kcbPo7KVX2SHC6V9RkJUTOayTq
bc9PdbBWVZ20kk+iQueFJ3e54zFcyAzIeqZF3CrelZgDFCf+2F2IwshJMTtJl2c48coY+3W6ClTN
gyiZUztIqM1IQqDDcJXM3IQ2VV8Q4gYxHfaTfsbU78vBJty5A0S5f419wFuAL7KnIOzC6ZV7ZPgQ
7L5kGpNJUzG+wJ+mGeMj+2QQ42MRGwVrf0DoyMdKfNw1+PI2y7rmoxuV8RKVf31WDKE6uhsGV+Qw
Lb6WaQwpSkZw9sQG1FA7kO2Xa7meLzm38/DdyU38aNP8sR33lhNMKvwghScNqhZdcSyO15Lgttd7
ekjEWTZCQYmFD3Y6L2D8SR3l9tDXgHGfXPC7dCvV2K9/xsq5gBVxjWGedQel/vELe9aht2dgdpmN
1k9j0ngOn0MZZTpe7rUxGFUG2o5ttUc6x3EwqADNHHcCAyP3F1+4Q0BxXGpO6mwRDDHlEVC6vGaF
UxiYfRAccZ/T0cWQEFSl1OvMXwHoKzte6Gx6QQZPIHqtu2bCagzsTzqMLiTdA8b4tfJbeMkczdjr
TVzQsyTqUM6yYLrrDqEQi2U36LD6vL52QaTsDCiS2lGAEu+/KJxZaMeaAWGnRBo2DKHGo6PxU+uB
yqc18VZ+5XHOjBx+OYsEQOmrozbAfweCrkb6VBTEFuNoowCOfxxW2isCC07bP87A+pDnKghX6yTR
upWf49m2grpEq1BhL1AI854+QJxqZcl8qcWa8ySQLjfr8zZxE5VTFishIl+AEMrfD7crwbq6Qrun
fFLpg0wnXcT7BcYKu6WCKHGrRHYXhrTf5GX5ixF7g/5aQ9P33tZ5+tYeAhG5/S7BeJ6d92zrKouD
veRWhyjADw4qwjbK1efTlrNXEjGcNRWKYoibMc8NTxmIif+JNIgdwACWsNkonYwf2l2VGGfxwAXf
59GgPhywMIayirudY2xtaOtbCXcm3jYkniimNtpY9Vl3+wMOg0rbxIQu4ieBII62f9kontsApXk5
/yZjmjzJ968GsvTJjenjzTpwL1oV8bqC8B5gDzwjZJXrKWzfoaksrGIfIsT7GeMNnbhC9kfrUvoQ
h/1nbh4i6FaPwR/EJTbLBeU9hQNdY8EVG2/YmnkyYeRLWDnNbz5DpiW+VuZl7tkB0wM39xRB2LEb
+2l0NRB7I6Nw3iEMEmURCKWooY18vkHSqT4oH2qHiThxFsQ18rIneoBggcZCzjV4rE3dcqlUabRO
vDGBd0yT2QCAixd7gSxyjU5U/mMt8wAPDzmODXH3iizZkFzWPtPNYgnNmmuqjwRgLoh2Mhu0JG5O
yK/aK0HTq02c4ryuSozLQHgJDBfUQOzo9XSckWNMI6vpCULUTf7DxWPtwKkWBsXOt0dc9N9IKge1
ErfT3tlQHmDu4uEyKm7Y2zUcE+7TJcjNPXQwJCcrN8xOXwTdB1TygTPxnli38L/E6GAqbHj4CDEp
NwcgjjnBPmHXSfHgUvdWQPC1ER3zbk5bfyMLXoG811aBnGS3fjOMImNhKJA3esgOuT+oqgYaN+tj
PpjHDgJsVzneI0ByxrHxwZWaENuRAy/vmG2neF5w7r/g70DSfCnhgKFLJfpkM5exoagnkmSS4DGd
UlCwXXBdKGo7kUIdhJ11vB2iNIamAIdXQvVrdF9SqDaEy71ik0CWuF4H7TRy7Ta34vWcW0oNmmcL
XRlzGbOtF0PPN7UCahFqoxCsO4MxtzZfoD+oLcGbus/1WrNkDmJ77m387iNRqkxlpkU7lroyNK0N
6zrrfZZn8vrbAb1k+rvkCv2794WwOAyaisqqsSV5DBLodGYyTUVEFYttMfIBwynebqcNKw7+S+3g
xghLZqafiHp7wv1l+PmIu3Pr/5+jjSoCZ+sVNewP0MJvNM63Nj9dCcVvLejhNidlU4iDH0YJjjJg
WsTJtNMsDQ3xhFfi7RMeGGljxBMMo097hTvKdgEE95y4CoMG8si+Cq4lvLcqcin7NLqj3mgvDjU4
19tUdz3svv+oamQityq7h1PvQIDIuG9n7ydzQUT2Bi2jmw0ESBgmKlcWwLiBHHLEOmIafNW+RYAc
4i9KQbAkbP4IwoOC/JmyAhjr1XgkEmtKIqUCV7+Zn8LjHJaMwVOKhOFy6uww+jPllj3LVDgmeNoO
9DLgTHgPm8lAFN7EJxD53sCao+NIbeSbCskvlV6leVjvVvDiFYNC+0lchh5CN0HZ7XN5DB+uWUhr
xesU30nIU5n7q4ERRCJdyJU1ggl0iBiaobMXcbRx5fMeUpxuklZN9xV0eTnSjA1apV8AmFTL1YD9
1UrIzEJ+SU1dDVKcpw6k+ZgTw3ESdV0bIxwLocljE3e4plWH9idPtFFT0oxuSOqdsonGMUQLqeyh
sw2ahnJXSMeeBPCWhwMGIGfWHJDaF5Vkhi36/Xjldpq1v0pRZdJNsj7pdR92At7JSodBVSPEgnuR
cXuWYScwmGmpGookA/QT+mq+HovzS2RLz+Cq9OvIlHPjsMDOYVsAHGZcWpBRs38GH+kW+ScF3c76
aK7MHdDShnx3lYw2bFFcUE0h/C5i4LnOl98LP3X2ziAgZlmZL1yP2jyj/Zqkzq11MSLzHTyLsg7m
8ty1y1w92xYWIgxDy4Htk7rxi8rMesOTRXWbsuMLaWw1o/o8Agg5lQ0+ILKZCkDY/7Rhom0FTJAr
UQVGqWrBAsgpTC7c8S44AHR+ZO6MbLLsOYSSqZZt9f9hrqsAlB0tBsmTCNy181+fEMdkxo0mynrr
q9B83EKOcwKOoqARX6HAk1w3RbSAQMJ+Ml1YSqKPzhzPGQR714peF3KAQl7CV4uY5m3FtP45s05K
W/G2ic/gQBMW4hbAeFD9ohLR/V8mS5H4TZuJv9L6ju7px3xfKf55z3TByFY/ywSX67+hjf9hwLMx
le72jcmgMHSlrp7/jq+QFfHJ8oWkkYNWdaH3ffz3C+gmrGsOEXDOgje4n2W9YhV/v3ONoVNn+Nt+
HwN1xTrBpdLyeoGreQgGzw3MdqYDhcb/v+nTlEBW0umjOuLBFT4mN8egkpq5i6F8A1fGR/+7AAhX
KG/sJ1I/prJ3hUKKzaItaecf3/GfT4+oeu52Fk6pQwCaw+sdTHcRjSoNLBbl9MBNc73Lk7HH72Rl
npLmv0dFnC47ul9dFAvmXTzNQvmILvNVmABe2c6jXEbPOcQdNz3cQMFJsR7WhDfnvqnEcCzmtqhm
c2K/WoZhPI+qQYygvdzZqt+Ui121zKJk6OZPRVq8AqV9AdJP/RByrrzIGBGAIV/0fM6actca6ZC5
9gTbkSHqv2E+mUfDTAxqUdO44H1w+HZwiyx+BKRBXJPkNzQUyPduweM0Z1HF4b9OQzZH4luR2YPi
/ltbzy5UKYWODFza4Ta8BCMulhvxizgj9wwKnb4V7fijr71TgrBShF+bQ7uZ4mT2GaXwa7g5crq0
ytbp+kg2QLm3TN+Buz/HqrAs0Z/beW2oit0zSEVoX5SeNiSkBanWURGhoiquZNp4wa3QDf29LMjw
6Ey8I0UAtTiZjvQizMtmSOk4rR4silBip+wIxWnRoYyJSSk/0f8aO9+lJRYd+7PcAduSSokJLQpk
XqF97A7jgFlFTCaq+coEhM5BH9AvUSYw7GilspRsN5/cx4vjloM9o28UevoVP7SpwCBeg2RdRe3l
DyrvkeKNzAwLUXmxF6mlUDtC9ze16T2lJc1wCEOUm1/v2yKZE/K6qGDMlchAOM0aMtVuNMQ+nDTY
x0u+OUbwYzssqdWmOFVnh9+7lbwJL3ASFVjtj/DoobV1KMwRSqyMadhb4jDCo3VLP6ByN0VReIZ5
f1SAdi/exn7tDzVQoNMou8UCvgSK9/aa9UhwRtExbpOgmV+3GqF5V3CU52OreZuqXJLLQuLOHU9o
oeSWupmeOmhIV4Ic3dq8lSoSLmqX6SKkrgjx6FEM6MNxwUx9Tm/45vwn2WO9qApG/58WUlS5wg1n
fwmDCbOiGvl4BXMCbdbr6b2HuuV9Y+eBjMGgUvqg0RKi/sfuo1iJcHPNh6G/WoyTgKdCHUXUwE2d
xFv9viMIpGqRls1p4STZH39Fs8dbfj7x9qaFA8Bn2WWMxOUObdxvss7EcQAAtF+6wpv6E2kbsWrv
pARfXvJMZRe33VcXPTsx2GfXEnIBDGDFd3uvCGe4KWOHCiYoTylMEkZkq+UUSlY0/DfE3BealJ2h
+/gplbnxhleIu4bCUUfmmRbq0oStvObPApDug1KvHWxfK1xAeOZ2abzgHKcYzqjTXeHaX+OluLrc
vs5l06JkJn1bD1sRIaVcpmiEMd6iG/onfTBLT6ljFRq13d6eab7vAk+CcBwIdFuLHeO9vH00q1c2
S9oLWurAy3JDrXeMAwQ9A3q+LMlJnes2tzKi3rn77R5T3U6F+n/5/Jec1eGbjgLFyOTnax1NHSR/
d1fCDzLD48tGjV+ixgkWumjE69pyoPDzD0hbvB+cGEwLegAexpAEg4kMu+oSKS+w2opH6uQa3IGm
hwisN4KFmRrYkUYouV8Meft4a25QzUxbWXdP+OJCXCKvrwA6Dtt9btaNaX4vfVzfYId/Grph0O+H
T+5L+7xsbWyi7JcyNaqh2vNdh3p4GDkJia9GOLjbjizN2KPQjzz+ftnTxieEnTatICavPedGRgKB
gytPY3zuKU5P8kfYA++kGuQv1dVGIC/KnOHN4PnUA88Y0Vi3DvFP+uCG11phajPLe09x5Q28bimt
U9UpcMvB75Wl464OgH+iHp3CJH5WJydkTbzHuXsXUGOMwHbtZrYfxOCLC8f7tPfNvho1kEHRG9kT
+M+7qodoSd0850ZNm2AGeYXsl15NaEf9Vz6vnWJ1GtW0fud9qGuVgSwf5NXvOnW3h+KSrip33SIP
pNIQykEljjD+tCZHzVHQldpA0GBIcoak8FZo7C4S55QpWIf8hOUcm4BwPsxxtut5tVxPC9CB72OR
WSJbERBxzq1BncpdCrDiiOCSEMtZWintHoyAwn+y8Md7uz2/x19UU2fZK+olcbLz/yXuXZWAoOtx
2y4bQMY0HevXf/eHCZBkeEhtYLplC/6H/F23QgkusCWhK/tRJh9LlHb46DpGxvbIlCeku5qGZK73
XQN+kxqcs9VPTIYXEReyGoiPHmQ7KXR//124V5KLBGwcpA2BRxpUVa+1DmGOcwhSZHJuuO0lcgEY
T5IdAL0XRlqvb0cCivks4a4yaa5/xpmRNnKmxXxojTr+iTu7gnc1I0LODWFPxq4FjrLAdBDleF2P
2taHloe6fweycUPna04/W7bKJJzr+5dAjptF1Zv1Hl+qvWCWg/Xdyou2hgdktv7tIwXp2M8ufZlx
kSQl/wl9/cRFzKy1xy1QEaK2LOt4leek0gILoxWCLacg3aU+rFxuhgd3zzqf/lmilvp8mKvEOaQ8
eQXRuUFnl583e6DJWyiIIlNekbuLjbTyMGCaBz8GuJhWLjPtp74ksHCP48/ab0kUlzrXn94ffwoJ
g1AM14YakV555KUPW/NhEzWG957fpWD6b7LTBG6XTydF6rO1Kwp0uXmEpSThFhjhZk5veqaHfm/B
Pr/0MwtZKd6y3l1bCJfG01xL2wERV5YsmZOW6q24kE+qHqXZPxcIEbeBcyvhurhJF7pGL5lTXb67
HuAeKgluzKxpYDc/wQLjXiMHceUw/tGhk72Bfp0ByCyCB34MRiMKGX3XZLnUk79oS+p37NNKTsGM
nys952HMtHsFOt76DniEwsdOOkN/H60K2lvfU6I7e/S7rG5xbq+G6BmBXVw/A4crYkKb23jnWjgj
ua3maeVYBOTL7yTl4WvvOwWtt7CKmmOpEmmepE1Fx4BDs+5q1EBG5fwsioGEVDvj7KeN9t9q2RFh
tZK1emEA52qzQsVYWe/Xiz6mGCwq6eNU1fEVdMw+N0aUhHnnDGNYy7JXLAO8sCVUxfau3wNWdeh9
jRBalsGXu8KnLE5G1BStw+q6GuiCWIn0FlluYz5a0JzvhvzHa4Mwv89H02VXwBhVRnD6I36Hwhpo
hY5ggYdrI/fs1DgOO7IfmA/zffY4MzLVd0su5GHAvC3PM6JcVm7rCeyBS65FzBlxW2fcIEVhZGnw
pJIvwRd0WfH24wZ0Mu1oHpYY9V05U91WO9LpzEo5X9mJvcraz7N6Om70rKwWlmqTOFupx/OO0Mta
jPhYjZNE1tXrLDgg/O03+29tKD/yu8XSicZqPXXHNzppZXXTqCBV8rHAgwlVUgrDjs+GFbAMv/y0
sNgW7WTqLurLgAbeIRv9+EppFeAMgZtOF7hg4fUJbP1qUbQJuZbKfHDfhXWbElEwykdPmJBRQm1J
d3jmUJG16qCKuKGgbMDlQWJZdo8hrUtoKY8C7/JllRp2oowdI0T6KmEEqp4Vgp9xl9TQy8IZjOxa
8XL736m8E9Oi6tqr3hpMSrqLlhM8YnQWCGuxBxXn6cYKfvqreL6IFPdpEY+s+Ym42JM57OuqCAjQ
rHXS70xWjp8o+VoFrKJeWrA0gNC0hZ0F6Rdwl0YZ1vXaKSjfH4AWoqP8CkiacmArwYJt/+gMMUti
HpRWBW89aHIhXCGppM5m6BUPHQ0aAccsP6TbHQAN25qtkeK4OQZMlSLGeR9l4jIYOWWHY5O9kGeH
LVRHEaeQNYMx+RxuEMNYZR6j7OZp4sdVafpd/76a3drxCzQ3D08Zcf3Q2b/SaAScBTPpbUs9BmyI
ORA/Qubi4jsCfhpQqPOGZpnbHip3xeMcIQDHYkCArHHsKacONRl8fYfZURve5ulDgQcNDEvzXBBA
zjGcVSGyprZB37cDfhyrNxBn85GVR4xxLDcDXgjmfh91WjVQUIJz0H5ry+yfs+ch4zY2Dg8kcBiH
Q3MHlfoM3UgWO0+e5q2KEgQDAVl4J7AkNmMJ83Bqs3lIX1SAoZmv/CXw0PGFEw7RPyTdxpC1YTO3
lwBddWRWBU1REj3XChvWt+pWiy2bGlZLQBR5LdN/MkoShTspi1Bt09EkzuHy1DSIcINcpB/8ztRs
oMkorC2hID7fsgCYTEtwsR2meiEpcIzPrFXGgzK+H5YHbfk96IYhkUUddOMa7OtUjRh4jOCdqgmD
D406Vn2l7QgA/mgKAGLPHmKnq6dV1zOWIXiCYpFa+7BAysiGjKukhmImvZVPsLci9ks6mhPmgYMx
SVT3sNR4XTCiBbxUwNOUuFJgjkro/bmJ7RziC7Ml7fgP6suoHhDC2LvLai2waJapSkROBtCoQVPw
5wbPQqx1j3TOIk+T1Cz3L7Ty0Y+20Su2QPXUAFjH4kzeTXQM6cayggJDSzV34ZjJAISO3elN1C5u
4eInrSAIGFoBrrzA9it2qvZ6cgPbb5dZ9oWjJSHqhryccltb6oknn2KzzvwHvOzu3EjkVyIsYWlJ
INpn+A+hUy/NWLBysSJR3Ddj/XmyZXuRRKMicZdd+pehAJSZRqh/a7+oTv+eS8vaUegUMwPxhOFQ
ve2pXUN2YRooLjIOORqWuyopPj8LO0/jogXM2kN1IcUYCgF+f0elIXmZL25k6QjkWXsbW/cE3PY5
JEceoZiOk1p9J/K9ojfUd3Nmkk5ZZLrMxDGwBCX6DHC+whsPC7RCICzj4WsK5AKba4FfKBX7BEBm
ZwvLLO1WRTx2Urzm+pwq26BZwIZK38N3No6ilYDWet8CnVoGDxO4Gvv5tx9aoao9rNMJwI+ClHPp
DM//pf+HcQYQ9vu9s/YrZlTosOn/VwOkSKjg2tx9MCGGlDTbcNC7DBfsFCu8xRtzqSAWLFKaiZsa
Kse7qVD1DSfL4KMnig+zV9oVxJYZBmBv7tA6EuJtGX8Ko5rv82hV/OIFVR4JaWDJcGYqL+XtrNpY
jRZJgTn+/9CW5am9P8uGioiK4HFavhO3SQfiylqbcXDz4nsGNV6Y96KM9vy9LQuzuy3ilENYOI6T
gCXSHCp44PRwxzo7l+sUFUWOsiR8TTNugmFGxpsej5RhTSjxlwJ6WgRpdCS7lNsyzwaQ8kgARFFr
Yjqhb0cu1W3gDOEzCyOZSVB9jnZjf1hDfLt+iDwhCERgtVwDAddiy28mHK7BDdr5HB7bPep8mHd+
AMZrsQiv6mqCAzmzcqGnjnN2TTWNeJ1uqNmWlzLirf8B2D+YHHY6zg+Iui5qojV7t6b9NE8t/33N
wV7bNFrWNhnvpqHKHu1QHmPyzyJH5Mx8Zt4SQzL7OARx57GU3kigrX/FyRmfGX55oDAMLAWWpTuX
+FrP/QrCcYtujybvIzujyroyS5dvZX659Pe02vTiRIAL5PszN024+OW3phH8P62Eqv/AyZswshyB
4apB23A/5j50Y4PlSt6ycBPZ1t1Ye6JndTPi0vu7z7FnRjgwOGGL95bL22pTKDD2IsFzgxr3YJ0i
SCQ8s2OOeHL2p5i+HRP+HG9P2h3zBEWI1qGcsEj9R8qbWWjx4D5MFzELGyltWzfMGsrAnUKm/HmT
Mt9eRWpFRcnqBcTNWeDCt3ebTiDk0wovmXB4HZTnoac4rSeAAqRGVjIiblqjP3fbmzub4oZSLgrj
JIAJATglWn/LIVI/w8xe6azy/xWY/6nohmfCwlp8ue3BhxgqFzz3ln00UDlnGq/+bZu56Pnb/wx5
0FIgtr1cVBWRApXy/jTU2gWdvFVxghSQKoLkPSaO6n69Og5rjkOHFnfHfWuC8KkkbddxShyJgBGG
qnKquD66uRNveDGxHtkuLIgcm6s9kJiFtr7GeEMI4/fiO8G/oUdWPBSu4D3Ijr7HTerr8Si6G8Kd
c4ySv3TfWyZAWQ17tBC4x6dA0giVky5C2z/5TxkZ+fSM+ft/KQVC+CDzjC9TuiDpIHEMngkT0FlT
QJnOJjC615CIu3xnSSgeQqxXT0LZ/CPCAXDLh25qMf2PVFG+5wUbZnZS0dP09V7yxAWFJYl2CXZm
UZq4usu752B4rQNTFUW0yKGBfBn47qOGdvsgBjwqHiFw0Qxi4M3mlg6R++SfrOP5jbEZ5PgH7abB
+ZjcmLXv6IxZxrARlG1JygyhmIuUbljP9PMmqKIGM4SlEjyAfuoKGJw6y4UHepmaoGiED4R8yCTA
M36mqHqsgmmxO4IgWvZmQ73kxpTzJIxgJWhCIUzkZmsV1geUiAPXAAmLxCAtcPn4o3M9R0hRjXQE
nJ+DwKt2xEnKQkcRwFYLTjo/KnWEk+SsOAEyKHiCNaBsNj0di+3Wp4IzZR2Qz5BfiqwLzUveRFPl
IEPHLtEN2FIUoC04AIjzh2vSwC0SsqbsxxQM0tqa/a7FRGp0KVVfgPKN1plMiP0xvSLERQvqxIBq
PPjUhNIWdgxcOznxKk5DX8HNWfmU7p1Psw8KIy7UijsEnIF2d270uVlW1yaKntV8a0ooyPqVsJZ5
LSjBByROq2Ck1FtnGy4c5HcKkmwjvDI6WMmLG6c7i3arFx5Y/CDRalpABm+OvMuT09BDjM0saLax
7fa9HFoWPmM7ITlxbSErUW9zIAg0D5JtxEp0mRMPnwtfWcNhw8Y3scoGdA7rsfbINtoyKl+ZgXW4
MAuow9Js8eNHYbHLSr8TbbQtYy56p7QEHTDwTzzH5oVxWDzX4lGNkGaRfqH8yW3Ae1GWb4Bdl1a9
/dIye1ujX+QM2O9NxEnmeZ5Jj/e0dtHhFR3mawWOpxXDRSTclfWtSh++wqnLg6fzk3rGuVkWwKXE
T5vB0BzHei8/AigLWNjwWWSxa1tu6p22ttRJm23i/88mr5kPgfEgZzSzylAGEgB7ZJ34P7MCM6oV
j/J7sFyPDEhgoi8yclWjAbKrLl9Wi+TCmG4Io6f1jFYX4wg8zycyU0qixa/N1UvedAsJfAOA0R+P
NzScTG2sf2Ep0X5xgBMxbgdjcmjDfWl/vFGUSh+vKOVPWTgrxj4mzYKgel31brsWxPzQwdDS6L6p
/0cusFULbE6RBJp5LnkbYmDZnsN8i2sGIJr5zAcSl+5sLWzEYTAFLQaYwK2bqUC37gQT53bsw9YD
WQXrY++fPQ+FV2jYmyn6Lw4zYtS6y9ZJ/Ij8Zt6ydE73jLKq3qbjwcmrBxyEADWeUc5b6lbTprD8
o25ksHXCGP4v7CO92MzfSqvc9NtgHOZqVL/ZDFcVJ6JtZe4rIP1O9R5wdGe1sLk8ZRwBVNAa80/p
DTTcWnhl8iILb+w6lqL51wzZdBoPqo37skclBOg587pqcuCQMDg88zs6oEjtIbgKy9aF4lYrL+Sy
XD5X5nE/QNTUyTPLhuNc0xaOjLqVzLaOF7Fm8LohHgDNchV0ZKi4OQuDzOXFJ1TFf7QTGAO+fcWq
LV5xhgYeoPEK5Y8oQqaKWUD/qEYUL0/hHmxIWkwoV4MIX3TcS7FVgGA/ygyiB3SPLdBsFxWbCZCl
xygd0PeWVNbMzfQypsCk51blX28NPEMiOPUtEWnMldqR5A/hMkZAui2EPT/HDb97EvIGGT/5ErSE
uvrGPu+gSrvIHqyMcnhxroPL+Zul0KuOu9+2vmMgFC47w1WnxJ7IyeU00SYcQC9OptJOjXYcHrhA
EFSVAW0ioZwAweE5lNYn8CGriQleOA0GuUCimukavxniryw6czWYYCBJb+ASLh/QR2qXhRfRLxQ9
QFYWM5EqLWRT9NnVWSehp3NmVqfKpYZw9P/v0SvrZn3t0OUGUk1Pade1hjzYwf82xjemxY6wzsFQ
ZQmjOpWYxFngzHnegSqsm6/APQJKggKNDxUisHgVner2tt90X3faDwk96O5YBFi9aWpwwnK/Iciu
Cg5RkIZG/4BODkcmeF2eonwsXUKqsFaUjHghb6fd5IAOjINFXTFJtLS2TcSNkrl8SOJ7Ig5VJf5q
Tp8itIevGWG8CvpgEumw5ZoEbfHc/bZh06LXPCYfywhE180Sd/caA9f/hcpV5bdwgykfCKUUQPPU
hMobtwidYVU9zneFBNNBXBA7rl1MlKoF/5vz+SkLask/IP2micdUKu49vneWQaBLGM82d35G3RTp
zkKedYrojB9E/bfg2+Ht3KeA/+2+BPTw+g1RV6CPZjcjL2SP1AAC1F9HQ6T4JKYVo/WB5hghmG9B
Uo9xdNVUO3U6XyWKjJ+xxlu+Saz1EVIsolX8nhEBbT6giOsGyi4Pp9nx002mhse7V+yN588OSAyv
nJcwdCUSifFNML2/dikqQqWCdmV3PbzUmqCiaSAbra0XmSpNZyyZGf5srE0AxaOl7unHXPDaqj1S
QMcDNqkaL8G/G2KNL1SEfpgiHT2iPvWDepBvrWh5/QtX0R9V2LiP+53pZVLfwIcME60mIba8ohCh
4GXuiZxO7IU0YV9JsQr3OBd9k4mYG6vvaUJ421FIHWO9ALoOQE4Ds6EldZ74wUNdzzE3zSPF/IYz
5LScCvtdj0Mj7mS+s+0ierceyOshTI4uq9TXiKyE2tA9YdNykUXWAih8jNW9J+201QbB+bOFWBSs
jyhOzqIoC71fowu1rkxOrNQhqGt5uxh9AXHznVyPnyeZFRQsziyzwDJdv3cdWA8Wzdbw7aT1g2sj
2vn7GZDXQRU9tkQhC9TgS80rcFNb+b7RPeQeYgwR+YyZsL+IWJbQXXv5HnyxvSO0upAD2KvaewaJ
AJRbLpUXG/N8rf4yc041ug/voW1tzy1k0S69TeYXPu/scgLZLbNHWSOCpcC07nFgvOquCbYg/rgl
a7GNq7intBWhyEQ9+tEWyJexJE/mDaLdvdocXxuxc+lZQltIKR7xtiRHHmOvaSxpWstwhvD2Aezf
KEeHgMDHFW0luXKNZB2Rit07KmeXaUTLRe4R22O0b8jVQbfjwJW05cnG5SKL0eLxudTAZK9MxU5I
oaI53T8L+yarj1H66tce6tDCOV9YW5VQTXuYLvGB8YxwDelLC4Yhp93V28L0azGNn5/dlffqcyaU
MuilrcFevjx7YWQgWaPJ+Ia0NfD3K5AnyQlf0Lp+T7RyUOVbgtqW+f0I+0JOQteBOwKBRgiCq47Y
nflVKg0BqU+t2v5ZyCZOvRuB2WbX4qsb2eqFDHaD9ig0VfSikA9j1Oa2AEaebmxuQFgvi+aFD90P
R6lEhy1WezDnW9lclwpDXn6SNolDruqBBfQnk6ZTRan+eRKLRDEO0j1dl1YrJQArpUFX0eFfr6tI
Svt2AO7ZgMylOfyHlMafqReTVmE2g75BInwUdkgqJAFI/beELCxJ9gYWdSu78FO9/13uZLsuGWSp
Mlit4wmSsbJ4QKwyutHGsa/THAmErLBvg/vTLamWLTe4HULODc30fgmofcOj6Ciss36Rpzij8YEr
wJlRi2RRkX75yGC1YBIj9D7ao8UuxlYeUjqrP5vUqCskZhC9OFhk1ijQDhs0ISJ1ViQrsOqNE+HN
PYAVyUGHl/2Y5+4S9TDuKOe9SyOzLvY/E7u0HFtmYZP1PwnUYpjrNgtgvEPtmrqdFTKCxFksSueC
Q8EK6q5wPxDAaxD3wVR4u4hsbDiq4UggIuQoz2NRwJ6Y0Vx/E9t9r6lbpcgWbxnRlHbUfIME4oN8
FbVIwJRoPbkn/+Uo2fO+lExCKzWbwXxbEUACAaS4PbhCFNmF62vPUUi+/Y6YV/xxAqoD0wuuHWBn
b7nElQKQVGhngmK46/R5zlWoypOJh8kixQIuwDPryMldX0w+2LKzvDtaYh36v1lLSGG3gNTKTg9s
LocNrdEZOmu6Fo6xGN2yLkIacYy+mnRbSLJ5BMU69tXz3iR+c6oMWiijlduX5r04bosxVns7XkyB
k28edLSZFYql6Gir77s1iiChJdoZVjtVHA1caJyUJzjTWvYppll7SHTk2llScfYgakkEda60LOmq
FO/AbfMnW88RNIG+/zL0H8E6KTEac3/gWeh9xzkaJk1rx32IlYKX5p63w/310A/4+asItsBK+nT4
aiCrpoi8l9eEtXxdssAmtn5olxxW9AClSIdygXFyPZTCyrB3hz0D5oZefy9qve/WydnCON9F1lKf
AaF5YHw2lWZB8l26e/9v66c/M/EBc58zXcIrcs3x50RQmSq3DHRbZPjrtqRZnEwPLRNYmfyayONj
X9Cxh/xXtxnuWvfhZq3xLFlqjeuJ4IO00qhbYfC4DMOy2mhV6JTvbEpi9hkVq+7O4iWqGmLXw6PK
23E799npcWxZkLqaJKGyToTHAz1/NzNh5/oi25bVfoS6ZafnfMAhED5Hmjxq5+RTeD1eEa+ijVyy
mUcdipjVA2OFG08Di50sB04Xk6ARR2ydavoARNl1hruc402OVIX5iebL5wX790A7TYPT2mdA89tE
z6SFh+r6bbo6QN1eGiVzzC+3u0PtP1g7q/NS5mPr0kA1CXUJIT4UyIQcEMHs7qh4o2MJfGBykXr8
xIDh0G3I2zu+JP3gMPoB0g+JA3uxLurj/A5t2Q0h413VeOVPDaIqL2usnXuvFGv0tfiGc0Aog4AZ
H0LBpeDkzIdAekNBuZJs7/AM/paFU89iNaZ3KDC8dp1wZ6wMPtXo/ac8n8XLUL7DqgYWY+Lb52Gr
jHrU7UEFPrC4nvu4jcK41sMXM62YhCI0UZJFOch3C061LtUYB/++fu7iliEFQ3/7lUWUmFI0+84Z
3AMsOdjJhs8Ica6pONu0jwr6MwTbLWnfBVNYVVU9nSuwBxLSbOlq4GgTWcQPalN8/rmLJgGwBlGn
xJ2Z+5Jbmha/L8GwZEbTLRV2cCYhDksMb6ftCFwFJ3f0av8FpbC0BZI/+Sow/W5+Zr2Yt1hE88/h
jwyijyA53zdJZNhVpTWeu7H2ioeiZrjwEt6W1yjxfw+fhQvnKnY8g1LQjpwFxpE8446W255+2ION
hbA+DHBoui0SNKzw0eC38sB48fmoPGhREZ+FigvYUcUwk1ClwGq7KSwOh2pq6E7Olv71Ux7dRbGw
sRPZkntGTpiqv58L/LFpLG1TGqN5sk754d+YuKt+PcEejSlkorRNObqUplmemRFVFY9QT0WKZpjF
ksojnwlwyu6MpV57qMRAwSBQHX0vSmf8bIiBJEwzwPzrTYo2mgwMSWHny0JZopOqqw9UHPEgoPtT
0UtZae/x5QfcQddXmA5OFKetGDn5vU8/JnRMwC9s+m77ItUfHTs/uqWqFAh8nUqPGJaq9gPOarjD
4MgCn+Vf3KIdteDLu7AZnOONJMG04b5QbMmcfKsfAc+FiOn7eeI/fK/1xiWLWcwaMBzP41AdMAli
UTpksaZ2JNcnWWrvdTbwKnWTGixp6AZmYAkL9b2UuL/gnVp6NMsp1OFEw/X824TAA6qcIVGpXD/w
ptGxE7+wvrG/wZuS9QN6I6G2Hsk4MGNFyMG6SAg+POlf65/Tj+HVOfxwEFIPXHLIrmX/xZci+i+3
AboBqV+sR/vVqNmje9QwR4D4Qrdd18ip3QbHAF0f1Lt1siKiuIBBCRysb5ZaNsojsPPR+eRriP7f
AswUaV7Gd7EpkcKYe5gEE7TlZr4rBn5ho4KdXhw8C+R3G/xahItYTGXM5iquzK+3Pd+tx0IzOXAA
+SJgmpyBHhJ9Y1RolUTohxpwM3tsYbVd08ss1uV5EOfKvPHbgkAy7DUnrQ8qS68InyWriC4uRhZv
ZTD9mWYb4hF2tL4ESSINuiNX8PI3mxDE14x9VEz37f0eGl0LcyJLwgFdKc3GRvSSqjYy5+znlrOS
G/wR+fZdka5hnczfEePYYWul4ssH4dQR8YZKMro3g+QUiRg+s5a/36aEWbalqFdAArmhbz66DOM5
AKU53Fra2Jy4TE13ItNzQlfKPwbWpSITVHvtt+Y7KnSFknSzGnX1L/yni9Qk4RVoyCK+47q1B972
ujfFyMrTy7paei855yngwXgxM0got5SxIAzbgDMFtc88h7F33jQwc+6CXCfQJnWOKhtIjkFow9Dc
hHV4beWbWIshj+Grv/FYVEkotYPNggXegMZIJOY+ra5kRgPySxIERMehabSIFd3VJ3he79fR4EXf
+FRdA64uyjIAh057YwOdLNywGj15E+4RVCA78BiOno6K2ghomc6eyQti5lO0mZlkKa4Cf+va+K75
bzs/Fl7l0XbTtGzjzugpRHR+fKtlLRkQtaUXwuRTKEUGRq3wFROHl+MXf/cI6y+P2U+tM8juJ30v
keFXa1mZdvVq/9Ty53pJ/F7K3hGEFHmzagyWLhVdnMmR8lnZVFfldOUOzhxUC8CYRNoSuwgj75Iw
bwThJU0HwcPPs1E8zvSmpYxo+QAmrlcXX8ZWAwuyZ8cXD9novM2bt2Im9DboHoiZrIR3IV8+j0qh
mjg2bHqjBMnRMCTpHfgqAqARLnvVrqtqipkzwyoWsMk22zXB19SI1FhQu1drp3Gg1PeTVJ+pDs61
cQ4PSxUGuV4Fwrh/F+q8SbDZOVLWkGwmamMQ/Z1foosn2MdnN3kvVdi7IsDvywYudbKtd984x1Wo
x+etSAhf/khV+xoHbF6N6kpIWJwNNezlgwJIF3aMciVXj0U4XGDlXRM53hFht5qE1z/Ww0PoVFPw
5waxTOwnF6iJeaR55WF/JxoTn8iAw9vjRJys0S6VlsFSYwak4nCmp8uUfMDjLbjX9br4C2ZwZ742
r3G8DhN9SZMrz1MJErpsuuLICw2CLm6NRwoPVTPYk5NjEikSh/wZotaJSoKybYqXsCtbh+ExYyN6
4bI6GJzpLUDtYtb0R4QdAF5nh1gOTvRHpd5yqRM87OqNLu9pgS/QUOt5g1klAR6ZRv/cJgCoD8cT
mOgVzBclJ6ZcWl07kNXcln3AiZZCzVhhb905Xx3j+zO0S/vw/ppCmNuLZ4a2+vD+cQbzPZHErksz
PihcoaGO0DhaE0PIYkggskhZ+EGp0zozsZ9vSPg4qWKbSeVSAKfvBc7XMRNoy+5gjZDf8yOhARQD
30qKQxClWq4oM0aJXG+0YTPX7JHOuK+hF8Pr1Ek8jIXHfoK2s6U8VqpnUF/k1eedCRCiu/C4K9/1
S+w1nQ7tBtZIt5lzg1MCxeoF62bwWhyN6v/G6sTYGmbbWze2fxbmECW8lyDobL9uvyGNA6xuVLYd
tuqv5umhZNDZ33jGPPx/w+sEfE5xsobfyEZQG+uzL1lesdZhMMok+HvsRwTB6aDfyfb3Cnpo/HK0
IN+oOfCg/hMTzEYATL7Gip/Fvvuef31a3/kQSuMlbkwBvEPQu7y0CyXdPHuZgirOGhhQNW/0mGiS
+i6fn+FagzuJLLv4rWiw1UXIJmbQupgGkfM44hTKTSK0ZHS52vGDO4UuZxVTY4WrnoJguoArI/nM
9klGOFAipC+/8iiEK2Cc5wUQVHCc16gIN8+UdM3bh5Rw3wb/QVpQeuj5dB3+RilRVzdOrgablkwR
dEsc8xRNgHp4++sN4fn6CH6pvkN2hfWpcSCZ+MHq9QM86hqszHGTXa+rlyRazPBaGRqJMboYhMu2
ZfpJ9MDYk+N459Fdc2gbvYD0G+BFaKh8wsG+pINOO3JxPOdZUT5Ep+snKcSPkn1rZ5u5IjFiMuBO
gRX2txxm95KphkjheaI7k4LMZUQOCpnPnzawT4Eek67G4hjAhVDqRBMdax5PCTmwCgG0bIvex1Tq
pe/fkQ/bApBAT71WJhnWFWLMmPOzwf2I943XuYjYcmg8W1ijViO05oz+vFOJXGeIR6oeQ/pBGqva
ZTYLKnLi2apy6ixvdDrFq6MdRFe/T9LK0cRbFwRTht5e4MJQPC507Q5eywlAhC664ePGVDlVA+EK
x/jDTGORtpyIpPTYul5bF4M+hnQYU3Jj55rS+q8Aysp6GluBtkwmrXJFZ88sa0jn/JK01OqzIMRi
VH+Cp7xlMafHMRYMsy7icbUtj2YvdwjmbE1YBnCFFp8EZ7TeXYkAQX6N3z+pPdzMr8NMBqXJnn/T
lFTEfAWW9Pte95B/ubrfohQzc4vgalVPsrSJ3Yq33IvluKjtyYYc3FM1vqHoaKYJzF2ObkuDmPZf
HuXT06/J60j/jNXhvvvf86AYvOI3BiOkEdkOfaNGaQ4qlu5A6mWBzqKLdklDw3Hf6TKuFPQK+I0t
VMExYtVYfnx+T2EJSTJNOERRQe6IDB3Ku5xHbmkFJq7JWxFeyB8HVEw9kpDLj6Wz0k3eVFEmNC/G
acAvx821NkZOcSqO49TGOdR5SC+dCoJ0C4vs6PoJxq/4RT5d4yZp5ZhbrEPAIWPbNxZRyIz+vIia
GpM0gJ5kNy9U1IXgsYz8ZYcf1XQGuge/6sWvqr8j8S77c8Ud+NoyHbBt0qpej1KEsic25duEKtkx
FCnrZcDySgT5qA9lSTY9Nyxfkooy9pxYJ/icZwcqg6JlAlUg2KeAZv1SDCjou9yXotmh22B9XjmK
iGIWkkpjpZ5/NuelWt3lpNX21jg2APXK4An1DlHelYFHEBm+nhf3U9DUe1om/adUgFaaPKajonEa
pbpng5ShRzHgQxVK2IaJgX1MqDAG/oTktc/xoTDboFLeXUSVqKJqQfWvqY49va6qb18ytAHYfAqZ
rtBAY75QJ0sAKWXLFkkukzpJXBv9vEy1cBZcs/0dv7hnQgPgJB8CuPx3XX1oukvYoj4ei4CfDbb3
Nf3knn04jjCyoEigaLgjNgpo/PmJtd/vCMRGo4Xt9op4TT2M7eI1/CmE7tFzMKLrVeCbHprHAA9X
AlmSMFJzGtvUwY6jIAjzlEV5Byl5cztOINxeOYuANEV0mBsvTtKwKOJrvyrUsbovn7f+czFxXprI
KmB2YRcUNT287cUvNN/wV1KPbvGr3ieyzJ1LfIjRnLYA2zsxbPwLLDsVwmAP/lMOrEovcKvSZWcO
h+iFWQZvhDzd7jm+KeCnBMBgsfdq4bHZ+2iZ2FYEXbEJJ+dcr2Xeg2jFJPlHMFWVnU91xuzZO6r1
lm96G142g4x3UidDxNqbbpa978O3mzAt8QMREcHG7KUJkbYghzDf7tEGx8FhK3BLJXvpxcEPJYQg
I5UCLhONrvjA1HChF+TpGN+aTOZic1P9+pytzJNbrKoFE4U5MgOWPJbg3LkA/s2ThvIlaZ+SOzWn
7LdQO1QhMo+6+bAJYeIGY5lPqZNXOMKLUEmjw12Bj3Wk0EJTB7Mh3y2zjwGZuvRbGxepzvqvLVzr
LrNZCi9RQaZe+obbNvetkm/Yc4z+sbvciFPaQ9eeIMOdAcwjcEUu2mvJATXQX04n7+kFrZs/UM8S
wuGwSUiVE3zCpYD8I6NWewnImwg2UgzLU/+VLukF6oHJ8Z7mDfOKan7Q2J+AWccdbK0oLM4Y2pg2
d0sGYw3r/GnIr66TPxbe6dFshZHx5/9yEkyBj1bsPVNWc/XajKwJaDhzmY2QmGmlqx9eDV0479Mf
xqmV48gw7WrRTRTa6JnXcw+NBSiLT+KRBtl0QpNW1afuQvW3F6aXkJkz5oMnTAIB4FfP3qYckGbp
Y9sMnuFcnAHihFtZyxjgci0YTV5lXGcbKAm57C/+Z8UmDDsYiZyoqsIyaeT2XhEdbQ3PrbqmonFO
XantDtwGL/fcvE92t7G61g/x9ELQJcKW92zP0FfBun+t6ga+FA+H+NKYxevZcvhqomFfjd3kQ3Dc
iBlKfUTkuhFOTXYCyejjDBG+KkPii0luuUntRvojSJ22ZD3v1cP8+dR6Fs6Vjs52veICFZf3ulVb
d9Dvgot3/d+tziSHsDjngoxQlAAOKn+FMMyuwKOOnp8OSqVHzLOgBD9JmWeIk8oKPtNJvpizNi9j
Rljw5v2cAw2WwP+rf/q+W4soAKS5tINL1Z/pSZL+bS+kWb1E4oWv4BMsV4xkEBO3rrJzhAFOdREx
b2jj5ObBPUQx1dNwjbKpEHJffy0e+3wFxHNnvqODWOFv3b6Nm6HGcY60moDT1qy8gbcreURYhlX8
y+yucF31DqI5u2E08wNiN28dvo3gsO/HbcCaRGfu0A5NNsPW9pXP5IMUPmcCLhbFYL8UuRq2rmGi
75Hc+L+ha6svdaKWokQAWdQ0ZOnk+DS0AbykgFjHzZ+KbPYUWgu/tEWkuK2TXp1HvEAVf1YPQ9ih
IOr2sDQ7i6id8vZx1CJTDBMPtwNDhUARjxT99CXEFm83bznGN1NfrhA/EzPgjzL46xjpssQiKnnu
aeooBa0Wb2r2w4sdaiGtA2EugolgVxXO038cWsOwOvxNoBoSKVY7XK7QKfJMfwPgtp765XSqY5xg
Faid3bf8t/IHklrmzK8Zjw7fETK6+kMHGDnJc/6rmtDbNBraHwoVxp47gWc+oDDFxsTCBI5/Y423
Eqk1XXnzmsU7kQMhMh8G2hNL6LzaztLraKvqqkZwLWUcotYhQMQfmXHB+j9ZpYQZJYWghr1QPPzG
34PdOvex+rSxjyop39MXEJ31oyAiSYmUlSfOnmhMxTbuNxhs55mpY+aHpc4PI+XES0MgNUFQ2KEL
3+v2dBTVfrxcmRt3V52KwDeqhT/Lwm0p/sEe98X/YFEsOnxi5BQhAxLGVLqGcBDLT2o65uzTlQ57
u150+PXW7SfRiSJO8tFh/ruULmFlePBu7HKxseNvAI4Fi99MDA1/0Ll8qgaWMByJCWU6iA3uSG8x
VgSfasJ3l7XW/+SVwKX7WosH9o3N+i0ICJmruUxQBsWhd/ceQLgdA3hum8683AcxZPeggksAefxW
qZQrobkmq3GFedOoemSMsCZBkzmggYjyVBrz9cvIvFNntolG0FndE5WN2VKdQyz1kVwHeLT2S1E/
nIWOUncMJl29XhXYFd47oe/2pPCloAI5iXH4xyGM2uErcgu0my/H7WpaQ9RMaK7fjYbN8iwhoKW2
gElaYGeWadZWlxTL50vMGtzzqqvVFaReYyPIkFCI6lYRusO1eQlqtCLallqFZ1MZkNLmXNKJVncj
P7Q3cqMtM2ueCR4zMxz1TvHp/A4Xm/1TQSx8Ye97p0pMLPwHuDblVyHf5bDlyWp0SHQG8aJbmE8f
MDG8v9XMXi44jecwir3YZHa2EnZ66nf+9oNriB1bOUtEJYo2l5G/Gjx0ax89StWYVE3+syx7sNYK
TFBx+g38FmHXR1nwP1CkXyLCnXaKK7PJ/Xk002zl4z+O7I/XzlwLpVkXsYMAMuqx7XyGBu1J2Atq
UToPhivuKzhwqM/U/ejajLCcIRM47k+vvRq6q5DO0CChHC7Et+dQ7D6YsuWU/DKEl+aZyUwxj0Sb
PkZr+2pDFdcSDGeOgGJ/4Nz/N1ejzfH1IVy62jXrpNik6yHLvWDD/j1Jl05Hljqx9RmWiV3jWAim
bO0SmA1cHYu+u196xt/0h68qo/UcddQKHL7PjMO43oxsjdWgvFyY+xt/udwXigo8UNweaXr0Z1d3
Fs+94wep0751Z5aHDwIBQKeEg1pLaJtS9R8gM4xpoed9jbYTcC44Rx5PB7RzX05myAwHQlclyUSD
2cNu28sftrc4NA41b8v6gFY6LYSGwqXVnK2/cbMY4Pu7L4xUgexOcHlvdGYIcEG55YImSXMmLwyu
upD5FEXlsjVUiWtfEl+oLUXo2paMOiWNPojrrYRMmSW4ghxrsTc154YUkAPxPDrFxyiUFXarUTxb
adY2XNhz5RZYqhdjzAvYGmd4bs1RLs/+mKK3MRs3FVR6vjJiHoVtiDrMg8c4LybaeVJVJ14w0lM9
XZ5v3qZYZMUaMHa/u2rknV1HQcXXoNheLRNwuRCMDvxVoashXCh4V0GX/zj5wWpOMMUUzZPmr3Zx
GCSRduPOSlb7B2Zy0Rtnq+yZ5srVrGCn5DR/XgYHMsA/yiSca7mGEierQh0I6a77KeHYUWMWbeJa
FqvuMYVOdY5hvwwgpkuQKOUq/iqo99RKD4cBfMaq1G0QCp8DEw4u+3Zave7+4s/v58bs6g8+xOiv
mtMhYSHKtRBKQ/h70Y7Q8bWoeVX+YOrZ8CbDQw2l1i7UvSLyMmwsn2e/RKFxK+vZ6GEm1Kyyv/XC
zQwAJ1X9xgm6Xgy5rgfv1yU8OTw0CZEsPiwpcSs3gk0eb4wgGg64E9hrgpxRpKPoUF8p6aIuUHny
GWRhFXgs+Eqr0C3BHTnEblq4vUsfDPagOZIrhN35nPHDfL0WTUdUd3bPdtww9c4qr6z3v1YSOshp
ulR3tddpj4xWknM81RHFrCAhwE2iF+3RHPHKRsi/oV+svdEvfA50HDxUk7XbnhXXMUGElNCR9TiK
cOMXaV5rydFzFlpsAr6vdTpenLKBw0mgccndWytOLECZ6Ib5ETmXbPyb09jNJHCHonK/QsQ93uau
KIgBNuHMhpz/1DYxfP8/NYC82Q4M2qmVIqOS9hy72uTfK71fL6ZxoxowymLkXGPU3Zo+yXWKvpXS
/Pep/BDgGuafrxcrEh4Cr0/nofJARr37etP4b6KoksaxADEYC9jGFpoK77emb7WEreHXeakGxaXy
WMAde3HebzHFVHZo+g1QuAQjKK0eXRzj1dsZNDiFjIBS1ahXetu839Qnnozb/hZNF3AR9Dj2foWW
N3wZcsXtzinxnMUpI0nCb5IBH9GPzKRB1m2tvcgdM2qHB2b1jvZSC2rLMhPt9mu7yvfhhME7/vFc
BJDqJ2YNUjfn+Gr5sMvXUz7EkiU5l2KbeEy3/EFTCKxRKvP63XKZNJ3fL/3pWQkdZtJmC0JX/fll
yEVTPxrEglHetI+eKIa8DgEQZVxyej/7BefdbJjBfWed1I46TybaoXn1nMBL3296cuYNRHeioIev
mClfvAY/0nqqHaAyuiJtbmJaVZqW+CtQaqx+epsUMwu2SwCDLTBUtb8WbgIdfKsX+++ia6EiqXgs
OCDzA8LH2XeHN5Jq1mp8hraKrd5fJg6rGsno2eAZgq6TIMLEyY8ALF114mKUgLOmxef5vN5zKUqB
sNiC68HkWfX+MTJ5rtviq0oIOcC+0JElZiosSSdbOKJTdgQ5P9D1WZCmZHLg2s6r+Ia3rR7s9II8
6uiHVXtnklDedvq9Y2EjGKgWMcCda+1RyTIuqoKS9oolJevZ1l7Ef9lKr4l7/jUkha1g8J/iAAtp
sEsFmMjOvPPwI0kq/BGAqD+wbIQEJ4iunAvj+muhSk5OU+3Kxji4wWcUFB+pkAJYqNUbCH6dQV+w
YKTGNDb2lt3I75PdydSf4oijGeOLtUkhZXT6Wg3ZUau0efxj/umXumI63dprRjNmdWPYfic1zaam
+9FYEAUG859xkAkcivQaS0f7PWI1SFALCE406SiNSpiLXK7L0hxKzJZVlR/mu9hMtGWIFBws+3LV
40lmWPCA9nG+E/YRtzYuL7Om6JRXPPHEm1uQ7gKp5KVuAPglgs8Nk2Uiq5aFR3PifIKuqZdoDBQk
It2JFePayrL5Cmx89pZ1ca9LfC8OtG8+UO2qhqyB9WdxURJ/y/vX7spI9tgkxL6JDQJX/V8uGR/d
XFpTGngxucFsINbyTjYbuJGDIOKZ6Vn7Atn/nUGGFVmdrjC+os1Qcbawvev9c9YbFjB3Yejyw1wF
0beySs+ruHOu7AteUt3f/aUayGFXjA6oVrfaEpY32eOuJRwbMvTbMHT71i60zCVu/otio6vtZRf7
hThTD4QKQHf/nvZUeZoRUArwDvQLW71Npbl5zmJ7MjYJcpm6w4CN1MmRaKnXeRaOm0922SchdLOZ
QeahYtxWHygpWfJxWir6u6vkIueI9hANu1Y3bISfiCkYb9XkbhFpFpjkRBKDT0o3GLxrJMMcWuqf
HAFyNQ2ssteh35FsWqt4/AOqf4f5sWUAHNCD9DzZtIygfvNLsOxrD+lh+QRf8iqG2HOYUosWF/6n
aRFPgtmTzsA/6KTXuZW9iTEE1d3+dZYJZW/SIfZ7rfrjtNKaaRFidDnb2xeybAaChBkoc3C5S0DD
NdTsiIqUeS2HH1Bkmz1t0qX6sJQXvg00koX27s2lLN5pf1n1Kd+xXnWi0kCBcBAXm8e1M7e32/nO
L5hFneYxQMN+1kFuehNdrkB3Bh0xfb34VH+kbD8Q82jSNJUPLn3rSz7ir5BwokxlJZc+qzbOaIra
KdKW3jBCln3tNMuhoJKUYtVRPfYX38sZ7rLr+gkQcJrku9vsR9MIcqFBkeOkWC+9WGu4wbcvcv4h
EL4Wbnu2ePDyBgwVqK2zDi9nrJjc6vDD60AVa9L2K7oC//L8jD0JsaAEqVrbTWJQ/yElzw8Jd4jZ
6N4OYYm6Y40JQRKXpZdUCjs0IsyyMKf/4BUycOmSER6ZYZodhFLld2eLHWTKtYaYzhaXtyT9UPNc
wctnF1TqD/Vgkt1OX0g576SaPjf6b1Z46kHYEA3wBtMNnpSPbXZewsYM+oDM5AghAZSUABElJ1sG
2UuVA/LtFJ6G5LdtYuGHhzoHSlSb78Lzc+j5EFBjkLY9E52x93bF0LQSyQFIcWEqsYUeCi77EKUY
XOJ4x1uR/wVnnzbiPoBypxBskchK2w/Qeovey78kPJ8DZ2h7B7yJi0jbpBJe/BtsF0ECopuL/AgV
XDN1+TyAolWBrU4cIvbA98h7BgOiyF50WGX5PF3w7VfWXsmjPObhIme+YlHitcR9MZ2Smg1SPGoZ
im4RS7ThZVuiwu3wQvElVe5GPbgxTTYBzg0Kh/SS1j1XaTtOyS0Szw4LXO0NTqUw3roPT8IorlXk
RHRhDH8/s8mI7C1Rz3+F8FDby8QRiVc8rkcQ7trVgoOcL2dOWTnG9gxM06QfpAOxfD55y4DBGadJ
3OqZBrSRR3OoKNAbpe4DkLttYFBLJSRP4NFuF6r5TzIXAPy3rdQQlmeIF2uTg7V3fb1b1aRryt7S
BA0SGP687PHshkYsqJzQCWbQEXZP0X/me3IgJkyzLNdzos4tcI3AEKR4lTMsebvFw2a6ClwEXwzS
qoioHICxGF/IGESn8G93RIF35egR1zyfKaeHSs8+Dw5fTNNlxKv0kuHH+k14IIb0WQLkNuaSsEKx
GAM3gVPrUcWkCHkUBzg40kxmcBfM97pcUY/d2Bng6MW2IovMri0BNtuQCIEDKz3cEcTS+30lbmpj
s8mGe/ajoNXhxORTEpcasuLKOYdXJ3ekqCSo565h2+pR/1OsdZBqrHQb0VLwdee1WvQezUVoJ6tT
vLsYkj4P/RU1RY7Eb5PuUoT7+zNVxct3K9YL07NwP3ui/U4wfba6B1uISIrZ/ObV3zxO+GCfavn+
E5YCS3jZ+774XrFbXOrWYwDLMPRPokbRp3Lsi1NuCXa23lpxOOMbcSkgas5o9zg03VrZe9rg9TGb
kubDhIeFncfayFAKzE9UUQ/8uR3iDCw8bXZ9CmgFgQ6emrTw9SXY8lhnJ71bKiY9u3wCbOy5b37r
7zGEU9KIHxE0VdKk3Gvo7yc25y4Da+sCzMVfKbyiNRtqhlTTgW8R3jEQUpgxPcbGhTcZc7Gy/IB9
2I/KZ/UOgBGFsCQNkXCNeA2ICmI4Bon/EvOcmOcYQJniYz8bt5Jn0qY5WqXdUaJnEmOvOR5Mm6Rv
cs9oUhIaeB0JrK9vgOqTAoAC2zgW4STkRyTIlqIehOxpy1Do738Hz0vzjjTqn52pcJjOfrMjoXuC
dfHr856WkEShFntmCPQaODJI1ZbFVGBrXzWpfrrqlIqctqFmHMaS/NcJi9NPThdENCaVUgi153Zp
V9+M42Q1bHZQkojVwltbFFQf2dHvCRqV3M1V/w87WHRFA93Ncl0WiVr+8HnUfgX69LZVndcXdtSY
zhehfqZ2FcpQ4RqT2tDq9WekVUo9BkYqsqeKeKRMMZqaPhKQqAJkke0tvVzub8+9t2GkZ+iw7Ksx
gRL44pQyM+V6KvuMfr46yEOWCistAi2GewxB1/2xbExQq1KCwSTWRoXOtbuI33YxZ0umaCQ0utSC
17o5lR0/Vi0o4E9e/Rjp+q2KBaAUdN3txpayEPhj1upuADkKvbUygzdmf6cKc9ToeMXMGijmpMMT
mundgFvBCVR/+A5zm8a68LjZIPjKUEXUOKhMi18yI6q9atBftZoAtBtjh2XisNdKFnLGYlgW3NJ8
6N9dn29BuTheOeHuhDOQN119JnMForhfRk4noKvpPWXhzJarPRx5teMJJcfiZ68rzV0sPT08buTu
Vz34YtnxCENeFLmEC/+rN4avXyuthfnJAAzdp6RaxgS1P6aypHNhecrOBm4oSXZVRMU4crl3wUAa
bv+E3aeJ6L3r1pUsbKszdzIZYji/oD/2hN2fMOoj62i1y3iuW2PiMsA+v4rG1Xb+iSHxjbUfHLN2
71srFWODwmfo/yhL94i99mtDY4a/v7uXLGtpwco2sYq4ULPDip+S7ErvhWcYwt7GUmjJEgdQYf1d
gqVAmVLQe/QBco1pfkn9j0A4Qhr0qUoyWOKEg5HLAxFch81XMr7cMJbart5VZa/EWxTeaVpyWnXY
eWMpTgp3o5JWyDfYUOhbdkc3GOhNdesO6a2WBC9DtAohtDGq0YCsvItG8Kmm5ZWspCs4Z7j5NGJo
bki//bqhyIUc2HW40gXLE48tE024SMVYLmE/WOXnbN5zgHO+iZUcoNWipDpXn/3y2Ot3n79/doPN
SgUEz0PW1641Dt5vxfsG2HP11NmMpMs2isTRFYdmxeT6giHPSLp7OJR/GCDe7MEHGFifRRN7u0/D
YAsm0znt6HiEQtOFVg6C6Ls7b+VLqVHZTrXAoI4TOMWTwxgz3YYJ/WkdqV6O+/7jT0y08j0A1+vG
RVC5X6cmW9WzgB+ywnzwzHyJUFkYIcKb/gPj2V5sB5EK6uGgKG5PPbR7yu3Yp7LPr5Dib8XAy2ry
PE1HAaDs3mB29cGMzMT0x+tWJM7DU/qO84aRCn91/vOEqoFxaqA7yfM1s3m5Iim+ogdsr9vIJKlJ
wQ4UW/v1knlWXGJsVp+amYca4kvNVr3ecB+ej6TeBeaZWS+fOcVCdAeby1ee7S9zb84SBR1Ykh6a
lBl97AJ0v2XBhdL2yhPQL+kvwDcoRqOVmtxwOYlbpfpt2iXHRvAJTkW5yYH1Ne/PvikBKS84VSnk
6AVg49FGu/ZhpiNMRaVJxqUwY6Yv4Wn4AZ3XDTe+xchx3HCxVkk52M6UxQL13Lz5a4Da5Tnz+Cpu
q3C1tMtB72X5VJ/cBO5fomumHK+LRu/zpa44NojJsv1EJGUhz0yblb3zJQj9EiITdv+XbcbWlKPZ
caNKkTrLkoxGKBGY7+NEFTgXAz4OHN2wgs1nM8Bj4MxPPJUTAJRavJzagX22Z5ipfwWbqmuQWBfu
z6InzYHfxWzk1XHvnYdeQSzXSV+XH1reaiJtcUbOoufHHq2ULNFS97yC6E53TYtRWrsSRZMMgwbm
gtXlXNVob9GY2Gb7kF+xM84KDLtphu1/qzS/vS2F0gAWHVkanjGN4A/hqMgFA6itjLMeNru17gI1
wDV0wFZrCne1LqTceL1c/BWmppmhzgiGUO2tTLwPjKq3+1FMK7DkmZoBJFbe5bxD6dmR9RVohemK
bGJIIw7Y0Hiv63i9Hxue0Lidt8n5iZ1oygOKGjRTUgyJdMjCEwYHMJi0/6veO2O+Z0bL4Gtwbozk
VugWuZmBMLIjMOlxEcX7Id2zj1UGvefQ3iM2JQNuyx5fkqCfUmFFF7qmqOAyKg3fyxUmMljiHVVy
ykt9sE6WmoP++RnPRtjQn/ztNPWjN/Ya0w2LZbKbcuHmpvBWWReLAm48oZ0A6E1Ql2gWHbURmEgg
CJkJKrRDY2I7tRoskPwEyWUfy1wwbYdZPczI5j1Ggigtd6xBpn1eKQEtP2v1zobjpr+ax1C3enef
vFXibhQWkAx6EJIGx0XwDpGjpxOsNTf7h+LMsgGyd2yDYoc9Hg1zg6dJclNcvruBGSjKLfpUwP93
f0yEbb3tvc6LhgxZRttG45k1DuOQTL4cGm89qbfmg1AgPN43d/xzOWN51ayQqqlAD+2P5qzwtyC4
vXCpgk4YOcsTw813a+utzaaJxyYXmGtZZT1y+O3Q7wt4205Yf+exJ6kBvNfELlcKuTdjpestxxCc
YNqtRUgi/GeY+A2qWbgxge92x04s4CN2T7RzvUeEJcGTJ0F4gGm0zymDHi81t5+HqB7uCipRaEAd
4+t0a2d/+Dr4emCvpswp300nOo588pKOty59TO0FuuAelfAar2yBBXWDpR320gg1jmuH6Hq9D7lg
0/n+7/qIIxomCUEQnA/hODuT2KvK+LWmnjFdyqAPVMIMnfhFnSSJE5cfH32jslaCdBJDQYXsiSoh
D1ZcmwbpRE6S0Wmj0kf/ywPuY4sw1iuGIt1lJ8qn33oOLZ8yH5+3d01wpYBB81icZeG0JQzJGI/q
1WPJ2udqf/HGsR7xXhGflz5auxZVqHrUHdtM1GpKhSVajnfA3yOwx68c0IBLoXVufVlu999qW10O
pPILG/35rswQ7g5Ge71vXpg10QMrVLGfn8TCk5npgg8LV5jqY9cWERAbGRBdGZkTRKC4tcTP6H/8
ZV4qqppBZ9ZYn6xcZ90NaQhb45KXZ3qvVQKuGsvOCRgpos3onQ+hkooO3HESAS75PcUdbd6XvV6n
Z11nyU5/mnnqCB88MU1zpzbLFIR4yDMSUa6DXtS8l+1HVQvlHnpGKmOck/WO8xw1HFF/fo4tvRTr
EIDzN2v34DYib0wnCmjvzCJtztofsyi8MrnO7X0b2xeAJXQB05tHVjjc6tsgWftxjr036JdVXV5o
XKn1+n9KMTfYE2eyzD2bi0tWVwRvi/6LIADVPEJCUY0C8CyWpUWSK/XrY9DXgjn5mROrXNXTafZh
GXe6kdpeYDLfZiCQFxYlFC0e2bpiE5ElL4JKBxOQjwGZF0r7NylEcklj1ajDTTGZUN8PoStNMVzL
5F0Z6kgCQFlJMtd1/zxkcBo5D5Ps8pME9aMTTi7QcyrMv2f9VDODRc0U3h/sD4ZhPrOPfYCbnYJg
VGuHB28KYsF9VlUgTjNqr0fuOCkoKgVL41GfW6SiuOSjtx7Fb/G5+IcgeGgwqW9J7kSjR/6v/8Jg
VLSB525d9UbmgnKWhvsWVLDfPoFKSTl0B2tiARPb8mKwvsmTqkdi0amLKfp8UHSN0Sskxfv2K2J5
Wuo5O/+OgcA0oEg7Y5wmBEr6RWD0DTKtaBHZtzqQALKm22zrbmq6Dinz/TaxTNlykiGqG2VPdR0d
itg44GsLAl4xFxjjmTc0U0GkfroMkJH7H0FwlQCyIlwwRFI4vdpXHK2lBal8w1Na6i8ayLACMl7y
DZT2ERAz3/oqtjaa2Ah13jNBAEufGhwyy0M4E6GoALCz54hsQAjIq0qHx1Bt40nufiiDCFkqt0Or
/7yUbCqS5wFGfIEOLGiFjtGciFH7P4Lnwg8PO6Hg3V/P2t7lML4AcSF4oQAJ6f0lay1CncGfGqaV
+EUqTUSkWc5yHZdFUsr5ACTGUQGYZqGdpRVHvmR8SJLNd8ZrZX7E8o0adbPi5QErVMSR2eWiv0Em
ql81t7NLkZDx5yctR/H8EPNMsDHsAG1f91d4B4yC5X7NQUZ7X0xbG7B6uZovvrDs5ewPVciTuhD7
0E/lN89Cc5FbkOMHgyCPGg7VNd2yAL9yjpwElgUX2IOjAsGWvfYFjm11xz7kYd1HpoTsDc8PraFO
dV+sGsRJ8D5gIrodQQF2FXXSYRmSMIyjbU3VZUG9HXS6SiMFDCj0E1tv3waGfXgsJ7asNFbgmk9W
6nOmEwDrj4neY2xZVRxwTYtMjFhJZI7krwj2rjnSOchc5Pz0aXv6X6sTjzJII5wdaELuLDinbFbG
CygOb4Tq+GxaVmXFztT+Pq4PaLyytTGJVvToaHwVe0zvS1RrjlqpdRsYH1vhGYtnNxsGUxWGlOb9
w57/6UIM2T3/PnoZrJp5wL0UKfgdJBnKFew4bEMGJM4MJRg/7esEu+hbhDpFfMHhdOvS+624ldaS
N5g1P2E4++KA8dLaTlreaOSx1GrTK4uwohkgFnpS/EjHaIIjxbw89cptqmhEVl4Gux3zLopvI9ZG
pAhX448A4LCXZZDIdHqRxWaq5PqLnpmndH/p13vOpk4wSVA00ZGlwV4F4dXygH2Mhxli0RgM+PE7
mVHigyiroXyBIkzkDHolSZzLWWV3obb2ApBjT5EwegnkDDRGwvQbYFL/y8T/mtKYDt2ZF5JBtOoC
/2ZcDwiVZ4E05dt5KMxPONGTqfO0BnQihuLqx80MegxunGyhZivZGj30R8cZvZ5M/zLd2fw5KHP5
7FqQMFWOHXHRTSva52mYfb8lQWMg630yOhVS2bHd6OKYMeGMB8f7R8RXk/iKM5ZN2L+2pa4njg8d
Qs2g7hGkyV0e2xkjwnaZ2Tte2S8Tumk2AQQ3Qgf1aZM896xfvgfdf7fei/PpMJin/6kQfbJyMt7d
48XoW1e19xpifi7NfPOC1M+vGF7KXPnSMMcY86MZ1v/Wdkl0wURwRsbROwCVq1UfHjG8HB/PMmmZ
yn969X4w5kRLUuQPrjzMxxPa+6duYQ2EpeQF5wV8w0SqzJF/i8QLMPEV/97x1rAn1eH7eMfn/TRh
BRbwmpZWGQ4UQBUIStrxPVNwoyIMjfg3jly35dAJmzB75WsVe/oOYmW9jTjcSuNxH6zr0rSTbftk
kx6FWvd2f9nI+TVfT0ThnnG0BypcoJALkmdOUUeDmFWrwCQFnUMyGPGFffEAAqBm7+BC1g3uEwoo
2K2ozTj9eCHip2rMudwtpBitlV8SrRfv9y3y9stgxKvEiCXz3XiAATZUGrhoD7Y/HDUoZUoGqLUr
oZfoMcQTZZ8T9LwHINwLLkgZ1zzfNEYeVc2sQ2ku32FJdsNNmN5KFqFiONJDImTNDbmhtrQuR32W
gX0fRUgTyMhgDk36FT4mjCBvlr4GzyXZ5zmql7MuvkX/SruO4AGznJcoTN1c/VLKNlzGwnlE6PJf
erKCzbeZ9vk84xA0nSVO7Y7Tj8rsshmfumGEQ+sN+UIgs/ttixUAjS8hMJ0ywk0diwE2U+6mHvic
I81Vo23P5yprpCjQbv3atO69iBAaz75xja1HjWOkOkKBN7EXZUjDtrcwK76jbS+T2zDM1QFNAAmb
kbS2y2nUJTFcbmTe924zekDsn+sJk5igTKvuHBJLSME/HMg5iMcJ6pzfmwn0huOudaG1bP05BBKp
QRilCaYvBp4Fhh5CWxktNtI+KW6Ck8N2B98KvmfjwNk+WT9lHm8bef1qkTnu44nkgTb8d+HZWt9U
I1VVVQBcKzjavROPSeKjtgiHZIiRNExNZSy6SHf1+Eoa8k41sqXzVBzhUHz3Gee2ae++pRm3U07U
Z+WaJ4/vUKzxleU9cdqy1zER2jbTKzgbdyyG9kcOdNH+Ht47qreiSToET/DPAcb60Hx20tXAFumQ
BC9auj8leqrKu3ApkiZfvzO1taRf1OOlewhsmi3gdEBFrNwgaANtVdxUT43YG5bKT7LLbpheLi+N
TVLGGM1pqlyhoNQxAanGHz7wJ40H4nmDs98f9pfowQjIRNcARzl2alb60wphfw/54g/3K83ao5He
pQU93xrJ96/zw8j3QKItdgFhJ4QS7J6xEmhj4CGqPf+0x2JciCPFmvTSo0qlIIdR4wssSp1wh0Ti
BAzDLhib10SxXCYAOlv3sav0Mp2GLO6okrDXtkwyankZMTPAnuoPo7U2xuW2YcnFpS3ZwiYnIJ7U
iM84kKXNVva2ztsY7VexuQhzsXmzjcIxQtas8NTC9GRHZIFyaYgplI1drsQFEI/aPMyni9y/TwxA
f58NrDDHoSOGLfTfiBJqXqJ76TxiB71YwOsHnE/7tZ459HqMpzo/TgHWalziL+EohzM9Umo1OxUc
mnpiyOM6I2hfdxUdC2SVJlxb+vcuoyzaNOwpJhvkjXfqufp1XsULToELGd4Bj1weYT1YRLlLDBi7
OrdY4PB3DWdPhRNkQnjiUbXDqibvwcyWjoUq5mOoEbyTJZ5TZ4BVOaBxb/By4M5zphMd1W0vNsBv
TBBMnKfMBPHTlqvdv8gKebiYkkY1C3TlKuDwCB9OCiVlF97q/c3xuWGuM/fsgmZza0KsKkrHXf3n
UTg+7VHvMioBjkkuSKa8Vi/UBiv7mOE8ijuaSzI0lyY13VDJ/kif/gw2fiiFH120cRsNiqtinpqB
1jbeRZnmnOksQ22TIzPMuKAtZdy+aaflFivnB3DSpMhpHxEbuCClr7Z2nWImqSE2DDBxXVo+xDSh
9vY/D5FSA43YMP0CEOW5MudHEoydwPZUvBqrTbAZm5Fw9xtL9ouKmbABf07OIwsgOAiihwpb9Snn
c+POnfc+SPruMI+1eiL1iqtVQriGk8end4nC7ADaSC1GOGNfwvzvzq2C4o900ZIolqXixYKY59FL
ov55hodfm5bO/Vpds9f2E9indJwRcwSBvvGBCZjlU4RIR0IvErt68l9QBFF1DZNi8IKj05GCemK2
JiVpiPzRVRTo6+bvzdjEaCqBwSeP3xs7AoslnlGTPzMcMwXH4kZxmhUfDP1QqRRxf9FXkztJfOvE
RDZXnz7O7dfq/AUncarn1uAarOmCGyKP1UEdpod2D6fsP6CIkWgkRj1rONIcK5S4EVUrBwjeWgRg
J/QC0LXNLhWW4RFxkgowMotPG9y08SM+t6sO+uBWaEb7cxqKpCZ1r/LyZ3db8sq0czWCpLFD4VYr
XXTr28itsds6Cgp5L7MaHfaEFktMZKWdBcOE1Lm5HBkVyU7eoLZnfLL3DSidZDyAclftesTIAvYa
asZC0GgGzXV6UwKy/iQtQARPQxG5uN2a+uxG9bbziTR+aeI1hgtOEJXB0OXv65gnDfeDLXZgM5Y8
5Z5P9lkIlKp60b4TzMHjpT2WZFUvzffyKpAYcu7vR6M83wkZjuoqGPy0QC9Br4OURailPZLwhfqz
BwVCW8z4PNtu/HIRYGGXHJaUJhtPRHW7GcF2R2jSVR/hjw2CaCuEAC42vTaSOy2vKIX8C/XTC1af
d2HCULBf7aInlYtq+wYgilfq3nlr5o5nEaYPYNgVf4zK6Li4K6OWDzK10S8Uo1Xb9z0YYAx+0vX1
Hp2IbWq5UX+myn5j0XNPKz9ktjmE+uWO/7MKxBm20lPw80mBN2dRhekgzeAicZgMXAy0kZ5ULIS+
h3az6ER1lM9K1B0NW2GmrYJQkm/SGUsN0hiiHzXfrTxnJTmVroLqUiwRKYcEdvu5fvs1GkP4dOVP
V0Wr+djd8lghfjW60PaOp69iEfR+bzi8TVP5RrKieq5+dKZFB4R7p05ja2TAOU7VfNNbHyx/RwZ/
Y1gAPATkG4LcAiHsV8usnUw+yIC6C+JLCq4dnSXmUzJEUyap9AsWZnfl/yvwbKbyTWO+6lYHBEsW
4SbE/KhRCOFRfAVyf7YaE8VofQuU3oZVBbxj4F7RUOQZscXrhlg/5Nhh4dFKDDxcKhwR8oTge5xY
j4AuJE8suKnaqy8UaBwux05Tdwz/D6QU/fsm2fPjFW0c2/gSZBVekNXWJGVb4ed2N8x71mfTcM7a
4c/UlrF5/Bya/TfBJ3ofzi9CVm9PhtaFrVIR+ioJ9sgDzbTpPvvBiT7mEv9aPMnbqymXioOjtP08
ZgWFH8wsWXgOegD2IVKK76pAbd1FxrRshzbg7b/3+VezL+k4JPZXUXSBKovjy4A6tW+lYfRQFbtV
GnKst3TpixT7j9PJyMho2pg6W+Le9rnPPv1XhWV5FvgMXvq8f8IrzD9gJipeGVu1eKWHXNPB5Q/C
4bC/ua4yjdfXyp+ov5kTlYLH5/8qRFTlJFpR4X2BCvoOH0IY5rJBJ04QC5kwTWDTqwxRosEkjUgd
7ZwUvzVnOWn6c1PlgCXsu+3iJ1lSzTALELii4jAjSJhgzJPSRwkDfZFoGTnrYkyFFZNkID7fHN6d
afoQPZNqTLsOvcC7HhS6rBzIE1XpWBHTnCKMBSPAmBWU9tYd+v8IL/ap6boNVaxzpmUXi6ExHQqv
xUzMJ2KfXn3Q0RJ9DcZiXtckX3j98mv8G331fo2Q1ZT8j3qj4IcVC+ObpritKDEfNy0T7qQPiOGU
ZMTucOXpwE9HcWyhsOHn3lKoh35bdtKMAEJvP/0D1oT1SpW3sw9TmiYl5JD3ca4O44VhGzkIdlyr
+/AUi1RxvSJarkF8eV+5P0IZt8Yf9785gEOYY/+LGkiDuUfA46UkNTAMBh0nv4JsI9AepCRsiW4w
55cX3cJD8+N3WSiOFYYcM1jbgRBuCIbGtF/bX2xPor0PKolps4E9A/sG5p1sxl8xJSKZuTERwaQc
Y+FY42xMwna7YId2t8bWVfFbeNb7/8pV64DLWgWczYFYelJz+GY41y9EH7raRWsBbYZfqUfNwMoC
+wS6Ld4c3roU+LblY6MjN0ui/h3VrTGdwKk7mi52dPk58/l7eIGAiyWQeFS/X2oAhCN4mIEaKC3y
Z//DNGnfM6Cehzjd4/DB7FYiWpH+cyH3xClU1OgJRB+ArOb+i5gP0zoJs2HLDaSXB8rCNKdwN3+B
0aYjH6VtM1YFF6ABVVMQ6coS68npa1VnkpSVYgoGZnpMjnoq+OczHzo5wDWPvba/Gqe4l0bav/Y9
ebEypc/cjfap8P5v5v0Vm7e3q/nn2asYdLsE3kZUfhDezLD7FOoNu5PByOpJWfoduMZBQ4TOozrL
DRSSDmd13ri8GubZ9NiH16nEj8dEbBHLyFMW3m7ofDQghBafzBIgQRs+fJLtkgd5Exot7eYZONw/
ESzEX3BQonjCEH6RaO13sui8KxXlxgQidgoCCXKwHWclpv+NrmIsJWeTjMbWUBAE9ODB4z+7ydBs
j/gryhqSs0FQ90NzNGSKzFMgB8+36eQWaLneavVG85MY44FeKVfAY13yX1nrXodmlJrf03sOpNYw
Y/GjWhxC8NGwI2gIuryg9aHLdJboHevSlPvEGcrr3/h5u4e8fTz6dJv3JhLsiatyoSKhOaXCmbC8
DQ21WZHtOuU9SQMXVlFmn2I6KPCni+BY8bYeV9Pw4VDWgSntg9ZA7Rczm7an87P98BrzNObJoKig
ByMw6L15JoX57ulYC/qBZVi9ReqY/tItWXnMoZ8PH+6naMhyWhjLGbS9sUXko4vMcVu9KpRluo22
8rMcmWrm1iPpoCo8NFSBqNMDTGfG8fJuF4tPftn97v3dx2S67HIKJP0uKE6y9sEjvoKORUgSVExT
OTEslkah9rkJ5KiHX5M6UK13KFatBjEhyuenaxMGD44cp1hcvq/r3HgMBGtdLkKDlhf0JN4voA9W
IOTaLETHByCG44lKH+nLaU9eDD0rcbDjMsaU7hkNyWNAxLnP9b4e1zNDNSX/eo0d5tOrG1si7K8b
S/NeyGIN7kVEZvP7t6DC1ZS+EzkXZ5U9pC9652+zaAr/6oVvYzpojHSRc2vOQE/3K//IQ69fsK5s
fDEkUT6iRx5pBh4BL5/3X06XhwUcNfdFAEP95pettlfArCGLr9xUNGQ1YKYkRTt9PWcrvktsUPLx
+9kAm9+I16LobXp2azmXetJZMkjAdXqk/iphuFj34IOFfQU3C3oM9TMt6YFHtP/vrenNo7wKwUFg
P5K4kNKb4VF2pa4svCJGvw5nc1uFdq5REyuzLkEX0iGKXnd+c4aPCmem9RD4P+henPqhfq6FzVoR
RufMkMYcsJveBWd3T4zbr/kHe37uBoGLZwUGqbM9RtPjlMTIXVL8WUlK5FX/soS2vc0WcnTAIT2T
AmiN7eUfXxJiTEDAioeKMY2/a2AQX4Xryo6eSlGGkjDDSdXEllBQrrJioQsuTl+VSbryA2FAHdqv
fbt9rZl5ctlt0DAdYQ4AksT+2AIBmJtDwAPUX++9qKaD0F9xazjAla20eYO1q2mxfypJ2NM1mhdf
sRIIANBQAOW/KJT84CYC4ysyO99qdAGXQT6WmpKC+6oTupMSRbK+efeBDVJW3jWIGWWftW2NyQyv
tUnuEy3RD98M+4CAwAFAKZ3EIyOcLVj9dlPWquzI4QikZrtz5FEEw42veg/kd6dNGBKoAe+y6umd
VJdXmja1bpjuTN+E6ma23/Q0HAjOaCHLJa7wnq5IqKClTWq3OJiJgP0dANHk58q6ZS347ZbFGAgU
PSFSM5/4p9ynMp3yFLUJsDfbt95e7PnQbCURcbdUjdN8pvCDATqYtOg9nKOsIMQYAlwGxw1vEgb3
uYFdNqKDRxcC6YPxi01O6Jz287rIRdRjJtD3HDFfqlrMeJ1Xmd2RaQbU+hfpBA20wbq7a4NXb+dM
TsOEHy4WT6yIcIj9J9QcLSe0+SSiFh5eID/iSLURrTGXgXPTwBjngSENCmKSUBvSWUjNBSmYCIxw
X1JLl04RjAdKW5N4VzzmGHA/nkA0pT8XpoBPSGuL58oRA2qIT35TAgNJRNFt+c9idi+rEfNSHq6K
QwhK/RjJ4hC6Nz2gJ0rJMiuQU99CvrQx69mKLPaStKMCmtmHmnL7PYKMRPK1bcJGjdz95fM7S3VM
8VbgnT13jHBu6T05pjzePa5zX29197lRIWLvwoEEmpLURVv9LRabMRiOK2f+T6WhqXmiPlmvKxLi
SXahUc7Tl4g7aQWnncqzT3lLAWWoTM4OFj/xH0YomFWrg23CbZ0C24Mbb/exwvI4CKe3J4+UxlJM
IVZziH7f72hWuMzzvNROQzXLoSm4PCrKlr/xoA54VizadeXapYM9QdbYjMRisuEhEtM16mxoeWz1
WTPirw+kKlLaEpFucqc6+0aZMb+coqbmPPsbWaoYKq5iIJx/tdkBYrK3EDxM7Hx89EE8NlcTLx1r
snxXEjkYe1XkLnkn8hqOf9nsvxe/QTVKSvxo0f46e7YcY4xHFgIafd1peFCupmm2pAxQjYEEaxAr
ceOjC8YPJ8BWDjLo0G0MZRTL9hbuSmUMSpdiS1QbLNlnVaqMeCZrVcg70UrHzFkx71pA3GFGCUuT
h+naqPdfhY+kZgDWOe1i/EoHgZMX3mKh4/f6CAIuaR2HUX+4KZmHpH05S4irx00L4XsuVP431osY
8g+zGrBEDtmLXrSzBXjklfNBZ+Oiusu/ODrulkBlYXEV21+vI5wdJ0+S+Wff+cVZ6IXNsPa2rhRR
ihlq1Qc4dTJDkL11Y0wpD/ClGL67xviwZkB1spFQgAnl1KoSvqBq3VC/a0DFBPHqs9NvQS6oLcrH
3b7oTBm0FvSGMjeHnEl4lAIP9BlkLYcSGs15v3u0D2OU2oaYz/HxXhP3xiRBX4wGZRkuAT84A5dq
wXJqjF77OjM10ZkJbG+ZgY8L9slMF08rHA+uA0DuV6Hicpu8gepFEDR+7URO+jryppf123+dYoSz
DC8I/XYLnK+Lc9Kg9VhcmpkfRgtFwcC3xGDpb+6kqhLKORfqclHyaxKr5sdPGstiJ8gk6W0o36Ft
eEoZ/4chwdRJI/XDoLM3oHsAJ0AV/jPuicbJWIBS45E4ifcKGFG1CynWAESAWhYnpJX5Vchsymv1
GNnTibWlow2hOA4E/tb+DTAGrTYmdCYWHvXW2vEl2GAMKoFz4lP/KsY8i/xSHRNvnPaEpNgO4YX8
dO7xPaahzJOnmv5D5ogVNbZHGvD5KvrXGkxZyYvTeQTU7h3PSNXxgsbdH/QLZQRZVa/ZmNoFIvpe
+KJMCFfBDxi8zxlWHIihwCa9rs5H9i/LBNAg+fc44TRFJQkB5WjavqpFBDKQHmcMZzO3ae7XArXl
CnWKfDQIt6HBYBgI/l0WXkqL83HVEbeNZmhsKFAfcWOChqRSE0XkpYpD97wxCeRsRYyD5LzISuvS
46DrE1ppjw6KkJPinsK9sbUkdiP1zpd+EKY2D1d1/XnQcXltnLFSSeFTUWpP3ZQE/N0QTvd7KGjd
bzgD+oNjr8Vgh6pIPU2r1eEnzrp6YEdx3s+VK3ppk0yd1GnY9jD2NHhfuQGHtBu3aPbOTWUtEXNU
F5sO6sV4Qo3B2SS90mKriraRB5+ActWKReIt7R4wkc8cNJoLtxPWr/ul9UY+qOuNSI1gHlcr9KWk
fIGoZD02TPanP29wxlFOczVEbaZuXvvmzQPHO538aj6gOjF/ETSCm+3oauGMd4iGmqOIZveUBVn6
g8n9K9H9G8jQ07IB7sWDJHdFlutoCSb+kvj/IbmSgYHbLppBtmEBncchTFZNJ/XN3tvAFGrZTBsE
hF+NzzL16KU1Xx7sWzbERrXwRpIYIbBGM1W0ykryJ9JNPQM3QUZPi3PceLRQIGeVXk5M1SQ+UNNr
cgM431cLYCMe0r5cRj0ghPVT8hw874r1hD4/baXyGI8zTqEpByxfAr4OcpJrPLKlw7KHUcwTYVtL
aIs6M288mfAGV7dJGDms3Ntzqs74QTbJ+3iRRWxh15z1x130A/ZSfwGqpbgjdd8kNOfceGm6EeBB
/+l1NLOGr11nMLJN/X4R3c0CczkGmNKUih00ZxMS6Km5YGBFyForsDXn8bRBBjKKd7n36o0VXHDT
RQl2b+x/Znzhh5BldGKdzk/6SArQ66aUTFjZEcML+MwadL00Se8bQHtDCN84OOrvn1DySI0vfent
1Hb3Z2a4loF+2arCl8E6IcuoM4boemGA2F2OVfGkj/07aLl5PvyfMwrJrbnF/npab6UYcJ9HMerp
fh56IDx2aEmfutsRmp6+IxSl/gGb09bHifSq45PEkfbN+ipLnkXAFy+hxcPzuCuYG0/TWUIpplFc
j0y6jalaZYg1bam4L6G2RncakAa0JaoEBTrO8MWBRmOyI6r9IK7vP6QwKKLzBMLZGEnj6hFc2oI1
I7OIh6OtNc6iW8XsdfOEFCqQvPFo8JJ7Be2RmZh7u6QiKvVq3pmCEYGgXpdzjQhNFy0Pn5+MZst1
jJ1fYA2POzH8d1YOvueITgq/jh9CNt8vNjRKVsyUgCmLJJ0/aIAfNUi+NeFhJF0B8NtKvuVJYMmg
pha4+Tyilok+J5pibD04l3+Aec0HTO5v/HOr7asLSOl+/PM9Md8WBcBASvq2O4rwP/Es4ighScfz
a7LQ/8oSfUs9zFnBgZnVdhO/KtVWstVqq3eV6aC8WUrcMv7ejuf1xd+eecl6t28auMxWndC6hNsH
XOlhxEXSQoYILXHRPnhjeZdFlZyLhWae166FMxzhGDk73/UdtXOvBo53GEPNbs7dDPh+w7wUXBDd
iesnVTMMm3CphspJHvYBu7qz6jPGPqybKAK9dIE8b+wtx1TupZpzxlZa6kQsc2iM0CxHQAqfhTwA
vbuvbfENCj+d1Fq229xUtMlh8GTImleoCjYHuZucKyNDmExJGTWlt6UKTTz7BREB7hOXLnPXJNM8
RK51VVQdif2wvMLgBnFIQQOWbmvG/1zXkmxxJrf2QCp5J7RBAqxpEw9FkV14aK0vIxw09WbejzW9
FAEfct2DZU6OCo2wpy22mC4f04PJDsA8OAJOWEDkGNzCY39ZIL2qA45O7A26u/OIrzwOeW3iYBU5
GiaNHEkyuMz0032MQ6wA0LVQvqj4qtksj0Bsi9Mhp5bfjvYwfH1HZwS3cpyaw1Jtkye0QSrrc3Xf
bKLiqF1NjVQgnCpRwD0JHsPgUz/jMX0KG1MsWla8tvcfwT2//hNyPxycB4+BY0qhxQv0dFpjpiY3
4n1ALCyxyhpJDoNjcT19STYyOQbxTtsV/o362dU2qKKvqwNCzd+xNrTkVGdMRtMmK3DuAOgdhvEE
gipFaXe44WoXErVe3K/ggXa34OuGpnQN48t/XSJ7L89ZwOy3PF0WjOWGomVhwp7ALdvk9UEp4wsN
l9txTEzIWuXsrQgcqEM5r/HA0qdS8I/eklSuL9DexYTAIrWDl4zgGmElFz/CdGcqr1e/QXizrY6b
J0Hal/6G5WJ/HPrOWyYb4Ntl5jmuvyAU1lyf5iI9b2896JcanRuJn4QH2lvPadGI3mg5RtbEsOEW
/uvEbeEAxPFrUjTOIUDrgKlknqBk44pv2hADaLEGFKy1KTwxlXxRDiH+Hcdol1W3hVZjxCA0F1v4
i4M/S48zhj7rrG2yKll8VXYg+ZC9QkFXQSrlm2yb0oOltZJmYh5U8AUdfRkIPcnAWydrpGZw/8ea
voMYeaVanDsWPZj8GmfXgOhXFFKDL2LBl2AqcR+QR+LjVUrXgQ+B+/edCtzqRfTgQ/i/N60KqcmF
Y3ode16hJdmYYCdA8Doip+NXohuPe4U9iUO7V9/cQaXhDdlc8e3LbbqUuXZv+dK7686Ogz2pvzjA
jT1PIi82B1qtqaBAQzgZT4zCNY01zm7EOgEnvNeK2Nmj4nv9P9m8GBJopMUD+HY8EQPINgOEkaR9
X7Soc8UDcGm8BPs8yCi6/g7I9uv15Gq4V7hRGLgXsDGlfA+oqInzi3b49c+VelQFR2V02+Z4Q1/v
rCxvS+S4rACjMjpmeOms+CkksU71y05mFDy8GtOYAzvnyxu1inEipxpPhf7gIn8D9nOHaVTSgzXq
Rzp2K8P18eyAKjCryfdYKs11xrZjLtrws++bD2895heD4lMY+z8BS1j9f/NPFbvKHnvlWcsHCb7y
/xpZvQ98/KUdqwa9YJUxNT+Vv+fy7u99RQyPYtnpdwtpxYgNRvOrP9KRX34cZTtkhW7F1WBlfGXm
5jS0DzqnpGTcACKciKckj9o7v04aXgOw6L6gzx5CP7HP9GaThkrpFuqHOyxBAOUMziWSF2k/0QzY
ch5ROBReLk1nfmT++zakSH5OEedm0GBGhuh91ZQnLvXEg0amH1aZcYCdKupuMbQBIInxXRyQtT9F
JulTfgZSi7+WPeBCR5du4Ervc1kQz7A6s5c+NP35Hzj4jOM7Ja+KB+zXg1fGrit/fhnZPTMjtDsM
A4XIJVaeLjaDIoPWrdiuKreF9vpGndUj7B/ZctLPmU9YJ5giEnCawKQrm8g6L9J3gimkXVjQmIcB
amES7MNAsmM0cBDjRqXCY34tgho+0RvYwSW8bYEIetR8t7XvYnSKpBar+N2usvPE3EIyHNckBTyO
yAt9IAaXqjQsiE8zutGeK+lfryB9S6XgIl3k0Ie/4bTVgyCWX5DeRPeyl4giQqsESkxw5K6xmDlr
ICDab24u/Rd/9AznW/dKZIW9LsMMOdddMdHdKTigPf2VT6zZZ6vSta/fmRvPz4/4RMA39haHZRlS
EQx/bG4ykwpRUmXhEccqKcQi/g13f+7ROCN8FswtVW0sboUCpBSYdSbPGdO/8XFElvErZP/pkWcC
3aiRYtION+1FJNCaDKkceiVlAIZJ9adiEb+Mqkh6aQkkuJpfeEicfV7Zs4ePb3I+S2wCvfH+LFuS
QRNPmy/MAEIgZxQXKjId6cwIQhfL8vJ1zP7JKSqWqC4aiVIe2vbHJX7QK1DYAUt84cTgQx0FbAF+
O4vgAyc1qtLdQYRlJeshP9P79EtQjNNr3o7Qzudv1e8Id4WNGvMlTtBMZpzTTtYlEw78Sh+RXOGX
YbAcfXjZyBgzM2r7Ei+4oYmjkL5Zdspbk7YIWT5ArcgwSf34D4s6+a9zsLoCuH3VOBFerXmuTPn8
yQKnIGG9wPToto210e927BquXKH13c+Y+cMq6uyxFjXqUvwAIlH21TTQ/ZkiR3+FkNAhzvaIbm/D
gv+Dp31RIMWNVvmnjCSwdJbO9ANGRyyBhOisXaBeAbEsLUfbUaK0yyqDqeXfB0tk34XO3OPoXWJy
fZ/dvYD8Tg3Y2XbPMzAyyh4+4y4a4dn59WMBtvqhTFEF1TOo5mq5CvA/TjiHdupfspKEW9mDU5+l
9g9aS8vLsdrcYA82RO2dtZ+jsWqxItHHEso6YttXuSrWXC0vWjfif8n8U0gtjcOgR1NG53Kl3WRm
kXsuNPhY+FIBVWtlHMuxTR5lT35Pvl+RhV8t2ui/lR44pYTxKUp36FSq9VXBFtulZzgwbCLo+AQj
m2e/s2JjiVo/RqEokMFJdfFZJMUNqXokQvknJrQu9tqO/GF0QXE73uJlFvvG9I/1zPH4M6iK1RZO
FlAFGhNAmDRoeUrPWxEcgLpg6f9hqLbW1inLdWdamK7Pt4a+Ap0Ass15oT3FrDvYBV3ob+KiqRuC
kejOlsUb41RTfOdsq3oieNygm6Tv7g1jkQS2USzI5wnmk0N1SiURKrXvMZXi6QQ42MxfrKXggWPk
Q4EHXRttRl9k/Iladwou/c/14YvgDV6Jv76pUoh5TOrHFwHiGMe1X7hDWgRLWjtyKbbof7npr9Sc
DIt1bLD+hbVmKIsfnsPl47s6DvbdhdTw75bCS10euIf0CL2XKnkwwKuKjjNBrixq4DInpQxTzZ1k
Q0qNcd9gF0VtFFDybLXC6ku80S2zCqVT+Kil/NVU34dGyzAH0+AqA1sZOB4LjJPY6sNWS4PAh53Z
9Xq/kZqxJQEAb79AzfCACJeCrp52bHdinhIQA4LUye35z06HFgz1cR15WSjyANStuF6HFdgt1CL+
7OHdCxvyvqcA4vp4jFr2oHbiSpdmGqmkkyQKhQN7/5N4hYB2Z9RCDB5IZ7LHeeBDEPzy7S1GLFU4
uCjnk/ZwveIeSRQvmGGxbNM5b26Nz4eqmBgLgFWwijGMJwRspfmJO1MutlBMkxfAzvoR9ynxuwS8
aqtaLbmTlQ+EfDfsWKZJ75OIt88fcnqAPSq42DLs8VnakUOUtgoCmOaEjqfM+obeSbcqFB/ELnw5
GBh0PQBDQkEXfGxX82P/QeuG25ibpo/e7tF3woHhiCnKkgUlfuitYJVh9W8fUS5Bj5IhDVDnDszh
cC9Q2Y16pxpMkgLjzqdUsXaFEHHS2zWAdbxAjD/4RnWtm3l3KvJCdthKGb43kblLWWGdx93yG9W8
zm1qe/IufgVaXKis0IZDU5qL3LGH+80SlyONfKn0wq+GMibovC1aw8iaxd1lQ8jfpkZ6TSrt6JEk
fMJcGSX2SXtHazqGaaDj0aHxzVwbV0Sj7DgP9Jr3bm55IyjKE3b/8WAuGOHwubaVvpsioH8yhW8k
wMLWrlCNgi7QqbqA+ZtRnIpX43RgWoUWLwx/ShNFTCOucX5pG9mxDQ8D1qslauPLXyYDHJQ3ujcG
Ie4QfeG982GN54G7ceVHuHdLgRaZOrNvfG+HN0/VSK/6FR1C1bFSsrRzc4WFJrCHw1BvY7ygouDY
XHHprHP+gA8W0CUT5MsXRF7FgiJIkYwv8HaWxn9yY86jxOw05F2eiEpjwB1KW9Jla3IOCDuM0Uj+
Abhk79gVvYkezyOHZjsO6TpjV5IV+wk3aJFKFODKwXkRpv2JppJkhy39zh6fmmRePVL2iwuuzrVK
ZTFla0Ba7jxUsSJJ4pH7p6w9jd1IUttm1Di+SXiesNc6KrJw70SXgZJnPB8id3Ih7rXhoyfyZJHi
sYnZmZMkEU/e7iTBfljkRD1uAOYWXfM530IbHQXnzYGQGMHV3ZwVhKVyMxHhav0oW3q1hCIFDGb5
im/YbgJUCbiPzq3+agig/Gckh3UBD9gcptISAq2qjgskyFARfiNMI6owuqF1dip6y1hSDVPjiDC2
wmJKGzA6dMgMcHNzTG0fAcSY3pSATS1yc4oYTybzZTWsWU9ffydwgbXitiIyEJr0NaKD9gmH2PsS
RqKSbalG5QoErIaB3tYGBab/60dAgBRshOs4/guO7YOcfzFtE6ynLmV3Ld0bvwZMaGFbsodjJ4A1
1rjz7g+2gCYcW5rVK+9j8GUZNvuQwT3cAA2Qtf3TO0uOPRIM+q5k7yhwH9zMSwZX1E1rG86MGW8P
ab/n96BMRvq4xj1zRItk+848tqYyxk4o7pws1gfcTzGq+dt5ZifZGaQEsUsqRIzsd+65KvMJ16vF
HHNJpZwLoXDN7YwfBIzeH5xjFnW+UNC+CFaQc3dl4apcajG3WiXDk292OkLLMqTxKkSHuJM4UhBt
u0vDvbQUIkXWcKjG86b4RfdXkf/sTdCQMdQJONkPofVfpFgR0bToEbMRiTqafBrD5XcbfD0klf9n
hZbVvGhl3kaEoZoh9RXj70oqZZew0D++6jJ/xX/wYVe+0gvcaaBSSMp3m5zlRxCaxAvdJxzkStir
8KFOv9096mpQDQqJMVzSU67O+I73Q/wt7+5nvGLbI54e+kz/ZDvpT2p0vj23w1PrdW8WwyiaWpXl
Inp0htbSds2zju1eDg30znenPwndfU5qfoxa8TkSwQbsbf4n0fuBsZeaWpSlXmCrh7zB2kfuTgsT
6D8sCVVw2zMpkwkjHLaeELXtGjVR9L/X8GSYr5O3++Fg7EXxY6/GbXbIFIvU3pKDDF6zNvGDJVXr
/S3+8UQ6Voh2Y/2V64CmybkMrqUM3oIbyf4eIovLHvXmT69Plz/VjbIWcZoFbZuFuHPsObaNZsU3
gZNNIfz9LHVqQVAU2vj3bS+UfP7aSsKK++CLp96K1LKlArtY0jRo74lJHJUUR/d394IdDRsjpLre
1mBqvGhpOtmLvMURRiT3qVcTdQScsTTA/+pgb1RUFNR3S6yYp8gGl1OzD8fT+6J8XiQotK51OVE7
Z5eJCoFMtU0rKz0pAGxCAm+ZJVcMamCdGi/VttBswrWI7Jf3mPr3kc49Z/aXB+P60InKke/XMg6S
RM6FxA+zsbPdM9Zhm5FHHsWp7Y+FD6SVXsAxU0NVan58LGGj9eFb4jBt4HVk9wzEZaalnAbuVepS
2Q2rLcRptr8rkQolIf4bo+YeNo/68rYu1G1MAKyAemuS6ShmFFZNfn+mv6LVQ4xNgnz+hBKiScjI
PTe/rKysur/R0q3RBqL636BmMfOXSEANIonP0CFTqpX1C+d5+ZLwECS+Crq9MLomJzfZOlFmDoOt
LcLEB3M2kwvmesmUSCdkG2jcTY5w3JHjy/uloXjKeU2cgBWE7oYzxthp/+IZJ7OOOK21TcZmhWdP
ZC/W54uDXoBL6UpryONd1HEYnjdfUOV1rl18WnzZmje8nrqGkldLvR91vylfFtnA0UrtB70q2w1t
ZMrBZDOI47VAOLr/DtZEH5ENwenZSc9dL31XueQ6kirahf3Yp9c65xBRoncsQ/HPC4WU6NN7KRNn
VQvwT1gruE2c4qJCMOu4EuGMBZDnOJ7vWi/bco07LEDXBTic91MwAmtY36kc5EKibIbpjelwJhjM
SNyrRnalbt7flx2xxIkHfG5AljcEi4ce9GVOiMffH6LfXWwKF6NNLcnqQi1UJwylz+AuJvK60/7r
aYReU5b52Oqkld04AwWPZCR4sXM3fi+JxUwOJCsGwdkZha15kA3LwPbnt7jmD7c86z3tuD4vYBQR
x7Wd9QCJMCMnklytIi+qmyVCgY8beGdPHGxthQHkbjusHaSKIYxDbClTAK7wXFviQ80zyqOfRFNl
saS47g/nIOOCOknb1i/PVr5DpXb2psIMsL6TJRcFgiEgr2PxS9msHZHLk/U4MXN60Auc1Ld4euak
PMsKE0BU3TDamoJVXK9Sm4z/7szqXeH2wZw2ZF8CFI9J8dNniG1zvq9eD2Xnm7k//WMu4tsJNt9c
bGQOgpBtnPPlCBgVCPpr9jRzB7QydPoHQZ7e7/qins8YDM12YnGfsEnm2KllUEwZ3Ej1NYAHZUeY
VpCAJovz2OfuidDo/oPONhD6S7qjWyZ+XdBuBHzkjCf/6eWrASE0q9JOjFrbhkgYshint2bA15ml
oqMiswYe6ICiG1AcB3h3dH2mhzFePLkl6a+HHD2met/oUZzb6xht09NPXVL3qejKkf7Y5CshLcZb
G+14MW77tZ6MGV1jBlULPeJnJk9QAAylGaMMkrkr4iTQH9pGDL7s3KEqYAVCwfIc2xTj4gRFbUMn
bZTQ32EJSOvBl2/21VCvUUWzmXynQk45AL0fEgw2JC3B1i6uwtQEWP0sp50Vssy3ohA0FYT02rxW
YMyPlAYPEQ34ScmRhN8IVMiI2NrrfeMu0d4Dx/0Tbk477LWjrb8YFUjgGVZ4/+XBFySEoUi7oR+5
uIGQW6AEHHDZajErdG49ZzxuD3CdK3KSx7ZFKLAB6UUlVKrkxzpfAs9T4EK/8pEFGcuRZPSXkBys
i731OJiVShUBepzWdVsoub5+SinsVG+HMmZ6du6y+b+aSNtEGY3o5PfEbAsdDXk0WGxkAgANkjCQ
orUlsOWsnBPqfkwpB1YrdSkYkroFryYEJT2mGUxEO6gcLmRYrJaKGzvPiXLdcVuVVPpEshvw0h5N
eZA18aVBkeGg572xbWETFUCH+w1lPYGnOcqsZaRXIQonEaF3j+S32dAueSBL7oBvLcqHrmdN3/ZF
p3VA3mitGDch95gkLZu19LAagIdQYD69YkSFQH6g6NZCMZsO74vNT6EJl/pYIXx0UZED3xwhY6Ma
auNcJWGvsnQeCwJS+xNbQ2Ffk6M1vvM4b4+YIt6MNm1Wc+rN9wMhb9TGziJYZXBrx1yRddmOCl34
/z+wKXnGD40S5wCmHpHi8UVInhi88MJcPULAP9+0yyYGcynW+K+oyzZjNH8Y9NHMlpVbRe+RVOhL
RPtLoW01YqBLreRF1Uw2qg8wOGqlpfjFGxI7yusoBfe4lxN+BSrR0VAjJoi7lS23UvZBAZJ4Sp1p
mZtuUHk1pXG5wo21FwFOwl/4tzcyXdC/XKQVN7jGn6wj5Hw+15DrMehYFn6Drz8vm9ALUTgPkRGE
fPbF+Q/KLcG7kLw0Z7WehmA3zz6ucu0XUMauHx65oD7fUzZyMInSk9WCraC7wPSueUrAPcVKrcLn
VkhsHAumyGlfQV1nlDWASoMIefNmlGm94ryCXxqaylS91aipxv0qUqBzQdYE5lPxOKkUk6D48xr1
zQtUXwzpSoHtQsQkG7zWgy/NuYmxVmyL8h9Li8rEL/pTV/zxLFWp4vDsOMQ5jdf1wtycCCUurJdQ
OZfo1JEAfCol6qPRxoqJ1sT9f085PgLHWLWR7Sl3kv4bGGHJci+DTUPpAWsStyWM9/2OykTKNn+6
C3dGl/RbgfJR7jT53+6JsNEac53G4VxHTHHQcmjQUMbwbsp/DNLlYbXn6dbprd6kXn7zJE2zyjW9
vUyL16qufUWD2iAGnHzJMY+ahJgMVpne3cSs7LvNU0XrL3KngQtep9UPCnGmfo7KR4KpWtNqVAeI
O5FlKSGgHYDYWVBkVF4ZGWpYp8g3zZbZsC4mHnRo+pqwXauZd7VYJXJggkqV96k42ab6tEzXgw4s
O+Vvmxfa6dneow5SNw+cY2PZUsfBS8qe8kPc6U1f0CmMOk2rooJ7SzivYEDnuz/cOVm9RO14VS2K
cqKpmj8zRJISZdKjwWFXQGHW8CfYG53MZ4CXPLT52xklF13HDwwXO209lF8onMh5TKUVrX55k8S6
lDcxkmX1HIgqQi/6S0yU7NrEobr16Y1gk00H8RMCK52ghzMWw8m6MC3x9Urqb/NhmXomx5N+OhhF
VkV74g2go1R/jeuohcEZ8W0nPvKNM+icFhexCnECZg87AaHwYpB5m3OEBH8mk4KTC9sOHeNZbUKL
MzJ6Yj4L3fXrlpknMAk6Sau6wCVzeE705kb1f38wIBMNx8cA29QrfiGSROCwzXepxUL4h2dueVWX
65WoZxGleToFrXxFFGMlfA5IRlZYNZWfiQsuEbJMZzKRIkcxvtVz1zN8DvkCfJs2hGiYBOdhFzMO
8f5XBV9BVXbhANrItTN6AKXZw3v9vd2WjRKSDrTMyFT/7YSz3RfxDtLrVFrsH97blEutK8SZ+Bzn
hNcaY/qdiVzYW86f4b+GXzG/64psEvyP9ge38vk7aHJUCEWctSYDX/8ZL/bfnYmVVFET3kKVZOMC
DiwWaXNSG89eA7T4OoQhKBdrr/faoQoFEVN4mivJCGeXWzUwfTuvEvfhWecNOk9bpyO+ghTDA5+h
h71Hggr+E3Bi8sKhN+6XcNulsais5rafBbwLVZFXz+3g3P2TuZzDWTcmV7sUL4fJoiJd8R/8Tn0K
XRs11mRVncxjRY9I5gwvHj6gqr6bjrUJFnraGVouXyZ4xHlsqI14SkLO0KOjUQvFhEHNW277y8r1
6BW5uVzn5eyFWhawpsuykIOBuz/43niVLOOmphZS7a4ajTP/glc9uqnOzSh0hmEcMGEVY2du1t3V
ZqZuQja7ISFX3/K7WTykULNAq9ko1EdBHYObn/4Hi53bp8fnEv39HN9Dq7eMhlFurWNvsVuEtB88
lPikYONbd5ZVt7+eLnZH8Gt+EVif3TrL7fmD/mRSDn2tzvHfXFQl4JrHAKZ2xIkdALrbyE8VYKnY
RJmotmpNqSGG/n99/3rHu8k03nZxMRFBa+TePkCq8XkMpmtP58d99PMpgM/KsMI2oXU2HKFcq3NY
Kc0pkE1UUgCkXIvZ4ArWURq8BBWzMlqTNULir9FkskcloiIdWgkePkxBWKU5Kid+gs8U4zOG22yg
TfucSOwaUI3tJXMw4UNxCXWHma0VVZilCE8W9g1OM0avd7eUiCyDOE7JKsUs301HiJRcqmrDCF+M
IN4Lb+u3uKeQrQ+9Zl3RA9q822FHRypq54Nsr8zw8YcixwKgMK89Sj7ZAx9OTcjy5G1Xjl6CWNv+
C4qJgH5MESgYiN7eLfCjhgV4kHyLVH5qJEweCgYLIhX0u5npDLS7V7BOa1KqSxmnVy910rdLOUQ1
sTcDUcb0FQ+g7U5lduRmZ7501pIr3rhMN4DGod0PUxoMINKirSgnyBpZKz5xcoS9ZLsj438oyxfq
Nb8rdSOqFOzfYQhU1mLcpbPhIAoT/0EexYJS0XbmCBIhMP/ZwtO5Bx9ktVSU3ksniPV8poLnIhnQ
CMD2KlCdtdsTSCzrOz+4OU/scXehYqKbUNAxHoAJaoaBv1b0H0erTav5xqJGb0gowVD7pVYsSF1t
xTzGN7i3bfVK8oAJeoOLEOXZVBvAqtsYdl0Is5Av4czzZwgc7m2Y8Di/ql6De53OipseA0E1GbbI
pUuF5FLbfWH9TlWouoDObHlMAqMJJXiHrG+DUH+iMibXB3Az14KceycMKaN3UeURI1maGgjoa6gX
GAN0ToIzfXBguffEMIZK4bT9Bfshzxpt8IdYfau3BNzUbyeXtPpuXHtyOyIGObUp4o8rFibAWEHI
AqjW67GDesiRA9jTfL0n/s9ShDciM3eokxWaiAPKtymVYcR5HXLl76VIOOYgWMjMY3cc9TNeYean
poOP7+C8uvWq8M99zr5UVwGdFmCIYKwT9Jp35M6WizQkp5cyjj/SOlzFJw9Yzphxnd2C9QLzFirZ
IfYpjodXgjHHdH6DvPG68qCWMaVnQHiHDciseiH9kcMM+b1TuYFZW2K/9mJ+Sr68Sm905JdSq7LU
6sk4y2L4ZOyOls5iR0Jz2I6owh28ICnpmBvcxo311ARIyAQQ/IJT0LZXcOqz+LQ9wUWBCS9OM7A3
SgqJZn0fNTow/2tvFmkYGqIjLSEuVYhvWE5ZbdhWWRhKYgVqly5uli5g6uzu287eqBRnVcQZVTRQ
pba232dXnEk2pfBqUnz/2HgEwtqBxsfrLetiqqVdDwEh58nYJFb/DHWyh2y+AJL+dWd0Au9TXOfB
H3NxPBCVUXxytlsiRDIW4oj1tH6NdjnSxfQsJThtlU9a7zHKk/fMpNhn9w4M2EU2oRXGNOzXD9CK
Qxx+SBlyXZCYofNeJ9b8L1/KifODz/LcYTz5ngw5VyR/5JVgU94/wDLcoEO7Ege9GFL2afX9PUeP
eV7EvO6xRb5wEfSqrK8ZE/QYGV+I0yPb+0CH11Z7Jwj0vHdowterxRKLzXHlTYPDbBJhAxKIqpVQ
pHBtnujMQaBlapXfNBi6qS2G+sGzBFSxkfIdzK3ZSun5Hyni6QWDvU4Y2FkYCJr9zmNCTrexndVL
0pF2WnHaOGxpEvywU8h6T57xut84CVT/CjhsmCIUTE6sHEg1YQDoPIsmtjgPXrMZilEdYAB/CX+p
+pXXNjOHEMCmS3XKmWrW6DVMaO+4ZSy9ipJtNVnK78ksGVmkM45f+yvNqWDZroHlUr6r9ZGGjJnb
C1mhQYDGai7OLCdD2kLi2E9Ydw6U1xCxqmnXL2kM3nm6YqQJrw7GsiKsdQ89zBDugsqcwODXN5P9
OVlbrxtrp5UrIUr4yjPAhQpto8QKhUqv4zO14Qh1R+xj5+aSux9YyeXOppLcmn/L3fj8m/miTv/h
c8xswXCaSuKLCzShoDnkpH4v7VQmhz1xMQu9vc61IXNxZndiWeXfcidKIUjCb4SlIEvA8OLSchqj
LGFi5Is8I4IdJgmN4Iegx/CtBjStCOfWnc4RXInwq7WGaFeJJ5G+/NokOdMy8fgNLjXitCMbt018
vlOQRYLaQbyv2sL9VgOGjbakTGwo1/UOKRmVJtBGm3J5ZhuHptf9V2gochiwHbK5Qa5QbTlajxs4
cRAKOHEsTqRpiB4dN3hkl74eZr+kGRJL02yGs3xXDWj9I99xLC2328AwNM+P/4ijtMsNunOq+ulo
LEg+5Gukoc1Eg005grF67WFF9OdNebVhfZZnjzuPLGyiEw/Ko1G16XCBOqtHbIda3AdjLhXYQ+ie
Ovt8JqG59dhM6ZfHOvG/RRawGbjfpN417DrGo/e/387fRz3XNvGVebU3QLTNkVdvbXzzYVaUFicu
cOmKkrZGYu+WuPoAfUvydG+m7SLwZd7joNZJ/W7SBsAYqfAkxrPLeKKZYCL2FKUCBlHEHCBSCUzt
/PXJC4QcdWs7O/JStZMj6DYFhJA57VlpobFxfU7LpbQtqZzVDzsMN5liXqq32QgPTUFxK+2Izmqv
rYO2OojINfuUmIXXYeb6HY0EQooNe5KGk9FZ+gUY6bm6VeNCmvRo2iZFEQzml93EIGzUiXaA0poN
fJ787N+1+oJpmm7yE1FZQse6/G1SxgR59fT9ots9FGTN+iS9Vid40Clcd/D5A/s0ncLtREXr/GWl
vqh36jxwSMGjjUfD7op5Cef4h/JHKxLlQGgVU0FBDBcLY3qXueqxQZWSso+tfShWeV1ibv8xn24q
pzlZrE8U9+fHrKFvC35Qfre+bkneJ+8dKjSLmwyEupqrInIHT+SPZWkXewbxctXpWuZN4qUwaZdI
gSr7XtyVqANaFAVzvBqF6nrwd5BvlGxDUlFctz2W7J1Uti2jncEauZIIdu/XH+ppGPg69+8TwsSV
JooEyf65ZXFmkHpJe8sJCYZ5NJj2kvEGKrNFg7y7CUYOrTvhScE6OJiPsp2YdGER10UcemBN53xc
xb8tY3W2HrnNRtOkM9GiF4csb7570Uy4ToyWODlwrr+FdY29wLKeXsP0pENoEWMW6v4RImPRCjbW
6fF/hOOXPtO0UiGxHUdayM6Vtlzirykz+iGO9JJKyFLdwAmnk66JcV8VAEyX4DGpgphcIoUYrSt5
Sr/alSjHJXpNEqOWGUBjBNaxbhGuan917GfVmSSzLQNWKy5U52xni9KDqSNDlTxt3c7jSBWgXEws
UstKcEc9DFjK7/N4aIKeT2RLjmSgmT3/3aae6nIUPY+MLHarh677mdDWRuOBC/8fmRIlG3rdWAlX
NHlZqomoTWrPzn7f1XMBG4XIgYWLxRgBKa+RRCXCK1loXo/IPfmj2Cc8Hy8EcUY1x2mHSgTY82B/
z9YFkUdaSvD52AQpmCn98qx94yQKODNhpPV1FJ3bOCILB62JlVdzUHyziLE+jG6wG0I4CPruHmrm
nvo3r7x+hT98SXWf1fmBd9uioIMNafiENNghoiUCLZ6Vai5x2Wq33lHn5t1vFbSJB9OWIZcORN9S
pD1BJduESUhrB/+5LInPMkpoVVnvfzZZd2j9ttTjAA345/5EUQX8DH+wPDuXeYBk1snvCrI1Nxkd
uTlcOEpw3PVEVse3naV83FkZYf2gLabqn5ynTU+5TNINUPceFO/hf96GrULrwBuAsahyAYeHPqZN
FZgJHSZ93NNVOpupStS7UN1DLIrs/KdqXcf3C7kPv0HSFD517KmaVdd4ONtwV4O0sEVYx9v52c58
HoLRcxAyCU8yUhFHBfIcopyL3q2wxu+oqg9sJCEQOW33H6BKJZVgCSbXDI43Ar4M3H7ZMYs32Qrz
nT4LpE2YbPeXdLXxbXC7FQKN6DTzXiDa15tD/to55Z5hc5in6q/jxo0ZRwHfyDyZbWTwifELOW/n
ONFEk8qm5UEqvoXCBiKBLtmjWGKzfvhAPv4iEJs98O6HypCJU2RZojQBGSR1REpn16RrR+EgLBAb
bzKk68+A/qyNgMVHJScWkGaWdbJLtVnrOo6F9c9Tcju4qtcBOJdAG+ET97AZYHnrlGEngC/XIrOA
5vNOcyV0v+kcAYTduM4vPKNt2WF5OmsVIcl4IOQ2B7PPVBYY2JUQJxFWlBm7ksUAgTYbK3SFn9w1
l01X29VzHX75bfzD99EOA+PzB1VNgxG3UECequaFTBDllAiCqBRKjGweKj2/2VPVYIBNk6oP72wY
JNu4JnBLEE9ZmTvXtCg6nODQC5UHYDLpv5wtb+TOnR4mJGj9/UWU9IIRpcWnLn45d1/u1sYoJo7O
1sCIlNhg7PCFqncPfRrLm8pMJTjOE14th7JNolSvBGAG1w8KHkjHJopWBd6fHBtyqH+LJFAoxPTo
8tgcYUs1VF5caC5SsySM2q/FpUsML991obuCdewHUdXwoJWh4PIssjyfaiJJDV7nB4ztIYy6TYqG
SgLJKlTdojnLuBSyHpIBHb5caBWxN4Kdf0UTDysndhPHb1X+4cA+6X0OUth2j6uoPZahdbe0hTc9
6tnkRwIU/MGqdNLJ/Yz9E1gGkdmf6TVJDdTTbjCLYw2EF+wyR4Zer0mPbxXzGA+0aULKbmYZEjOJ
qaNEkxkhSZiLhO7I02/9exBxfXN0KAdHZYcSzhJJ+hS/YkF1AY7LkxkGhtiQTY0HS6nkC+q9y6Y2
aXCHp++9HA7sw2LrFmttlA2Oid7dRDfc/751sMZ5WHWtSrEB5S8l8Y8iqq94bfiqW1zx9g0QWGCN
j2bLZrps7mdIJCs1bvccBk2DddCGY/GXSuWbixSfebhVX69EhcaLw2EtVTH+gkHBSjduRdWpJWyR
DxVL51hIUIfP7TaBnpk6upGu/gS03zAzhTKu3NI+6Ou7DJB4cta6l6IQTKiA49H8Apk7VyjXl2X9
B0RH0IhiDukAMi5t2wJHm5/fMZKBxNFd5VK35YOUAodGzP39W3QW/fSMcxNLrJC6wHvr0UpPcXPd
ylUxdiPEyZNqi3+/dd9mnMLBO68ohh5tVytxPJQsJn1ZdUlz++epj5eGyJntAt5z5l2ijFjciHtr
N1+5pHvfzUHmNv4Aei2mKqOjkzgmgGZhH0z0kUIJwSSSpqTV3rE/03jvGvI3yA/7OrCJieLT7/i7
G3mAYn/Pmw3V12VPlBjk0dEugYXwdGwU9nHTJ5NbRh9YskoabQeSEvbCGJXzHAmPcBcIVZugAb4h
g0dnJ3AEcG5KBr9vOy8nhftLo8xpa6ESC1ush5hHqRyRViBf/EQLlmQtjvABp2f0sRR58O4Wy5fM
aElrhEFFhWvDLOTpXADdYCsQ1XGHEg791DBwDkDXTEVDTV+wEflNxBrqDd8vtlufF+yzurkyXhxg
Zl9/5JfS+SKHkB3SdlShE/wdKKHE1+b3k4U85PA3wRLNABF0xlceZiOdygWgMvhb0Cec51hKQzga
ltFw2k0oOgR+eVWB4JxqrS5RIAJhv15BkTpxALwwwHZW5WqQ66xyOBaSDSCMgzNOFH5FMXg4LABI
Ait0aH1qZM7MIfS2kiE83AD7HuFJtbUNftxswDi3+c5g0HWl3FtM3JerlBNLPeN6v/Ex4yT7J9YB
EsJNNhUSWDsaNF4k7fhQDhwS5P9uC2BWNmukHrB7KLFpgZFrPW1R6/nRoHLyDVhtMlP9E44gUaoz
RQb0B6OXDEMRopCsLUSzjILMaFxpKQk8FM5GB1RoVYHZz3q9cxkKegzo3Qvo8mVtIPVVpUKMiAC4
P64RGQo3OkiHsAwKBFLL9z6+hJ8WBNQXPlmVW/3mCh/TIl1TakCNyorIax7H+IMOXtAqm+Zc0FJV
QKHAkrr+dKNXGGU6VWJsAPKHy1OJuukRbXv5vEj94VB/0Si09ptWBvSbqIowbRsEe/Cx0UZCAJdD
mIiKx0s1M+vC6NClxYMtvI+WXPaAh2crxG3t98Sb/jtABUBH8U/9GhOqSh+L/tsFwPWfqUndfZOu
23jljei6qvkEu2tZmgwGHtGNKZhhS+Cg4kFwkVdhfTq8jRebI3EUUwMAf0cBCDCQ5bF/ppWeqi/G
HCGm+zcQ0vgpO1ulasum/f34BdHjyQMNy60hT9DtoSp77Z6S3jJgeykSeYopDAypZMIfI8wUcqEk
qsDc30K57a8kmWTUenfzcH0sXIYg1Xm70dWxaNewPgvm1Sjtsm+wfBL3AzYj7OKnCiOpEMufn5ny
i+02PWnJFmsK4l1YKAozXrNmMdr+eZv1CBynbdrqs5YW9jWqz08IqB42wCcdgLM04SgdVfsh7Vjp
imGNLchypBieLkNRddKYQjAaurXk7UwAFY8oa+4YtnYGFLtC0nLqDyGiDJQqzcaAkKIVaIB57X0k
p0RDiWqQBnTcp8nUMzKQY3Y/dyiBxcOM5O1SL8MRG5o66yvFp0COI1BlRAXA1q51qr5levOIgvHK
NqWpNzfHY/BZA9uu6bXufMLQVv0OuCqyG5iimyJyfjNk1t1KB+3IRaeW9t7gazV+jlEA8xvTx6AP
Tc3fWhCPfyVXNqIlamUndK6IxWvt5cN8XheZvQG/J9rU4vyYxUydw+DsiyLdv5J5qpUEl1NY1uh9
DqWLUDCzOcT2QdDBnvZQu7Gr/CH08LVAg2P51vbMyw96Ey9S34gRpOunlZWKEYvRG+rLoMDbmyCw
hosrh+OA1lZzSTVnMSUBl5ig/zxhqt4T3mnluyjoZmMzv/k3JCXS/r8m/bpPzTfv5UPAjPelJ6qz
vAPn3XOLrzkDGBh/XdsM73tYoRxL5HPCeWEUJ7p5CYkE8qE4CQgZuz+wtD5y//uyjGaa2v/oO+Pq
8CFUq6raPr6y2AaKAvUDwZ2n+tP4qUV8GO6/gbmsKfxSzq+cjtesk788ljS2oZTRZb3Xi/GAsMIW
EbiS5++TawpyNZcmNTcFo3iYfisGiKzZouNeHAmmCsZwknYkAZ34WUefAyIJO9fMHVjHrgwMwAvM
wsh8O2/P/SI5PdrqEeEcBFNyqKloC8wwu5JoN0qB7VAKOLua8leIma4h5ZkRvBOC4DMt07VeyXmq
Tcva8CkXCwD79rwnDUeo/FRR+p3NNC79f/QsSKU1vD5SCWstfpcOyyn+2OGA4j1dLHhXvQFLUP/V
aIcW399Z1aopZ4cgYy/ILoM8rZms3Lz2WoITmDIgOQ+w+uzZ7OMqwDcj4JoMMHlmPMwieggkgZ5v
ZRfAEleMORfo8ZoP3PTzGuhey71opj3my0rBtd6i5J40jVmEdQ3/wKYpTkrZUNDZnvpXoi1aXMdt
YoiV6o8HITLy7wDMIwrFI8LXAgaRXoRjQNuD8cv5ffmbZItuQqWVJrauxBpPdoPZNMpyeRVNXQPZ
6kE3qyQep1ppZdE0Y0mS2qzKJ3tSVRuDMGC3qH6FFKwnF+nWw9Kbt3fEBNDGwJqmdM/6HQmr4fWW
ikOkVh2IISyC0Q/x3JPLx9YMsG24sqxHvo03kl3sIjWsfsm1hyF8qHSHLNiA2mMUI5vDlUflU7tw
N9TCfx/+Gxj8RmFESSg4abYilAQ1V75m6qO7nzNHKqOwwbwFyw3hJH50yFYozy0o9dWeEFcdleUB
BZ4iG/qUOhYnP2cxPL16+UWRetpJKpswLYzCzXvhwLciA8UmEK9B5s984jgXVOheTIsdFh9aUjpv
Ec+wr/xhbg7FVn9owIjtooImiX5JD4RfTmAJkmaT05JFY1Zr588GhtjeEuh+LNcnGdMoC0hwkJBG
vOSyzaqWYnE5FOz5S1wRINGtSpnGQ/7AeMJ1X4rxBrRfHqPyBzA2qOFi58s53et4+Lu7HOYj7mjz
4AoRQhRA1G8pbvKINzNIMqWsL7KOsoo0qyexyGUq0Ns4clpAoSCDjCg0z5gZAdJzysn6F534eC+h
erDBunJBHYdU//fWrBaBS1d6qG+TdFaTLBfDMp7Sj1q25R9EEZpqA9aqNwu9mt4eS3RdBzdyzGPH
blEMZ0OP6onJV/EPjhm7tExrb8KB+G5YifI9wyxsuEyDpQkHJieFbjcg9eAbGv44jXoiOgwGxK7e
dTpQC9HHOoBzW8vu8Au8k2WKHWwVLLkVKEHgmZFvLRjJ1b0YjVUoM4d6qAsE0BNQiprSoQQrPrSs
RR9gd4OiK3whqXfpBbyagrZkRgHEHbcWfAitOg+VI9ST/jt8Jp3GMCFvzWXdxVTW/OafgN5IGjSW
HOM16B42fv9V7q3bv0BLa1QN7uVo6iyaIt7CFaMD/mGa2f42SAICD3HHA3kNQ9ED3EgnESlH6bqH
zze+308VQupuxEz7wlkorfhpxl1Kodw5YJ/Ql54D91GoCsrCk5p/Ys3YuWe2e2PxItwnYEg5UoeS
ZKa6+wEBrZXVrPMxuyHFcwn5/zftJq8atrwZrHNuNrYi8J5tInzOZjEGvHW2I6fODxIo0bCxiWXl
oM2jR0MuQahBSO99/lUB7eCRlDyIUef4LTdCceeSqzBXaqn/5NygpLXsE2ZuqsRvVGqVxX3m3aJ7
vUEeBoiVcu2GEv8NJlk62/s71lf9etFhtqjjRbQDDto1aYR7C9gaWEeHZLy7Vh9wB1eg1BmiTTLZ
p0OE8vWhi3rsb7S3sPvCWY/FCjyBxcm/ZUmHx+wVdjFWWNVzM8jMS0LjX3Xf7zwuunJ3OhCj+OOt
UrY86/QSxDxjgeqqkGARHqL9fvidNIeqzya21OS4+IbgcUhpXGZuFnxgdIxMyhbqsmUEZbXmbEK7
jIT9iSt/Lxu2sOFOJ7wsmZ1zJ7cEmzpitTmAIQMqTqNpbbKWTZAyrjhhqZ5yMedI/Zo2GHzJwhGR
eOsJkskOZ40Mf05SP1PgI31G3t/My3V1S2CTeUXzYmpBwpr73abiWjziDCrY4wSWI3CbPFpPPhjy
GYUCjWDL2JZdR6t/ED0X9dwLqPnLGyzlU9D8lYJtr096WTinG+a/eSnssrirmQobdXdOw12ibsqW
4ofdPjTfaSNkB5l+GqlQ8EzM5C6sTeyDsVuRNRdgkxiDm5lexw9bB61yk89M7/4IwD1Nq3cW4Gfi
nGAfy3oGxerDiLYdXQWZEn27YKZiqd0dxEG0bY03+qA6LYWGKs3XTMrSIE3bxM/ehhD9ZbSLpmmV
UDejgx3TkC+xmyGER3uCNhu9XGG8NX/n8/KRuoTKozxK+eJGAe+cO3LGWrueMGauqD7nUzy1x18P
NCZp4YPfvNaRmIOzUf2mFF9QJLNjImOHEDtWb+p8ScdFjCMAnR/+zwMhnQ+1L0GUDg3oEubml38g
MaM4QN9svcK3OWKeB9i5+kj6ijBsq0HR4Vg4rjrXH1hDflbjUrbvaAxq9GJEQTal4ej7ImaPfPz4
VxZ2TLZyXsRv8/gwDlKj8d81ERzxwANyCnDx69ILv5zy8iq8XhE98AvalJ8rbtYfUgciLf4s5fsG
WD3A1h9nOe8MnKvxW3++no9VMRuJQqwvGmj12KuVtpaz0R+x5HBmrVOL3KBaL1OkZbRZsyCGRfNA
Ms9DeBS8POk/aiTSJvDpCserX9sPxVZFm1UbF7KyBFXu3CffdO/mNjBu+lrsqM9uetCtEmogkq0j
H5Xl72X0xg10aB6dkwDBR+9n2bpSNATtJC8msTotoE0NcFgJ2SDlBdnYT6T32MtpYkIIGCZhayxO
CE6AIkRBM+PtvpWKmjCdisFA40xocxaCgzZx4PANCNLHeXZwaA4BG91M99qzzuGD2Tg3sHv7N782
kcpISJBtimeLSQgF//es8BoIlxieIjweOBWs2EXKCMUyPo5a0fbp4HgnH+zvk7OMDf+T4juXNUpw
DOY8CM37LOG2K3O1h13SVOVLlHp6chE7VLGwYtYR1L/LhYMuPUBdd3HPNAYiY2O1w/+9Pw8Fo256
mCxc3ax/27sR6CO+e9UUGjK1fLlOy2W7a5v77XKOi6j5k44i3xAHf09a5fT5fsdxgMN8Mpv9rW+o
2NgKWO1ketLVXCjLbqWz0WwlplEGeL48Zr1A95zCsrpqTHE3XRluOnUZon1cUXgX0Fk6Xmcuwmyg
QPqHsMlWN3S4g9chFGfL2ZynsURamm6b8LKOqP9gpufNAuobt6H6hADp4hQTaen6Z0/PoCEuyhJN
enLsJk2x69T0SOfTD2FSXCu6zEtkWz7ktFXVB6MCNeDZH6qfXuUtRAM8/rdkTfoyG6oWCKyuYrjt
ZZ+9lblnIVTqVUdgLBodmmpksgJzxxKlq42Tlh6YeubL0UxRDJeJEaQc6jwtj86GIz2XKl06+0rz
xooxZA3EmBCFz3Kgn9eltDqXBB8LQ4y9CmxIvjXLJIQhQcp4n4vzjwOpbfMzzBJhZVyWp1wIFzTW
BtisHBRUNHLZpFd7kS1TduOV9rvwDDad1XjCaxVeCVGL46ZXJwlqDk9YiKFm7285VgS5PpcLP8vI
I8JHnLjDWTNahtd+idlHkEd/K7BqhiePJDFnfzXCro1rNq5p1zo/TV0uXR+oz0ul5JJgrtPXs/cy
41lnwCwtVkuWvFQR3iio0JxwXP204qDtPyRT0duUkLJEe97em4VHLtf2kmypslVU9+rV/+94dS4Q
gWabG0uG/IUpCREFCqExwZrslyFeQFuyRdD3ngMcEViGQdnMa+iEevUwHCIvrGpMVsgp2micwg1v
lSQAXht/7fb89xNIpuIMEA4BnTAi11HpKWc0w16nUulYWn1Zqfm9639siASobqtAC8dm/xX9iNwv
MCcqXLSuRWmk8xwRISzhgo9Qdc7ZL9Vg7aDeIfMul4S0ZNEotrfp732XcXVQyhhcPIkhyBmTUYU/
wCGkGr4280eD8qvfIwe9HqUEPTjAwptOxvgmb4uhLsx0zFJlYpLcEasBaXZLRpDqYD4uaDMfgKWu
/JxJVWPVToPVjIit4NWz+kqwa4hFOtScBkqxKwQdKCjbVMwEDtwnRvcVuvY0Dd+35oX6V3q4tUcf
2QkT4xK951t6Cq5j6ZIOiFmkPgB5p46NbmrTQq/B3S3/7Y30kr8Q3yeug6N73kX+02szqoWGfhE3
FgsiKDSCseblK3PjgQrO9A+3rs/9GBdx7RhRveGAOSJ1xJFJcYLLCjBv6zMGhHPiBMVTDVp+gfz2
8ulBiLeinpPXs9u7V3bCbixW6wKO16XzSm2tOlkD+DwTTkdQSXK6NcQ4AX6NEKdGJ5YgK1zCUmyg
MHwhSSR1ZE7Em56kjCPRAQgbODiO8I1gYecPsMzfHroB/jAah5IGW8TMzAVYr1bMsaaDuxv2FDFh
dxi6JHJYGX4WL55AnMb8j9vvKY24j9RWtfcw2zMZVJp2tlazylFbgahKR+Qli/VAoVnJrlxqS1mb
+bPWNjJm3w2x0wMqyLcB9Rb7LJwiPYlgg3rwr9eDGcXagN54O12XF9IfKDcfXLFwIzxe2ttE8F2i
vNl7mkOolpGeT39Xd++HtcYb5k+I7bx/JZevTpUBnQxazPdKmF5wmublZxnczf/qtOqjK8tq+aZi
Zjah3eKGvoolTY2q/d3celiMfzA9gOKifaCTpLMVReUGy4RJnJmwrXHhsmg8arzH7ijqp3INYIMI
W/QnTtrP3K26lIqMHuUcn7hO0uIgU54H04ztFcpjE0pgciGbC05zNkAmGsJEhLYR0D7odRhlMxDT
epqXP3oUT89Czpolq1NUz3Vw7jHJgwxySSvBB8mhKchjpklqetYN6AZUP1qfxQHQ6vVllg2vTTaN
RqZlAMFpF1LgKM/WXaBI3nM+rXt6Iy3j75M4n1HYprJkMfyMJEWDLnUAdDtllWR+S6jG+P8mkOAq
Jzc0HRr5tjYiE155jBuuqgWMbvJ7XcU/x3j/kSz8QhiYxYZhha47YdIrFL/P3XC88ReAT+3cDfwY
5EWiMX4TM+HVvosyrZRL1fpCpEG8yMG+3RUR1w1YB3hyvTbD3clM+YCbHPdGbVG2Dj3JHf6CI1N2
OVItwPz1jSxu8ihQ4gyrCnEHIn9hZzJ47/61FuaBqgA4kdoQeUr7mk3bhxTMwIHJcRTiwY8bDQKr
bJtkeQ5qOOvtDvWpkpViM6ML77BoXrFYCKHIKNZJjrRClVneVhLHSKT/2lyVwLxCJGodefcPo1qJ
sPTu9I9MaWMKIVF7EM3pwwI2jERICmv8fV8MP2K4369LhoJ8S7CzsR0Bwo6C1bWSphsz3cVMT0Dm
BGO9W7ymQIhw/LNqZh5R0WuSl6CfS6UR1xC2tmgdAl9tGhqMDLlyTx/lsVgQ7gsVqpIW6Jy5t57+
IJVyBFgsnSG63yEhEwpGmNfEHTWJo+PlseIWxlRqqiCWn9SuzI2z9UXVYkDEDgM+dFHZnZsSrO3D
S44XY6JslA4zwpW5LcGv5znrT7W+/DOndXZOgfnHjrr3X4HpNun6QZrUUe/k84YWidcGl+F/3bHS
Uv/3/rHDvwcnjPJqnmk3JLCVSJ8Brigb/7Y8pdlbk2Jfl7afvBu6yR7ElkxEDkfUGQBF87tkdjDg
KyfFOu7iI62+5Ujam9GIK6cpK2BSBZrXgkpn4op25k2fxNE2sis4G1f11zyqJmB5YK7tLI55Hfo9
lQwIYX09a1WDnnD/2N4aRmVVPRPv2bmWTYki8loRqoV9PZbgD9YHgZM2j24dBA+A51MC35cTcSHA
3YJ+pgfG3STQrnWzxeUiUb87Yd7Ubk3zZ9k1QwdvTWu4ZGzd8cclwx+GH8m/AFsnllRyt8hARCQU
J8ZiU52rjwvU51dmzUy4hK2gjpo/vvNChr6BA11KPJIgXh+2v8ThxsQm9e2h30l1L7kwhuaZayDc
hiR/7suvN2B/VbS1Y6NCgLBGaPTkH8EoUaZmoA1LQkufxa5fzzYdTBn6OiEtojeyz/Xbc4rFahag
oPtepyK1QpHU8OgaWtD3Y65Y+Vi1TebW19Zrlbc+hz5lymk6lrQpqUKrpq2Mm9p+DwqltPB+dpxv
UHGsDL051EZ6ofQkkJzSpmba+JXbIlisXsJ7wdCYfsJcogvWzFCaMniue0ZntzygZpVWs5xl65DR
JM6Qbt8KZ81mCoQgEC5OmcfJGW+npfbJ+EVlTtQS9nYEDl7GIhoaFRoSoihMexygwEkHOmdnJ+Mt
wAKaxk4416nxHbyFPPW+FISNDL79TcXjopziE5Zxi2cUatipA71xLkDE18lV5QXWw1hS4N+iwok+
uJ1nyaHvaoVr0QGQKZb++mG7kkYJhr40hUS2nbjuR+tXXE9vCSftQnO5708T+aMWnH605kLRkVLV
gZoWr1mrWRYcgNPUlDua67J7xvrPpf2m+lDhWthdBpz+ce877DQtquI9CfaefwDXlDIZSRTpDdsS
w9MgUINukRI8xopv4fCQ0Nzf3lLyMf1iFpNk1dT31vQT8/vuqAi7BJtAa7L+1v2Wf21toJD6QzKR
pYkW47sAMWqBLCKqe5zk6LXiko6Z5gNb2PVDQiI4LH/1wD9lQgWZivJylragd1NzlIkcWrB0wNge
AZih1FavDbxOK4sLJX9jDGHa5sYWmfzc99ksEfsMqj9eG2iKU199sqUW3Gsvwc4IsYkMgINTq1pJ
uFz5kLv5Mq/MUeiwBC6ty1oGGJ7ggcRssLNITNex49YxvqHb+E6H674Uml+HSHAfYV5fpksqyxnV
mU3AiMPW7KvdQOVk0pNSks5ME0erVqBLnXGGTcG22fow2MVoJoDH4EUhk4jk4b+Hei0aec8Jo07E
gVxu4kLez9awnv9YNvmczxB1MSdrYhuah2Q5RuSA+iACds7oyVWMX5cjMxj5pkzLG2axskh/uYwj
b3gRoBzfBTNeKIsbJ6AXUcv/2vf+D07GCaCztoFnsCCOPvq6hgLrwvJ8Kw9SqfxIYjRbuJR+2Hsk
6oX01QDtlkQSI0AosL0NKmzXDRiSZuKyDI2Jd1bMZsnuyrBep7bMS5RDPHdr4XFd83AEV6el8p1h
PyEfw49qD3nNcFWipHZDc4pPNFGS318DN7ILNvj9CisRIZo524+LCa5HGep7HNckxB+sLW8f1Hf4
P8ZdbrrlWMOc5w48CrIKHZpPvxMy6bjTKp4etQZQs/AMtNnQGTvrAIJ1rmTJxtDGPkno82h8D38q
OXc002klbdZTvw3S8W5taZWk8nStXnpgUN8WKAC/PKzUvZm1Ol5UAbuzsFQ2SRI8SyloNDu8ROAl
Xg8x1dyTWbiGudtVEQOQ7Sry7wbHsAfr/sSWD516x22cJvScRWi9o+bhJ3ZRtMvF8grqVzFovBRm
A2i+zhc3iM/NOLbagxn04gYJvPztDb0UVXOFb05y1xQy1YsOc+favpPmNHX546cuYeUmtATaAhGt
ITDXPNQE+XrWU4fcTo2f4Je/UNO3SErxy2Q0ajfYuxdLRtKyLjO50iZwnF2vz00gaa6d5VD17lOX
W1zIBkiv+upKnWUt5eY/renjZaFPpWP8BKH1OuqLG2TsKTywEcZidDZb9H/uxkenVj38uD6TzTt+
vry6lJq8PtY48DK+bwLlqxZjW/f06s7DpPijqvRBb0xH68Ursbi8hwiQnlqXDpmTzx+HAqUquDt/
31ugMW4pBmzLW3NKq1P0bhBP3YTnva2ZrobPJMHwJKIjH1GTKhPRH/FA+aysUkg5cAwbwKyEKIo3
kFcwxX2hmbRggBmIQUqnaBY5oWEywhZsCh9QwPq/91BjSWiTvIta0r63+CXV8sGYdL91kE8r5QOO
wVXZiCsVoiKBGc/YSScQIZOnrqNp7H6n2SQyvpZggtWCZ6Wh4jpdLw+/jgQZ3W9rYOCrNAJcJXu3
lsdAJL8X9aBzoN6dSVzyX6BpaBV1SEcUKTDZbdgo5cZWOG3kH81PTuyveLcBKk0y4lbwcJKDX67b
+uXUhNzqlzTcd7bTYqloXXPDbBlxzVdJt77QmY3oewTo49JLsoJm7Kq/JlFET15jZ8Wg1HZ3zUiC
8fXs4exkCZPgWFQMFzocs5swIwubeNEqyk2Wq4MXf/Meh5MnttM2RXtSQaG+g0Old82wT3FmnZAO
81mRx4fjxanInY5aVve4dpdcydgxtgAM5zFEGLOKVJdvD6KaDBpKaCyeDvPcvi5Jp7x5ZcSWIE8U
f7XKSaPEMaxn5FKpqvkJK/GZgn6XseENm5BaP8Zr8uWt1NWQNFttxeikpkOvgnIq9nTRw+JjEZip
UZH3CBcLSWBJhCEhe5sTbuKnFrejUo60nGIhp8CC9AlUxTmuI2H/Thu8Kl4EwlIkj9ZeaC1gV9lD
gCVKaGY9yIuP36e2Y3WLpSQz7PIZh1rmCfsO8yh/WtSAc+OtyO/NBGXO22dz4YdtX4VbAFtQT9h8
01/J2sVmKJSuxpvrgc/yKjve1/zQpBdy6hydCmMMSsB98+4OoUiVoz2RsBXcYIapZH5rQWp8idKY
fJICGS+nCgtzR84jVyjYOMJ5TwhuSsJHGgdnM5RBu2ZVD97jdwnRqIMnjJzQxSRaodXlD5SS8PMy
fdPeSVSrSjXQG914F5tL9s4Y8OaFh5s0ylCMHhsmQSLbu5OXTofGwC/5OfnhzOlFNrgz5KXmUkho
XgX+7C3hqQNCEGyIk3FzLEZlOeGExyTRLiFbW/FWrS8qFEhFr+F8R6vME8f+sjljBSYRyAvZRSz8
360p/r3rTXKVgDYkrxwgY9samamKcIsIYF3x7Aru/Y6M8Gr8+0qd4U/VdwQsUqioDZbSq8RuBBV0
2yoHLrCDU3m7qcDv4DCRB2ps8yiqowja2EHjWE3GEjX4Wx2xrZMjXatxS7kDpmaDG9RIXPOcHKm8
uapxMfPoDXwazfbefI6uQIyhHsRbGCEz/cNth11EUxhBKADAU6SEE8l3cMLiiu8+ZBg5YMa6Fn7Z
uUjYW0bcuO4cPH2SBw9YqNoASZw3Nynmg/zL5BiVonK4mTys2pA5iiZbuckSm3ov4hhnsnuObqdX
SX0pQ4eaWUFuAfYdtTSCOGlVVGSrCDGCHu1lfNs2m685qCL1OzQsovLtULbuf94GfP3tyMMS7ySP
aSSUo6q+f3HLzhczc/sEVLS7joZrw2OAsIG0/lMQ6+XCQssYgwnZNzEAOOw3rKTdSbB1hOVxBomj
qlseqDd5N4021lgbiw5TVaDPUy+e2UAlmZLr+MqHk3cFgBONy2Q4SPq56s4eM7p0GHc12P5dTHqk
UENtTkG/rHlcVE/8xvtna3XEmDY6XkHNoFphI4+M2nGb0uAfji0EtSiE9NsMntAa5wk7MOiwKTyt
N4IIZZIdojTzUgGWGxPU3f7brREVsAC4WlKRdGqieT40OSEBZ0FdA6QiHnAuZjld+ETfBj3z8lk9
S4n8oXYxnzpy1i5ZgfJ0BejI96G4xl5lXuCMrCWoYneT9t4YJt46a2a7EkB/hpdwJH6xyRNJlQpx
Sdf5oJe9uqFji2SKV/brI42TZKs0+7SO5oTdNA73tOkpCdFKylNcckOK4lrz35PUn+mv0mItUNK7
08c9H57Dn5FBLt+2ZVuiyh2qn/t6UaCVCUqpoEdCydRjXNIEeiCVuj58SaLjfdo7xWbFjsysORdz
NZpCIol3rR4wAgHdMOqioX8xX6x3ycLuZk7Lg8/KEFmGuMuwjD4vRQuQeuT2GHhQxF9Szfl9r4oJ
c+X+XXMaJ76xAxMJr1TVicJczmKPreKftar5g1x8dOxP5dQeNthTKBxEJvJoKaikLZBL0nfMOUop
vhvvMnpJFHjHHGjL4bYD8FHwmDhptHqhPw8OhWRLBpwDXx55RzV5d+A4jVReBHG1pcCVJSfbYCwg
GbFHzPQNvt43XkZo7MqDdEBCzumPEe3xgUBPBK5DplEixcpwQImLXJZaFNXz7njKaOuEjUVMbtBQ
uvEbhNSh9D2aonHdIYxku/WMqVTEF8DBWC6k16s77N7LywV9WRBID0YeTFVRacFHohomutdqQAa9
uwaow7g1HqWWN0DfdP+nCQqLH+lZITUpXK2nFTSgDQKtjYJfb6npcAk/4Dbmn4IHK16sgeCbXv6S
7ZjNRPq7MfUi2icjRK2Oqs9DzMYo7Cko8Ihh13BtDThBSufquFJtWgE2qyvpPc+W/sg5mMkAFjni
f30JR/3wJLMagGScKm6mmTDdW5xgcc43jeToj3lNuU9LllR40g1soE8ns3X43b9z9jaffnlevuLQ
THSN8dwF3WIIl7OdPUUuSkOkl4EVdT1HOybf8+diNCXXspcOyD8J/Emem18k0f0h80J6QdjO4mCf
BUQ23UEdzAwFQlqrD8dmDutp1a26NVxwgaMw3nbyc3zD7FKmIgpAOrOPq36Cq5T7U2PVNIPCLWTl
U+bGYR2vlGJ8LSDVxH4kkMdftaq+9LyulWYCIPZKVmBL5Ha32UDmuUKjkPg6irQgNeKdmGc9h5rS
wgIo0qpBaQXn1Po5Lrtye2a4ZzwmJGqxrT0+ZS9+Olay/cXHFzJU6UZl3KxiJamcMrQKeL1uptNg
7V4mMQvjGirFosoA4Av/VnJ4xzOVo39e1YFmaYX2DUINqbEfttxFrb2BbslAKfHrSxqbqfbfkJ9D
XwhwNqgfkUTIbHx4Gq7qLcn1dqn2e74Cxy3g56IXiCKJaeQJuT5+92aGSGci7vuS8O0CGRO66Egu
NQ8Vuot8SVmKRXYtdb6x0Xj74Va9DpTjJmWsOpnIZGsOqhUnyaWOWn2gQMBKYFCCEzUhJrViDan1
DSiQLeNxrFr+ocnU0Y4FJC9RTE6G+O9dvGmi14Hu+yxlxHHBM3c1tEPv0kD7acI1Whnpc2HvGinm
fQa+QyHTnOdxv9RhtXw1tYsT6ATA7EI4pV763/z29mug91pW/q6Wi/or8G/luShqboqCN7a+zGIh
oTH8/o/O9Zk6Hs/3/WHT0GtYJXmoabfONVaoCWbeN4ISouEpeYaUvcD1OU6RKKCtPl+1pgPfgFE6
OuwYKj+py0YPScBQ/VjiPwtS55BTATNY2QMeUHxxTC7sQuvjiHmzd2cGzfmsnGt8nvxAdmEWEB2s
S8R704tQvfoZNU0deKyNzRI1rcpCbh080g6i49IonkkrkG0qqztD0185E/Ta860xOXHlxlns3nNG
w0BC8J/2I/8khLCxzuacxSovcGsBc4xt7QYselzPmcB2pVqteQUCRS0pFmeW3yVtam5/q8EHrQs1
GL08apRUK2ud7x5g9lW8w/XHknpIOUb2W5ti70Z8bUuA1Egc/vkpYeoLtwg2uBOwZg9BfHST0aBY
bHTB1AvJ5OALAyjgMrTgthd0QUxWD4wnvvdCaABLNGIUZNSKAOtyYrHVQuXAr7zO4hPK6rvWl3pY
If34HlB/w1j7FtENFX+nXnmQGs8QWgpYnewsErUyaKwo5p/ZxLXketB5jCPgr99rTJbZdmVlQehP
6Gv7lep5nsw1nrW4njxAScBfmsotCcBdiizUB8qV316ZyevFGC2fkL1AWp/BnLynJbysXGFa1liy
j2u13W+AZAFAL1UiB2qcNVtjype+d3mnT/kwlewYkJnPBgz+4sNYvO+1sZrJbrYHpupb9BKgxArx
YyDWbmzfRlXJ7KnYrNpM76ycEbSsfZ/6ii1dW6LpbDKlSmUKV5uR9wpUzzJqdRm78HDK9xRE5tPq
kOVUePV//fzEUaZ+3SUkQZowbkuMOY0PxWJv9AjITAfypYzbGtxbaK6lMCq7Ybh8C1wpoX+94sYY
ak0Yt37kE2f5fydr0FeVC+xxO8mBE7F5DSW2+4N8O7imKifsLJ7utdYGZe0GSUUgLwcmbt7asQuz
2hi9B20Jwrjg3XPvoS9Q1VnaLarWQ/rNC0BBrG8Wh48AiH95u0BYPAog1A3pUEUCBq2ygOLcTyrB
qYevBzi+Ps8wbTbe8QNrj8lmdUKPW7LiUg9I6xOOJZfS3ZfwFXartpMr81v21rZ2Ks6RnqkgHIzO
vpUiupDFTKkMbj218Lwu5MatA525Uosxm9fyMbRHB7fXKRUw2g3GcEjlNwRq7Sq4/0XXVDBJZ+6z
gjKAcyqgJFyrXAUC/+VxXvuC3m7vp5vBr/S6NP94nZ0vU0k6xLZ4HhpqJiDM9QBVYiFjccKNaS4P
8Bb0lWFYuPyw2rSXgHlwvgLdnAEh8BQ+H1Eao4Ttzb4nS455rH1yQ9uxuuL67CkNdgStG5kDIWWJ
hXhGlrblXrtWtwJwva7uHrbmTGYVgAMAMMpAvYCvfJmPGg3WZlFMpjcL62HRb4E8QgfoWyqFnpTj
f3VOgtZ4BYEPHGodMUX/NXYCqwVXeRytx+e9NXxzchgArJuTmPlxCc5aHFQqCUsuSwNfZbvEvJz6
EASSE13WeMd2Ad3lU/bRKr3mHsLf3ER3IrgGac3CvDbcWoNow9O1GU+gmj4TcXA0KdSsUpMKcbr5
6quiLjSrQOk/vaPiVgGEDo5cB9fiL+ao9PPyaKG2VxPzME25Ay81DUlrD8h5f+CMG1Mz/0DhmoO0
Gq3RgYMFWE6yx1sAmjktlMf/1dnm6JqHRMO0bTvMoZrsAINnvVTasTcOuHD0ErUugnYWuzBu8Ykx
IfNKzAuH951rh7lGVNM3D8M4nNWauAzZDR7yg23FKNry05euhE/bT/X09cW6qcxM6EAcDMWrPAzd
R5eIQrxqGW7tMvLJVzgA499YxGuE+tE3PzlzCdQPQw2W2VxsfnDnL/ll0RaZES/c5/idcpLULbWs
j1Orf22PHFWcul1i1pjuLXReYgGm6YPdRbVfq59r4ut6vNzQbL5ut5qPni1ttTYrOUSgePYrrq53
sC9F2kbIS9lMhzycxBFXrd7eEK/YABpvqgngedxgtp4pItvXapP7UwDj1JHKeoyhQpZ9g1wLfTQd
Lfh6gjbQDKE5x7n9v2ELXFrhyp5IRrE/z2KUKNlUEYUGEkhcklR4nsoaxnbBwl+s0ua2My6keBTs
QvNtDeCjjMOB/qIhwiJ/LaDMu1bfzVG7RPOaq6br91el19VJzeinI7CvNGwo5O6fXf3n4sZku6ek
yoCYOuv8MRp4iyxamy+Vaqz9A5rhFowQJj4YIxMMI3mTN/RKjiA2QiCv4wnfU/o0G5oI5XW3LV/q
xCOV+638lNxTB7/mSsiaLcMIyYwCCnKnvd+z7o/P2V/eQl4dcWeX3TCrOxaxeqtcfSFDDDuOMNgG
7e6qXL7k6hGXJI9Pw5N0UjcJQJBqZW3kfKrgV8wwja7gct7J2llp072G9ZPhgK/0yVbJRuKDpfmW
o4qw4IiVu+kxIjN2Ff8xH+1V6/CmDmjm2sOezGntEcewopX6TomfG0sQxi1E3OSjiZKYCOxRyEl4
Hz+rTXTg1I9uflHG31o+yIG9w6DKA3v8Ba+qlYDL/1PpgPJ3Zg8yA9CIkvqrUjYJDFEU/6t1KpEc
Lhvc6X6vuA4IcLZky2NnA7PqsrP9nS3YXZ09DVZFYHAmQZY8rqInCYWOl+snXl63l0cdgzXwuXxH
C4iX4B0pHFer3rdhLj7F5d47wBrw56UwMY4tHvyO1e1yHAjo+CzuzbyRf6HsOqs1Q3LUPp3Y0krL
ZhgtCdnkP/v3PcTMkPtYDC/6YYLab4/QqoTM8W8HeGJZhwlTAaL+lwxGwgR8+Es1HPEzb9I1V4vu
1w5HnBPMQIeq14Lw2FWTXI+Uscwwsoxu/8S0GY0ucr27eLG1b7U0+6dTY8GLggGn5ylb4pkUwT7l
okl5Lnsx/63KA+6Ls45GauQp04s2RI7OYmO6p2pULGwSSh1kviw6K1GjU62pYjVLZrCfy8DqkHH6
7d+9GuSSiirT6u7WcTN/OirQCmKEsguJaDBuMg5bP6ncGkZiOkYqxkSSJyj9AzqWofRPGFNzL8AC
h/vy5p39ULrPZYOLXwZN+omvVz2sgCoM7p/tyPKpAAIT3z3h8NTwlW28tzvJ+p92MmfzNOW0G694
qTPQkXySpvGVHqt4taickXMIVCR/rmuQ/BdztmlV9kouAECZVYbxS0kugXpvH0qzzqF3Vy60TZBl
8qpQQ6rq+Pu23YmYeLFbQ/54VOxW7F35+wRZSKYrB553TEPdjVnwwOwpAvxR46GCa3RVlity3shJ
/E3zkJlJa2YSTyeWZbJ/yoiJpzzPoMCCdiSOo3iGY7rf2h6y+K3B91bcjhxP1MluqZ4SH++WiQ4W
NbE5x2fU9dW3CjxNVCRytFMUBJH48HWaMj7ireJ1upsDGXUSwRYbupd6Z1S74rVEC9Pn2AQ9eVsA
uKDfCTHsgizQ9LPuCZWENyvDwavZvZbxutOO3mPfX7eIRdnmpm/YQtcILU/IFrQlwNC4P9suo35X
UvRGNoeHjcPF3veWCTwNILfbH5wUVwksH7h2EWMG0vM5xiwLzYANa6Xm1i8Se2OJx5fR0fXCLHc8
neThowyfTfQTRqlKoi3N74F2tYtMibVrZhDS8bgzqoO+pmCGe/A7OADC8A3NSibXaeP8lah0gd3b
Xj8rJ7rCfS/u3sk52uuPZ54PMVTmF8CPq0w2wmGJ//U6+yvzoxDObTTZtvuKFaleGZhQ1srpAjw4
6kzXukbcA0zgyly2yO4jMePrkQ5OTht1WaduHhc419McGwMqBIlDODB+7eh64+J8XOvexWPlHiaH
jik+8YMgDbV2TYdxGDZE7y7YbL95qLfDnsb2tgteOu+uVp1tUtB90oEFZLfUhLpdiAleTqwWNWX/
x7fWL+ScaZsRXYtpQ4zecc/2vojDNjJ/yA+fZJyNTLJHCxjkHP7urfwCD3JV5WRrYkymvu6j8xMB
LE5ENdym5Mc9V3BRKJambEr58empEo8dVD0leZRgziOgRS4xzC9BD5SQgXHfaJlRCj/sEMLwNFQE
Fs/tGE+XspIxYHyAxjlGWqmdrXOgdxngd10PuVveSxy9cxcSsESnF+BYc4r9AGiM1b7OLunY400i
i8syPs+1x1fjkrs9SblPagL6Tt5OZRj2yiC9qGcUkRIilTBvT+n05NMB3I67DPm6YMtPlpNas08e
DWKb9PntNbAXs9JKKJwRqagow+8ImZdRBXQ3SiW8qohqQB36QNE5yzOhkVdmpKp7w+eNPRtofFrW
vTMHIsWnOU9lwT091yT2+xeiN8ZtZp2TXLwTfWVEJDc6KkLIGmTzwRfrcqV3jEQysJCvBtOA8C9v
26mNJCNHyu29h/40gtEa1C0zu6MK63CDjiR8p3IKpnUK7CqRgJ26IXa98WsFZJjvQ3dPGDpwAXQR
DxPiiBOnzAZYOhzus/H4LsDTf3CVfWsgA3tdY+rKCyFlG6nCMIoXZ1eb4xpTArylgu8Jy+kWUkvR
SKez0HUejZ0snygzKCWVUo4yTB94xx7Zoi/2Ku6kURomPA/kE172hdtBE+5vWz4QoiYewdLDu7a9
h1hpwnhb5/CLYLPg85nOhFjJ41HKisYTqWS1HhhhZDj0kOC/omxOjOIj8w5txycx67i2EgaLYo6X
P578toAf74Z0kK+PRf2N2sFip6ZrWehNJPs1XFebzBO8UbWslfGw4TRZQGalgCt+QF7zsxWisjY6
D7+O/dmBWSgnI6DAq0Oe8Nib1Wnf/3IfAlWsaQ2q1fiwcekzdOM2PV/XxcCmw3j5Frfjr+nkw9fv
FMTl8UtdzFTSZ6z3K+nvFMEquTfP6JJxZZGcCuZexKY3WeSYawLy6hR0ZABtSowN4TAK9AnTO5r8
izoSND62ZWpg6Nni8tacL9plEtnHHH5aTpSbGCEMnL79D2AVc+eKe36SVVxYLSwMjkoANvr6bWdC
RYhfrOczLcm5u35d4tSK2rzfpLQ9TyJMISjODNVXzvjYVgDyngK+tJRtaiwI8+goSH5y4aUU6QJh
R0J8oVP4No/DWTo2XSFguSBlCxYF5zM1ks43xQFv7TsmV9IkHgCxJrmScVO7nmzhdpnc8P2Oc8SZ
FtHuph0C+5KnMfgPHwUwar1IypJnzhGPEMcwExoP2f3PY3Yw7nqpHxSc56IuokiScntXBXiT+q4Q
g54v4L3XxcIvPnV0rZqUOQ+HxpdN1ZRnB5Gqqk9tHtGNcbSIvblsjkzGQdz8fkhIYiqzr7f854eu
lmSvUI7D7t3qDMSRV3wWDeGNlSgdQZ9rdt0Ag0z3YvSCehihpwCHQSGJo8xIcbwpJQnSS3XbYNks
IpZNFZTlI/a1+dUMZOlQghffLuXX3uwhskmr6FAOTEEzkjkoy9lFprD8JeXmP3Gt/TVIsMcbefzr
avGj/jnT1WTdrm0k/sHibJtid/P1yIkOZZZKoLKFuVj2ixw20lKXobkUAOZrf1Te4eP8RSqybJv7
yfk1QVh/jarXpcvS8ILdwCfWcqFKkCV6y2ma95pmV2JPw0eqekE0S2fURjsffvvg9h7fqJOdfSg9
lAabSmLwMv1PtaQJHJoG+GLY39dszBvZJfsQpszzDJuKshlnYB+i26vrkcKV0aSh6JeOzsy4RdT9
OIr2V/vb4skAARsSU7wcfQRa2Muy2499SBt4sApm2UChfAF6rGqyOAblJvMwJ5c/MZJTCoCpSwuH
HpHy65+Za3LMiqFD3x4yqUmD9d0+hUBMcIPo+263RFk8tqM6MVp+zogVqLnQjCQqFc6zMdAn++yf
x8YrVvgUsc6yrUcImis/+t2zTJxrAlLvOs2l9eM7LAvMebs2ecrcUoAh50uEMVGHPh7ZdDh4IZCs
v49al8DvcH6I+wyd7YklNpgT4lAGaGOvhFOyidAZg8MyBYitJ4JAltu/04Vu/DbeHaSh5pUWx5Ye
GdxquGd4jkTxs17J2/gswqDobR1nHzp1Ld3kZXonalg8dhVU8w6MWEJx0/ENayzN4XHRqWaw8Ovt
wkO3HiZ0veqqUI3y7xJ5Ftd5fqlVqFG9MVd2H7hP53rJgdauZLthmKk4OjshWgbkIbfMFED+0kzu
KmLbwO+KoqWT9eUiwDXqsu/uCCLcrvFRGlDFYEUjAoC7bGQ4HilSGSLTYGRkFn9UlxYaXr5QkD0T
LLRUoAhhv+M4BueiG7sBxP1X5yNa5AHN/dqlpIhjJHb/4CJREA0SqH5PMjPJ49r6r189v7opF2QR
9sfYVGPpnd9/gmqq3RsXzqG9gMWf6aezbsID9z6JzOQuEw6cWANNSp782+wHtg11vmkWd5+bncXr
wsqVG4eEnZ0nkGGYC2qY9AG10tg2vnL583dFPKUfQY0XhZWUPTwfLIRha7OXJJxZQpbDqh+u0qXW
ZpidJ7jQpUIrCUZHQLstm+wuIQgn4igozVQXCHYiSXe1a9UMMd9HoI8/7rAn2FchZraRKTB/kB0q
vbZV/mYVimCxBxuFXJ9QsksxBiEXF69JT8ZUINZo4k3ONCIe2hfyXh0acJqI/HPkIfMTyL6wLxrJ
53imtsPWWNpHZBwR1e0U6Kh7G9FmVYlMIdbkHdqjun8qcifb3pG947v6jWI0Yam4/DrJJ+QS/FVb
NXOjf6nZJiz/0WOSDLdsf7Anv1zdM8Zlk3kW0wOfwuG4oF2QRt2TspPyrDpAnGi1nuA2BA+3mvBP
yHZHksGbBYSXvov0jYcz9n4NOVcbzce0gjPcFmQCFRh4ZsjunZd4l4pecBJpbcd139enxouHd+5Q
s9MW84sazzxf36jzXRaWhXWbYtXIoO85TwceUA6lEVPvBQqSNU5Ynnv6fWjMH3f1t50l+qg5flfw
mzvTm/VD3tW8Is9HvKWH9tEJ4MJ8r0UF6NQifg8rbL0j//RB0YbcGsH5kCTIFWlwKTNWrpvP7kkC
uOg9uI3wUb3bwzpveBTCXOOiEI5OvzYWTy52B7KF2VIPYTJkbqxIGvRNpT0oTIt4xxxO7bVLzrbA
PizzD6iF1xjp+wupZoX4GG0WlD+mVA9B24kGH0zNBFLWIm3U2sPyeBDIN8ews+5S1DQCgOtmUHwl
S+sPHme+caJfeZF3xm94Btm6ObOTGpHQrB8nOLN3XmllOdSrzDSzAGuUC+HdvvPA6tA4n8Y1zhZk
8hKMmUbcTsP4DNoITT9IjA/69ZdqrvxLwETSpPraF395MZj2bNoGG+5g9dkR2y85+8SJl6QP9JmV
FtPdTbeJnypjdXI2hxYL7HmOCn3u9hzZn26OHZngYUYUkb42cHuscU5YHWxtEWM/WDxUyig0MIzv
fK5ibbWvx926LhMERJ1R1xWCEFxC1LjDC1Pp6z/GCcMWVbnky2aWQpbYr6o3QBNEBf/Oi/1BVYf4
R56tY7jMYM2TcSUrQUEFP4HET4JTK8+5Ov+gPxnGrH77d32oF++RKfDDBdbsBA7aPz6zH8eaHEjs
GsMa6fNFKgc7q3JkcSLslcxrcwfdSWBcp7s4otL2pFVjHtTi5BLm9K8ucNpmp6na9XM6NeDgpvxS
k2gba8tU+4vmgllVpuMt2QggCoxFDEq7JlWTxsNi1EMYZRgb1UTWmDTnnaeEQZKddMG7hSiwp4L+
IGUMErprqDaoewmO6klIKA83wH3BVPab68S8a8XNW2UDuI7ZzbSwamGg8gTb9QJC97YkhkQYLGA1
YrOJ+BTpP0Ia0F5kEmo2zVX/Y3exhRSGi+MLSkC2BQrsuUb4X6JOlpPiTPzGRK2XBlub2Wlud+KI
BdINJJOG38qnmsCLwA/3rSe1rbEH7IOQHOXUNUgFlyPzkx5BWsMlX1t4xsqgV0nNG0RKCgR75v45
SvtJyf4kNnjKN8+Nz5l/Z4OM7XXWe39RmGibGiSvPo306qj85tVzg1h6HQ3iSqfX+KckU9uwHUsY
KGD0PWALoDzpN8ImF5U6sCCXBpYhPKinf484PckBZ6AqNyWgRujYgJtyYvWw8IN1N/UnN1Piy6Pw
ulYg8uwXMScvyIpwkSzAk5Kex+cNECxuN3bPEcOEqVDRKNfCw+/VHXJwoJ/efeiACH9wkBHGJ2jY
efPOiHxPXMEhedMebow8bJfB/FazP2cRo0AKgtwXNdWStzZoIl3M6HM9RV3CrC1tQCvbFjs/3RAE
yFM5BYE8xeJoUkmPMh4e8+eBVgHAcERN5j3JRG9bDeiuhWXGtecH2iMIQWdsZ/8QanGTjk6I6Zp/
rVtORiV/rGrYqugk0s7fRxjqrTtEbCKU46iywqtrlZ3CISieIUSSGx9PExSBeCPHMf5ww3FRQVH0
x/o35x6nLFIA7XWWId6PX5Eh9tucOuvz++Utr9Gt2DXOlklPoaSjr4YUkSa4MrKprTjxj3ozBzNr
UpqkoclpIsyD3pk1G1zlRMFH70D/9RojmTM1hLHiAxsLS1/fUSwwUE4F5YuYCbv9ihgHAUsyZko8
ILWl+7vI8vTFNRV/PY28kTchmMxKs5tNfaPWf/3hawfiKQnO31TlaNQ/MTvmOlv5ucxYCavo8eo0
SrEcn/0lC/1yXipZOjO+0NlCXa4z8MQJc1iqvnhpzRHOX9PU8+Ifb9qtwFhIqg/Gi0k+P9NsWqln
i9UXgTAEH8GK7g87WSTB6FwfJfdNnlInuupbvGNmuwgYeRUWv9/UQmj8oRNgT8oC1gYclZCHdJCU
9CudsMy5ahvctv64T3eMAsbfggXoHCKmtdsP5E+jhhZZRqTAFca8JfmhtsLJIJYwL/OVwLRaGZrK
Nkp4WbD0e4KJptsaC04BUhhSSwHNJNcWO8BOckAIi9OY+tHjrG2YWfxGSzWiXP003kDQK1lukTHj
emch5+rg8x1+dnNSc3KYa4/Lz29h35Qf2vbijjnHSvrLxXgsMWjORfIS+i0hmZEn8jAdvyioqx3p
lLxU6T7ikDO8NwdHBXAPgjygOI4zZvTUecEhiSh3A2I5M6ixWsTgd36oU2EyoZOh5fkPbwly0DS3
qcrtJZi2TWkc79dyigZ8DMKeJE8QkPqDAapGuyHTEAsy4OsAgKcjXrwgEqumhs5JucHcfDe6JPKc
NP/UvLeT4NEKPd35PUwlxJ+p0f+dzI+z1EO8PNQo4aiqDsGzh56cYEK2JJmQhDzuEG0Xk3hVy5X+
Lp8nfKbjbRzR9Ob5lDz/RfuKD8DJQNgnFIwA7O156f75PVUVGCDbk5PArsHLNMb5ruI+pJeVYa/H
fMfDZHZvOvvqR8zXfdQpvO8kFC5CyHsfHgBuFyRZFOPXIdNffgZC1ezsZsbl1Ss4mQjgV03G20N8
HsK+zAeaAv6YmuwC/uyx4o02c4hJhLvajNde/AOlX2JFfW//PgAwPP53nQSyy0+phPKbAKivskTt
AWc8DTwbMMUPjQWmvhitIRXhYokrYobdcgsDHIg2Vvzh7HSz0HkQ9NQKsoAYUwUnPePdvyVUlf7I
ZdedxtlUShIaeQsH3jmk4B4A+LtK7QqTwc+zoF8qLhpgiioDBwe3MTVPHPNTb7RZUge05pdzdBcn
LTYv6OBySH6mojs6XpZuYSUniuaYp75FebWtjscfTX+wh2ooQs/TVRGunMLcBijZRpgXSZPOgh0X
lCyjpFhseTIvP81dERqekUfD5J8+i0OCIwdmehOwNbjgdcn7DhR6U4ehFHGBEk0+PUyQyuzrQQrU
2OO+EUHs5Z0MynVy8VLci515hPQ8N41YCGB7BBC6EcGlRZW6YMCxGHXaC8LFe37XH3e4Y6NzDH9m
lPexXxFtDXlxUV+uLL1Wrg+l/2Zx7O/uBKcuDEGgVIbriDcKoa2xO/tItBsIiQlMMk8N5Z2U4S21
//1l5UsLDpS8yHLGOFJKJUOkg3UmeQa0N30oqScneSNd1pVAL9P6eOFBJK+1cMZufnle8zBc9ka4
vOGkxshOp6li8rnjs4+KpaW7a1LW9YIoiNPFAfYc4Atp2Ul3o8ZLAiLkpi9l1Mb3UJDAHZUH+3qK
KO2jEufr+FEwBW2IygrnObSNCNtXZrGQ6Gt02SM3D7QebyvrZ6KI+ftxYC4XlNfC9XxLC7Fg8mGy
0537Nv5R1R++cWBUPK1sHIF7aGCF/BPhrNrAwoSTfGXLhSDhGfWoMuh8NslWWPNJlO4+myB6QGx9
gwk6/L8EjXtneDwLhvx/Zq4NP+GjPkZG4HMCfDdNqx/gOgFbfeREF3pNmNow2jD/XEKJRO7598Aq
zAkcMv0Ghej1Yk4MdBLY3Q3h8wmJTDtFcLUqesMLKooNKGMZKd/VwBLUJZy/pZ2dEoKwCVFc50xe
b0D10iaZPxCKlVqe52yWSEnVn2aXHwpnOyW8sGXczb5f460pyE5YoOeTLI/OMrJHwqPd4kVcr96S
LkLBgIu+IOX94Vs076NwF7zTR+zMqN7tPpyGB5epev+Fj3dsREyaGTNstM+nqfOHDRflnBbWj8i+
W8lk8OqHddT/hJ/mWBfVtEkvEIDV6Lh1vuJdQxCFnjp7c/TbSBuos47i3uzHfdVlGyWS2pyQq/gg
P8f6h8IbNv/MNTmUSZY/oA8KtNKLZBOud0nz6l9Aue9LAXRRuY0A+jKEuxWgF6yD56IdhcRnRrFO
mm5poFtp0Ydh+LT+0QjB3aa6SmC4sNWWsmcnQbcNq9uPRpt4eWY9SI1FXxxmcaZTAecK14l2ZY/Y
Z3ue6SKcd/Whd0SiDUtoyOmNQgVU52SBoVrIEpEsFMRgGWo9wWEXo09OJnUb/LAKFQxeCVCZjX/h
0tSmGYWcpP8PQ0P4o+A1+zYt93pImCETMARyR0A6dXx7tvTIKQlAzKEQk4tCu4WAvR5b8E3oXBCb
tc4mDGix7gvMmwCbhjc0CxP0U1eYBemNP2xhEgS0Z3w/qCDhujjYiP6K08Swhv39+QNrEfRsDRU4
nT2xSfh/4asvAJlsg3Efdnz7hWbznXp04emqmXYd8SBAWH8md24P4F/CSQBDyOSbDMH+GhVXdOsC
wsoa8phZ3R+VHdi2OSJ58iPwbGEPDunW+tbpAEE+XdgBfLKgYbWQ2loNkjqHPmfdrwh3/rss+azR
CbTaN0warPW35t8KuEGp+xz2+tjZlP64ZUq0/hJ+0bNyt+ZGsNO4NUdOND1eMBwPFQEhOjFmhjEx
k7cAxJK4w5u+ieSECLkI+NkZTZpA0s/aK2ZJFEF1+yE0dhZh8slLQ6DBRM1TQbh35I399480QbK/
jgj1OLrFPZUtJF3ibWOVFAehEblp9pXdMJCV6pmSQySXEGHJ7JjOQiL+zAHCOPcvYyRzUFiXS4ST
y0qiZh75XVeDrQNwzirk93Mzziu3sR1hgeWfZFwcKXSokOQzpbbwDhzYPLDxqKRsFjshbxlZn0Uj
4qHkNzfbNusFERAjyx67NWyS/WKjJHTecssr/jTmKylhBB6UDjns2YGuPu0TARTupSGDY/RFgpi2
9fRPXaVuFY2mktiLliqEu0dbMSa4vP8zyBSLOboqhOIfWKt6yO59RxZeHk2Wm+4zORCk8jHXn1VO
miexjpAuiZcBFwy0i2/nARSF83a8dBwAAr6K/e/8x+/yeIQjPTBBR2aWbqV120rqTwpg6apqWocc
itwZiWUyjx67BroTQ96nE7dJNvEC0vFNZTMelivQcRWMueGRLgqGiuCfPNGtN3XhF0pduhodHhq7
kuUi2zGuRt4FC8VTA8d4iynMIKxMsMElkOUuF100uUu0jZHi6O1e8NAbSSnNWMc1N6Nc9pg3nzTm
pi3U24RKPzosuObxrFVVxQ9l/ZDYoh41NCaRAeLH0JrifqrBSO313ERV7crXwy/fBZOdLcuGuZFA
pE2c4K+EV9wxDwcWBs3aTqXiQMZv6zwz7R8ZD17a76mbr9kbglRWCeSYw1Cy3YeAHtWoj27hGVq3
ePfuOC9gvS78K0rKQvn5aRurWblCcn32l3bRGKZ6fvO8H29XeKeRXGZaK6dy5atvszIaolkeF0sQ
BnD22i8/rPGE9ptf4f5mvQriWv2NUC7oidPyGjNp4G23EWyerCg/PckLKRvnTbJzPkUBsAJ0bokM
fuFWO3oZ2GNpfYPGiDJAZ1WaqjhhyPwgvKKpFw==
`pragma protect end_protected
