`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 59072)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpIZbHn7PpHRhDrC6FSsS3iOStQ7Tn0Igm6lzfB2j1izK1cBPjM4rTA4Np
gE2tgChiDq36yjdtyVtcQa4ctPVdMW3QmO+LYDWY6ee2FukqNMZFgUqodsUeWn4lfZVj3aUAyKgu
g7FRn9NMjgyCprBtHoEH8vxDSbRBgwQSRVw7/Tse/7hgIxxKpRCZ5zW6IODjnJhEFCPmb4Qnpfh+
E8VyP6LP1ACz2ZkcatQg4GHOr4VqZOI46s23/NOtmdFdAwcuOUyBLfaBuCwbefgGeBGVRACbEU6a
OkptYwyBwcS8lOtZGMxk3vN8L7IQy+OLfBVf8qZpyEPcyD8WKyuSIAdMrFSM+3MLEPmShhn17zJA
4i2OwUtJE5Q6SgIRaJcp8bxQ8SA4OJU+AG4PqVrWoNmITyLJRaO/Z4zBgti8k6boVVaqIKTbIjr9
SpTBWFVq+4K4xk9XwRBXNRwnm86MOqx3g5LMePHzBxpCRxSDcxv1/8EEI+bdPjU272+KjpE6B/Np
RLRr7sESCPCKbj//5nZfkkFxsdKjKTqg1xUxBpui6k2khi1io0uUL/ugAZqjf+pawImGUSIGyB1/
KMGgkMZNuD4Ywga9CnI+tH02sT8K2w4yzZSoPf2cB8qLdaHW54SCT/+0vDbIlzdnVMt0fOQF27WU
Py/8Sk5vFfVWzQYPzT1rWn6ryQz6LJigfboClzwju63LHxpxf9Rb88P5vlmCDM1896H22WbxeQ06
CRhDyXZ/OrNIyBIHqCT9jCFwjyJknSwJ6/frC9AC/Dm5i7fSKfdMTIphKsiI6Hs5KVlBXcmFZ0yI
RhT+ibFtAlCMuAMwtqwVsEVx3tTsChI6cI360ucb0KIj1td0X6jSZC+4zNAbWPUV6mMPt082dgFD
/O4ApbjtbnvOYrdrET3Kd9z7AiTkr5OyO6C5mYL+Lq/z2y2pRLUWsVp8jNzjmTMEW2CPmzXRXa/Y
9YWGyRTT3yEUnb1k0wOKFJsSqIHZXUOllW4m6rFEM6I6x8S6amGT1JJKP6CZpwBne4KXTyP54V/1
J7paKmTwOJtBOMOytZRajgGlhdjZqSaqrEs7owTcZVU5clAxMmZV/xTGWUYcGCARbL8KuBH7KTwF
lXPQMS87GJgtbMveDFuZphPiR7qfFGRC9EkyWmyLGmJajJua9sXPdYOiL9+uGj6l+NCV94nCgvSY
4/6YpkP5n/tWNxtfryuwzIQKAsmRd76foenvhsaD3nToR7ZiYUOR9+nP6SLEOSs+MbVRie/BEZxR
q25Zme0/UBYdlICz+lGGQlPw+jog+zHl13hE69t+JZdvLenZE+mzi8MEF48sVvHFWC6pZhQhmAPk
iz6MgmAVxaVJJdy4fqGiYbtXuZDwu5+VRQL2JUg6G/vSqBL1nuI1d930/1TqNPiy5sdkzXpFgmb4
9P+2+E/0C0hzCJrinr+cPP5DYdNndM02wMTILeNfuDOyLcX8wecwhxbPnmDWPdoXwj243tNuqPcw
7YBWTBvCIr2aM4vaoNj1uE1xHxK/DZq4FwSPx1zLPLtfezBNNJAT61DuArdFDdJxVKBc3gGJoTUw
HTJkKiDrkuoY07A8Xz1opYbnM3dBnw94wYOLjOvssWeAEwlshY58tOufRglwzYhf60aFdCais8Lh
+Vnw8a51UeenPPH+2d6LIuwCVh5G4rDOgn6OUOObIY27Pfvh8VBfJPkiW3UR8t5MRFSy9vW5g5gL
hn/5K4LcRL0uto+9Ohiaaj6gb+0Z92leESNDcm+lFdvwxZG6+rhnL8uacKj7LXhpj/S9/ewA98hx
sD+YLqltsppjJQB8Nc902kzoJJts+ag2Xe9ZGkfLg4+SHnX6yn/9axdTSY8basU098Xr9ioeJE+0
AHYkiQQcw3IIx6kHj8ulvPnu41hcGxs23TFW3i3BnFMzon729qad5iW0xbRBV7pJ/x739zpHogYK
5bSHpnc5N4eYdy1YH/rRu2cwc86OTx6Lt7W2wCXemEWgnV2jy1FqNg6ciNPIp8bUC2aKK0t78s8n
4lh9SVTsRpeuiBGDhBIqYXvowQMRXFh/qHt3bmt+XNDPMyFjsYZ+Pa9ZcbfvxSmSU/+c/BtxIwsP
Mlu+Wr1HLUuQP32RZgypvRO4LuwVjXLqMnZhUYepPFK6hHzlY5HonIDnH25Cx8IXeEQ3adZXpuOG
CR8u8hwTWstBMVD6JQvj3KJ84sDDncCIMQ02qs+SS9qsFNcdNTj7HPaQNpDL51HoJ/CgbQG6lio2
D/LN8JBXdZVVFPUCNA32t6eK/ZEw1hqOpQH/bG7njaR6ys07u7vAWOwSTkykkUia70PkN8eGTRNn
bHIdmu5b9pnonMZK+JoVLmGQGw2nRJKSwNN6MWTl3zDPQNABDp24cVYhXw9pZlqtGWS62/x86nFU
buO50Ew1mDxZYdkf5kmZJ0IY30CGGYnaV4YN7EBMfD88e1X5kELCzBi1LEvTdyrk17cY84+71f0s
4I8bgWH/FCBMwe7N+CmqgUVPrGOvuKGik2Bj5HTcqjppnirCSBIsamP5dq2jytxC5+X0UiGDCuVe
porWKL7bMtH3Jr45vzbjDN0jAQB54IAe6bPQrSFU9jLc7OvIPfpRK6MiaQDMS9LfBkszazpZKOOS
a31RqydTrupO6npSOuxlNE065GOWUZcwG26VZbkT14XvKhKJfZ9KYVudig3MIsYj8uJOOeh0JcQb
BBjvDn9Y3UmqS1p8hh6d5HT4stH7HSYJz4jQYTAHBAAg7SJY27xifr2UjnUMOOVr+APH4dGHpD0c
MLZNwvjrEkxhhZKwlWtLHU95N7C2ex/tuFil8MXYnJGUm6o0RIxtjhKOEmwhP7sd2QkjuFdWsSzT
61gwHoG7YhHHL0X7+2JTc1za8DLJSIVaypb6FJEHkxrlicSnc7jAmG2KDxnt74kBY0leY76N6BiM
zVtjcaK9ttl7NFper7gozziowZyyHQxDUZQeEc1/Ix666FBcZ7bwLt/rS7vc4oIKdiamVAexCHjU
XLWDaV9WZGQPENmWFx0pyIeowH3IZ0/1v51c9xltfunznR8b2hud30xShgftf74kk1z1+yNTDMLd
E1NQikI5AY1YryCNlD8hmHCCvt4oboE/rTPrbgJgx2uHqSqyJTBZzDHPkXKMdvOZz6Vyc9zliDua
zDlKQ4Jq9D+Jzzu9WIHMFjguwfdxNt42OHABuxBqVBiC8fM8MfJTY5mor5rNm/cHFvRgaXVGzfpE
et0acrhD2dL/UKjxgikZNdbp+ZMxsKmjXCFXjma/MpX27+C/5U/nP2ZyrqrTNhGC6ox1iMJqsK97
0ZNDgT6kQf5peQheClZ9aNDLAwCLcV4ngWzXAp7CJOxtb8nNN0hNWEPXlWI18H4u5xQAvRfnzVNC
J23DDHeKAXQ+o6GgyHhyGoTwNb0SGIXkO5U1ic/pMuQySGrDyO3Od58xG6my/X28oEy66xKmezaK
Xp78P7xqC7aI7W0sdB+dnmIx8kGL4K5h+S832O/O/AvYnEuxXkCWesBvkSUeOSnGoz9D/sFFpJnH
pkJnree1a3VioA54Ctmh47m88iyuaFaUEQHfa7eITNR7MwFZeZxirfum9mls87I0nQaYR3mEfwrs
XXeUSMCjPMGuHKBsqJd/j1XOrepkc73pvztHUSnVFFgBLwKSrl/53oesWbn6OBCu5H3JcAKO5Tdl
wOouxeSXEXXbKzA4+4Hs6SM/ThA3/dQo4LEydWMPfJvMsxb+RVH8QS0DLKido0tFpmc42KRR/RAq
sMDr7qeA8KL1Cz3KQOGq2BmCYIa1eqJnK7jmkemIhB/rVO4ZKtJecMGRYDKx6s8w+PEqqrkp2EzZ
6l/kA+KCjBn8xBWCBPzdm2EhUP4bXigbmMOYk4cflIgADnynWiiBOablEnjlisuaVSxEsregUCdd
6Gq3OnW998ZVTHFdpiY+miH3HIH8IIQlYM9y4noJ8YAo+m0UMp2dAyMzpF1zTtbEabcDGKtNgjkh
g6byxZ4oltG54cUNE9Fb4yROaKHtbmtQnm9UfEAzkfTtJ3W/rz8XMedg+0BJ2KsvVPb0PDrCbmuB
YbkA7nqSJYsfyuC4xbfi2hihxUNltkMl/pB3EnL/QZpQvTHfH2uBwWMJLRHah/5PNLC327Y+fXZJ
8F86WClzUXCThVq+XO/x7a3PhaMx7UsPnedT5YtzC2qYFrUUhH5jQQyA26a2SSDSNseTsRENLmLs
XJSQfM6tJoGVbzFy+ktirfiYiS/eAId+aZzxEL5uCH9o7G3ecoEmQ1HdSdHdFfc3Zp//NwZC8IVB
wOGUb88HKSVCtI39JAwKRAqG0S1orBtkGdEiblaVVMVaCoIEbcUsC7igZrCDtEooJ136Xri7DjtQ
vmQLtPluohMWBi4jpK458nIiFj6MI4mDKzswPgikBwNYQLfGwDEjol4hA7qePOp6wlhvFzdROWsn
vDUOjrwxaiWU+Cq9l1wHHn+OH6nN8uCfPnv2lacfzozwTy+7Mbdxq8ZQbIzrT/y9SrVEzqrc7/ZM
AOEoruuD5eMrFKLcDBdvlqcnuB1JBZvXpB3fm5DLxlG7K3n2hms4ziVn4FQJ0ej9htZw+5fFD2T+
sqmg3NLiG1EZCUexlFNKSBKt+nCbVMeR3osR3z1e2ZeQ7WwgVRnqGbIHImf3sR4p2yIMdek7Xcww
WmTONe+9XTMDWNV8CNY0Y25qjXXyfnUDLq18NjUZdSGywMD20CKYhrYyQLvNnPZwiVgPe4i73j+D
mk/QSDmQvq6UaVZa90W+zIIDuk9VsYUME8QNABcNLdlrnalsYck8S1KixA/gnSuGHOyXgZA3HghQ
1AFpOCW+P7MZbzGD/4FFng95fomOhVAkiTLyy1SKvKY03lAguWaMgAbfTLqYBLo0KRjR4lbIst3x
FNCxKosLSASPtV+fQaujHQiH7YAiYba1QuLYk6lcvFcxPKlWOU/C7xmlIhDJvP0SKaBPCG7Y49x1
ebaiqOO23SQAVNAqteL8qsYJNuZvCUsFQFi4oo5X7xReY16K9fpoAS12WPzK0Vsu+t1sSbg6v5+u
DUBZJ3flJTQgDCkOcUSDBv+vjUY3igIgZv3gJ5pPaCPXQEcB12ShNPSgDteXrWqdAT+lowZZyUVk
xV79nNTFkDsXGDUzgb3rlEj4usbW4qJT7Mf2p5eimIZdIIFOx9YiykTCDuUAlUYsKJKdwqpkvnw1
hYpxpin7YWMFGtf3mfy/EH73hN5Zh3m/Fc91qE68Ph/dR4zsMF4bTmkPJIC+iOSeWjl4PbgUX2WY
YvPObD0KipedeaJEdTX24HxTLa2bxPJUTwlZf2LCVTfVP1I2tEAsdgxVw85iYsiOs6niXOAPjo6u
h+ebXOQxlhoS9HEqMtXZAdJhb7FZPh760k15IOv4BHGZZpLT8wcJd/rvNi3O8X3mauoYs7p8mG+S
+PdRnVfmcNrCn98gZD+LFgWUMwKVSxSyoZlpUzMTWaz594kUTPRa9ci6UMG9oN/ZY3EGlCTFYLC7
dpchtddYpg7TTb5LuDCWhZ7glj1bjKTX30s1r4nJUeY6RdfoViN9G+pOpdFRlexiAJmMDp8Dz0Z3
oC4SBqd0RkZ9qgqinsmDGVa7qxQ6X24PdeKqVrr06CQS+tGN4oDBtkJFaDF4v0hA9M8yUnxoCiSf
lTiEdl3DT9QyyxCzF7V+qQrU8+rc+jK20rtevI2ortAqPJ1kaxiRsyuiT/BXC2QYI31tKsnB7VxT
TqLoyXSU5ilRdxZd2sRULNSNO3MNGlNoFSj1k7R+zJIIYwDg388nCdaf/xmQ/Nzk+eEJ8gRfYIoQ
3ngT+V+O8F1WbqdXJFUhY1u6OxXoFaRpF56bGfmgunCNjOIP9tv2SDdoMjJN6iyKr3JmDsFnSrI6
7s8r09ML4Mptvl8LsrxHKsENzcHoq96izZrMSDndNFJGpcy2/p+lUIQdMCAAH1aXJWcOYMsx9C5b
8o3ia/zI+h9tIQr9NoUtyUDOSoCCywmObzBUdwd9fHR4inmf0EDLBdhKHhfM/usYhDtkxliG58Az
qs1mlt0sTn5vc4OAxGeNhK1WVJy8HE4ED5GxF/t8cIypmqZOEQcohPY2iiDL0lRGCqc5KK3V46Kz
HWIxFwRjLaoH4tZY3pUm3owEiw2i8tCqvutlOnp10aeQ9qMZLwvM9fkNbvCMVzKFCiEDHJE+B56z
MxajKX7D9u/DThhCL0NY1aMDTkssjdRinT1ffGUtRF37D9yH2nW5xoelz2qsUXnxNVHh01E7sACc
qWXuplI4TxiqEpo+gN7jw05v4i84dzsKPtq/fCbusrhxZsDH5AmRxKaa1s6ai1uXvpZpFJx9aNsa
uGNrsd3C/CZWsXm0IW+fIkS9hOYd4vKUZIlPViK5aocb0Muf8vAkKFw/yUctp3ihcCxfZxyObHqc
ClU+SvlKFe+c3qW6wnRas3BrOCRx/dIIETXYDDGCSyhDSn/vsK1UWQ3Y0uQkpB2fvjBDq51BREyD
AhZAWXz/hovYH7rrnbRKdJ88ezXruZQ1jJuPNJx/lTyDy1/ZLCAoQZPzDg7yGbi1ktKybLHB7+um
vxnBEJBdIRdGP+m4yo47duCjmv35Iz7ZWYLB8BZ3PfpHPvzu2eTv9C5UYbryUGuARZsgv25BTReT
8d8f8M3cTr8TbMq82p1M4QiLfg3SL+fueySfw7iIVyCsHX0crjRdO9vcPiJft4RprJ1CNcr2L1LR
rV+j4cL1E9XFQXtz2uiM0MfrRkxp7NhXWfQrPbCcyuM36oJpMN4I1jz7I3QeGJ8g7stRATfXGgAT
nS8VcMyamkXM2uEZJ6V1FkO8GKy29NnU+el31LUjmuGATMPh1+3Et68VLi9jtivEsJKfhcVOULwh
pLa7AyXdrsxEgcIP/YouAeLziE6sAwMI2bezLakyzZHDKerK1PYBxRvrhqtJH2LbXCM4H7tbS8KC
rKI9DslvtT7G6kEhxYbCJLHTMnsjvAyKE6dOf2jo2Lvuv6kcjI+JaaShzW5hdZzWOQlkupcEGItf
IjQft+2QnEXf+jAt9pWQL70x6z762xLeDKBI31bg4K0omCerTrPEkdn7UaasG8exj2HzCxJUwh4c
esYb1B/5R7LhsGc4Tou7cbMzWcGWhweFex6fADcqpgDLMUIIgYrLDTg6tNc3R0trV+P+3mCa70vc
1KmLGP3c+WoJbmE87klCcjAQUFTKZreipobs07uJm/SGKoaqEKHjGUW2acWtJxDlylUv15+aNelB
SwJnyCaO0fldqyF5s/Ww2zaVs48OLn6VUlyojxwHND+YDmQPK0tr1kxnhHeef1SJ7R8lekpSNexJ
DbI/uyu71QD85s2aJFFuHP5pfB+P68INEoJT5MvxXYW7UYCBjk5hntQFKrmedc/W466RlhTe4ure
ctZe5wkrKwnRY/kYhmpomzasGMbTy+WJ3dWal2zorKPHi7jajFlBhEythoBNuBwGJMjECt1yVBKn
B9SxbrklAQ9xDvFX2Pk6+tK7dypFV1ez7d+FniUeH+9cwbcrEsm7CbKTdzYRFzg6O39xWa8bKdXR
hTpQJIdd9pSXmpOKAJgjCjuz4QDQ7XbPZfIn7078uZDDMBXvgkMo5+iyaxw/J5iz2yFvAh2kq7em
se4poTGE66NgwejmEP12u+ds8bYuuGpAIC2Y+hTkrffhA1/T45OqIBREXRRG/0CWgv3qRNiDF8vb
M8RbSg4pjOf5wHZhvxxNPmC47wbTWv/7jNtGqveMJ4D5h4ZQFMqVRqpqh97ocwiJj94OfWY15cwp
RvdbEESpt87qHB9UuI5lLHiPMA7/cO70O89xTPqqUVOoO+9jrIAhUhFsYmWWHNBtcFYXVc8o6a7v
nNim3wgOpyEQk5gEnLJ8RV4kuxJL18HIK8VWOpMgf/18fogThVg3Vznxg0jfyC/9yDnwjDB5EIvo
56Etjs5vN8OZEptkAEAVAWBE7BRvAZbpDlRURFTVcAa9p9ALUd1KnDkMtVdMBGW5TUH1ukKTAwwt
Kead8+fWLh/wcyATV8n2kcbVZ1AuN0OiuAUeuxpxVM5CJnA1lK6k55XUgqn+evfMTRquqhOXU/+0
IM4GhtprWnykst7gq+f4FrjlIivbuukXYS4G9d3jUd+epYQ8J8YedrcfbLC7GGFTUw+PMDHiyXj6
brhXfZeBQWuAGXvAl+EkjzpzpxxsUU1CCyzVhkwm/0SgdgpTa22zZKmcll7cCDFXP4+Mgyxpbkej
XjuGqUEG4SAzLrA0sOmfyrnypdqT+ypaJn1Dq5W0FZxMwxFgaUwytr/Qo0lHj59nUD9IKkqCQ/ep
N7LNW4BJ/CXTeHSjh2v4PNjNmI82B6mVVUDNIyBdTKxiLGm82wqxLFkq5MRsFF6RxgnKhOLZUxab
/pmY/4pUPUAvmUykxYOskxV0vwDy92zvHUz5SHz7NDQ4oqTBmZAMuMuzNk7J8az7ksjB8Lxz/mF1
KMfurfrqQhA2RWkJkHSlVj5zNIBmICysFtg1FUQ0wDyAL2E0sp9Wjo9eV4iNOEZ0N1ZZjL/bGyQQ
sjWqMEgH7pLjleWtGtvY8oUoc26VLZuOUuojUO45PfY8yjry0k9lKGyBd0I0dQFxx/yT8LiE3xI5
BLwKgJIwB7SLJGmLbLsUBg5puRnd6cGoaz9BkuCMZ/qP7Bk2L9AZqZRH0D5U4IWOLxuC59aTG+I5
8IAvMUiwk0J50qANt7zQO2JNbQs3JmF036tOnDuVQsq7o5FgQcWrnFP9Kts+lwefHAp78pBnR3bP
UzFhrTyOyt1c3yJ6QNBgD1GlOBGe2A1+460cH0jOPpNpOs1EtR1kbkOmJO+0XDkvQszTflHxUrhK
s2v61rIyEX4BIFAQUEhpHfV4J4jJAY3dYfPKoDs6yfIwHFcsFSARzCcRHekXUUQEqOSyHdNnXnOt
ruoT0vaMkaDB90zlU2gRZsyiQyGRUjakKoa+nZgBcNqZJiLXBefxkpom5Z7Kl9J54GeDD98dEkGv
+Y0WMiuQ7dxW8H2HdmtDPD3CMck7Md41j6V/N81mBRYlszD2WaD/dEbRdht/DAVLKprpBfeTgy8Y
nd6taCmgvgkjmf4lIQxrgOT4PHCwZpSe6Q7BE8jHSTFHQY1e92nfHzmxybgDgvHxTVY+dV5h3VTD
hgV1iwg2SmRv6rEHiPfM4J0dp1X+nL8MnKAAi/mK2Slgp9ban3HwahKoNMIWu9qmPWhv6lxfmDmB
dReahcWIxF5quTgeJIgt1pLvUKOQgsOgw22vJ2uN+TBYQUo3mM/T24ippZFfZ5tQOxz1WAK+0E7G
3OvBpSt+jFcOd4SGSw5PQHOtsPvor8reKVNfzDDHKYiRQmD4Fv3mlpYb1QT5ztz0RDxWKk4fACb0
c0ElF3MTRFt6hhhnhmkTpp06XBs4WvwzaAGwBP9V+Ly8U1QX2jFV4Cy0RevGYOghVxriW7macUN+
xgTAr8oHjj0hewvRcecxIh97oMxQa+BKuf3cYcNde6Bhvnn909NbB1k3yP/WquxXGcX4+JCG4nV0
P/7loJeHzE2KmRSIp+nEhsumNOJPDmlSEom8F+EhvtGwF7uwPOp9mD6H/tI465uo+YH0sPb8QccL
/8KO78GKEdsFFQsPurbS8ZaEUNLtZ8Dob7H129K7ph5f4QjxNjvq4iLtFzizXGiPFNq2XrAZv+jm
tD0RX5vEQa8Meh2moTzKAvXpBUlcu2HjUw85gWmw5DDjl3eP7kaiuYhv4cx+0HeWM9w89wz5fzpr
QNytK8aKOc08MyCYrvUHpwzqbe47dF4wSB2ztKvBY1w05kkI8B1PilVSbLpo1zrIBU6HJ5TWkHaz
m9turm/K8/ESub7cnUN/t70tqE11WTVd075Uc5LarxIulfc/lDnqvspnQa4muXwVJ7KDViPvPj2u
ODWEyVfGyqe7RSqnKSa8IWM/2fclN4eTrrLhsNyB+zvfCGmx2/LsAenbX65zAhlp5+Hft1vRshdg
xRRvzwJfnrTfitaV3iQ0g3EnOraHRVPPrnUzsTHXujSdJ5IK9vUK0othQdaSFOt4Lsiigy5zZaK+
UU7zXtNCh4hp2V4zqnYS2xol8X5D5hutx3uISfZ4fTypWqWm1qxbYH7iIafuc63CtNpnXedxQUDy
JnZrDbxSLa2PW5UAMTH6wgqFw3HiilPA0o2D+Ase03cVHbSnWmFI4FSXTlLaPcvPb0NmDZSgbddt
2VVeZ7d6Uyaxwz86eFiOgxN7TCWBHpjKSGDzTKlwP8G8UsmvY8Sl3goAWrFNvbVOiTSICPhHc3lr
b0mq+9jZ/tbq73Lz93ch4foKs4p601MYsf59ZBOeXQvuYTRUi5gyKX5VeMK4XSepogMQ5DkoCwq6
amU50IivhntsfFljOXLS2uiChd5DJxfnboTLFdIOQJaFg9kyjpUk14FBKsdtDIAfWPegNhsk0wvY
vu+IdgsRBiKOXmD7z3g1QQ/dvZZeP1meyWAEj/67BYmrmdkM2Gd9OWkoG2wUoQSbjKCAAldqO1pM
RJelJaFJWNIPvSp7CNXdaj0Nwnnkz/5iDaA7+S15zy2DUKge4k8eeoTn4eOUmZZtWfWg3bBltcaP
DcBLGnLqwThiQalITBd8WfxOEkZ3IMDRdHw7DaYfG3VvxxRhScowr2nC0AEtHibYH2RdShU83WcD
lyqCGWlSIAOrXUuWHzylCMv9oCx8YSdh8cLj3/+9mXL2b3StgfxVb+6hcZ3tquirwTvbECwNmY7l
9qRQWoxADknCQbtn/VV0UTs18+OXGE8mxJQwXApgLFZeZIDmqVHcVYIVqSKBmhK/lHxBSX/O3IHs
G26cKGQRkvwLUcZsZ2npwLD7TGBLJelNoCS5R6WfdVePFfTlvAuVxj2d3NJXtV6C6bf7mgZnojEs
C0DgH8ozSwxc85x0bJur27wEnsZJedzOhawvohMtITDt+C4gta/3OzHGPCHrUxnGYApspGdO1mD0
Z2rFmI0TyXF4xBVHsocZe5lKU2YNnJF4Ob4oi592pjccwGF/Oe0ve2TWyAvkTGQgGrHxwPDGJlrX
wzovsikQs48j/0dYaA9B5UJTEV8YuNydasg+1WyAbRLXKLEf7G6pJEekZ0rUFDUs61g/jT/164Zf
aNvm6zRdu4YP0zVW32nX+VEoIP1Y1yaAVX+V697Zfp3tSUTteto4vr40w1TKfwFps6v6P2DspM8Q
JILjZ0WqilTFlGOj8eOt5GxUDTEhMPFO9K8IC1kA/In2Lbw2CdfX2nqbNLBdkqjY4bn0bgr1tmoL
+wnIR/AROI7YZuM+AMv/NykgtdaXi79zpyZ38p6cZWKzcH6UsHnCZxCxowpTvqNR54WF9dIA/wJc
WQZB2Cna84vKenwRFKF4PWh0bufaXV+3DhLsTbKxF0MtYfzmZKi0knQBzHoS2lpFfHtQ8TcWPGA+
Q8+wDnLLT0cmI5WRuLI50dZim73biIFntr+NpAo32FUSnP0RwE7TGHJoNctzz+//LvkYWGqN5pyS
zhT1efQbJ2/zneV7CywywTgVHlE6ltJ9/215h0MUDFw0H9546t6PTTpNtSBT+r4fu2VJLqiKv5J/
sTGCV0s/RW+JtUpFqkDneuHeRW03VV1a544FICOTRShFA7xuUjdQPHItrzUQreaesXQ4PSdPgrqu
VcGp6qDwM480GXdZtLEcjCyA5StQ9RmDGTQO4dFnjayI1rnVC7JKRmokbee8CWzDYOm2TyCfaLjK
f7nqOhWFEpJFOdoIRv8M9LQGezYCAWyIjCr0s0K2ql/2P3LgISSScJdIP5+eiMluSsrdbOvCmeeI
MgPDNxK1NpK8ovfVtushnox6jdUo0R2kAHt4VD/mzZmuHuz5GR1uG7YsuB2M0oyDAanr2X1alLQ0
bw9l7cL90nJr4z0aQubRU+a0DiKZgThZLoJNR2WOrFMqE93NX8xjmNAmRUWgKTLS/iyXVYXM8Ri3
U+XrhgeoUWcXC86uJdG+ZtgidgwrG2/JNTXxqlUbe02yDq+BIeYYp2PCBqIwP2KAc79+X7M88oKY
Ecb5eh6WO0SjwmTXplF8kYrELTQ8UfccpoYBrzotbRP9XvhixEX8Ey59YFoPGLjQrVgi7OEFumEL
Wh3NQjWviopfZAcVDcOGfvIBJHDfLoJtiQpr4iYyQIyvJyDyggL1vLNUS+gizCjA2tFbw6i0z/2q
Y//Q8GkReFJ34DG08+g70gzFNiNZ4Yxa3r/iqp7I7TocPHZmojSBIXZ940xSWKXOtD5lQANzHc8y
eNzJCCQ6tvZbUPHkK385/1boNFDLICGj0Sm8rdyirmoa89s7aQ6SclcdklbPnegNJad9IrwNUmzx
mqTQJTSVcqquqOd9aMUDfTWNgrdzNPmOhGdKyWMP4zn67HBEWjIlLpImUjaa0quct41q7g9AdMlT
2fM+a7BnMRMG9MifRMq02yp5K91uDFIuYeJEJqXGxlh2FNOWED63BKkesTWOc2Ck8mYt4+1SJQKe
XPP06e7ABq3VQT9m8qkw60c0IY85e616G8ph5iuHAIU/6Ctw/5s6aglGpyiIqpuT94H92Ch/B0mw
Nz9pbzyL7R+kEsqKX+fEuXzcOFjkhYTFbNtyuqnNPu8QHjzqy//hCCCpWZFT+ZQjZszTN95WCT7s
UsL+fwONn8ab1wsLATiA8g+nMBtZggyLweQCrERjT4alFXrEq+3q6JUcePdy8TKeDzIqyavSdida
2KmR8lAt6GQrpdr4IFZfW1o5jcFFbDniJ8cMB3M0RsYXFkGQj3/beKtaSY5M0sGAeIeW1hqgWS0x
vTKbf6eJaAd4ZK4ATM4C77+odIJg1H3M5wdP41K0xFXG7tyE1ghZTGvy0KoPJyG8r/ahBLKVYGoD
kIUd4w5X4gJNakkOKd40IhIzGtRaj1vqQKI5+n21Y/CGaSgClJfsWJFTUzGQJgTyepmYTqdFQSdH
82L/UXtPiprgj4V3V+ofQLqAjwn7/SzkgiAPxwGzLbTh0xLfx5k5jIggMOJdIWTQU/gMkYn9vL8F
H7sGrf8Q7knNxju4ONfkkDMPd3rshgdwyiCdFs05mY8XdXYYBf7IdAj8b6VPnf49gJUhCdTVz+wb
xx39eIvD9UIzFulgiIO9ToTl8DLttNmM/DG8uZxCg3C+cIQ43scHxkP9L23aNyDeXIFwdys24rxJ
AgMGc9PdoTMDqSYPKErkm7uHqrZOoA9Ztb3QdUpuZMraTecrp45R20xm9I1wHZwu4oZ2NNFgQKBB
LzjJZ48oaYmQMyfoHc6ZBxg5/f20czL7dfiNh/Gx6Pl47WtYPIE18pqyEvZ6LL/niMw/GoRebNW8
RLGW0BF0JaBrTTlc5bJvpO2NuS2fGemN4Se16bnhk5Fj5tEp6Ug8l1Cy5dNhstV2txMMVvBgHDFQ
rxvu13vRQ3L2nrgIAaiFP3Oa6fgDttZOOpFnjP/VMRyWtUr3PtJzlTXMZ5k38Le2P1NOzbpjUukl
IaS4XUNkfTU+HF3tVY+OWfcCEA+iwPf5mlOFoQIrAUMZtW9xEX8GGHXdGelH+wEuEUVTmvG/6Nof
Id9EywaAW/mr7pO+ohOEoJmDALa+zNSGMmMR+10fFasrRKClDYE3eTnhvhsaSJfQIoQS2mQKv05K
+bGoOYB9hWT5EqlDy8b1fs1TXcaCbEYU6HvRLfjrccgX8AnLn7wA+owZ2hXnNa207D74yGQQHip6
9ZPga6zA1DOElgfVt5PL///tvk++VUi0JaFfz8gw6IMYNl2lU49R2FQYqJGXj1IM4LkUXtOwXexZ
0JoXs+cgmFq/1cU5YqZMR5/IktBiekLgfZqdKkUbFURF6LOOu35+IYxBXRZn6muPMEMupUJdoVXM
805xoMU60NnTozQGMqIfYeg3JX4H/TbB3p3cV/17794Jw+ULq2BBx0P990Ii1jb/pBh+yL4oDKXd
OOp+KeB6bJ2R35utU7vFsi08MFWsKRusnSEiCYaZHXou4LaiOAGeTO2To6dv/nJaEx1y6vJh4Up/
2VlkcNUGIpDHLwgbCnFvuu0RZ89HOlo+wX3j/cN5HI3V6KjyOubgswgKNdNPCNCdqmV94LXW69bA
vtP2qtK7e9wBPZD1eGAoR5b1fNmc76FAhJ44WgZWOIgVsNZmhWusEbsol3F8Nr+4HPwCI9XHogeu
2a94e2dwrNKrchu3WvkXuW8/BLQaOVqPAWjrsKdQqRxoj/EPZXR8Zk3eK1jasIbx3vV181zwKUAg
ve2W2uWF3Ts3rGnD+1rxDHamtIck1Vd2fvcHPu7HiPDo0IcGBWoPylwgIayMnjUkaQyrG+D+TF1Z
Dzrao0DCNu9D5fZvdQ5ESjxT/6QvepyA/IvGrLvigxbrxH8/RcC7AvIoV+t+uCa0dP7bwV3MTesa
FByB29UO9Sr4XoRKZdV4SW6qSgsmZwnSSD+BTaEeIay+8LExPd9lZWjeSFwp9XkA+f70rvX9IFyc
VYHp2BbnwW1xo2i+LoeBtkLfawJvQ0iF/N1gOsrwHMMEIPEDsAuKEKFeaKsOySiq5Xr4g04vTyET
otHigZhcnNss+lZz+QcrJjhTg260fNgiOo3xNvA8TZd0xC7CK78qUvgGEY60Z72CTiW55ldWWOfY
EphzntmOuGLf+KRB1aptZS6PsZGlblJ8LwirmWZkTGWG1C20PxJ1bET2l1sThqz8SQnGXolV/CQ5
x3XsRuzO+wu9bNo+DnrbzTaOP4diPX4Y4RWUzR294OwozItfCjTjrZf49NtohcEaklg76LoE+LhZ
nN17Y9y1FCARrlsE0U41ZflQerJDSattn/Z+bo9voHSrwF2Yqi3vU3MAnrnhNV0+Fd7rWetRiwSK
GfX3O67X9edPMsvSbZM6fPbGq6c8GJde0CwPPhWkGvjCB2z+P99APAfRD8NFSL8QgxnoOdrHka6g
PIcRzSA2T2EJTAj97712AuezyVJHuXwVMy3oQ4w1rrigeurshnaqjvQ8rInGfxD2iqkxsHRwchum
+9nR87ygQNU8rh3diRP1muw2qDaNSbGJRpIbM/D81EYcMOyggL1bRJFbO3xRaol0qdiUk0tEHxbv
lHrE/CsSsSUnLMlbCuB1hMRLKnSBbiTT/5MDXosrkI37vUnnqKkp2JTNo/EtwiQryKZc8b+0TBcK
pBcE9OmdHl5RCNrermSuNmhihjXKz+N538+8fhnmN02/n9vX0f9G2A8m9Rpv6GAsyrkVDQrlkIK7
tbSGPYhxwexuKof3SGfaiWGxl1KJMussXQfSSJppgGztpjhwARGKLj9+Lv/1UPANlXpeVvpRT77s
N30AzXQR7ESpGGLttdKSDl2SGO0y4v4GbNN/gUdnho4sbgGjR5QRXHK38hMiJoRCJ0SWZW1btIWl
LNMrRkkvUNi1PZFBa1Q4Z4DdCTkD0HRiPnB3/8kJK+B0a5TtTc1Ra/geMJPUP/iCrJ5iE8kUATdv
ozt49xWpJ3xvJbW+AKTRGvD5yb1Etl+Neuf/YdwjORpWHll0H3FSFKEI9ZGcXcmxgHYDFv5fLAy4
u+LIlVb1pDQW6A37hL4rVZDeiHlZ2R6hfEZbjUYbwWmdadSBk56QLi+Pf41BxwYgO7pqbIhC88uN
0scFmKzhXeKL9Tgi/zew4SwJ5njHp+r/1kxu53VXQC/Aumgc6zyaoDW84I/2WSI1Oqd9jZxy3/iO
t8K53dLdHC5A2KymkF7l31/E2Zu1cIyetkGlzn/urU905HrwgZYd1fdqGQRuySep5sG0+mlbIS38
yYCnOGgsa1gdn6gpym0MZCL0BYRIbARNsy1x0ejiByUZzqiXQOizr0YyAPNBSmQjkiMoy5nmsv3g
Vby7MbwVjJ/w/q/GHIZL9RlKJTwwsrM2rLlCtd5dghb47Gti9lsuZkm2Ogu2ysPreiewoUgzAa6q
nK/rxxPNbwSgC1juMT62ZllRyXDIQYaJw+22BiNY9wR+tAfXgG67bjbAtlnVs707outYXqMqvjrS
0yHqbZOVT9pDWGNbmSoX95Hvw6dGotaj/Ow3yKP65/iJltJSy0BKBLrsxtdpkLbj8MqC5bD+ydRO
DjFfy5gxmotMVGORTSDwKuFIhONW1SgPoTCu9RcKiZuue9ndX0Jx2V7hhtRoPeCpxGZnymXPTdy8
zw0bB0GgqotvlsunU3qDkQw/N4nDCehv60vck6zG551D3H+7yFXeWX+ESHpMDlwoW7ujG9XNcLgm
wwnc+7zbC9pDzK4OVtJsZqrHQxn/3kOrtaC+DRntWjpMGiX7BBw4IPSn4PX2Mo46IxRyLdd+Ek9I
gGhlt/cJw9HqSvpBHdxsZgh8/xuPtBZ9AlkquwCgPOcTF8gp8pEjaZbEFA9z8wWRFYlbmD5np/Lh
Gm3f4kjgvlCkfD5T76Hvq+T7htd8iS8dcq51tswQucDdx2AY+btVbsLbaRGfjeYNKaf3YIQpJ0Mg
tsQ/8bnUuYX4BsHyThOSOOEIe8wLLeRtIPQc1UTICUnw8PB30tWMJnODlu4yUtO9slOQB3gn5m1z
QBhJ+696upoGKIGhLnIVZsEiAGJTwCx1/ScxjM4se1iHmt6a1DAIhY5p8oQilTswK73d71xtpWcO
P4oTphhqGVtTLw0wddIlqCOKsxRdZJq8udv7uRb0pc/ZvOMywB6jMr/SXHWSJQ46SQ03RK2k6sqe
e6gRUJFsXTsSxtTBWaLNz6CYc6B97lUPxj2TWJz0uI01ihEdHh9b8BNImfZO4hxg6eu00SbiUcDM
KlYLuDMwYxBk+WF4dVHwoBavdoDSMBGV5nQtRzrXgUYMMaMxTuLKDzOLkkPYoCqBAhTBVu1AMgK0
5syI/15F3m6uZJGL2xv8uXz5hL0/lhRhg6ey0Zaq4HuXEq8vwAf7IcXRDNNzNm6h2hD6YkGOCA2y
Majp537pbQVzJCPeRecg9eKfNmN0sLgFCBUQ59Mm03O112llkU3Ah+H/kXLqidgeVPQDey55ifvO
HFCcOj/Dn9IaoAC3y2Dm/J/I7aLyau7ytnCv0lzQ42pQEQ9/mxGlFWCwsU2xP/4s7OSbBxWrk2Oz
6XjLzXS0jGVjZCIu9x02dVnyBx6cWDN9VXFzuZnjWvbajUXEEDXUTCfU1YgJx2mpjQYkBmJtpWDB
cEJfs5iZIeHxFZhQuHvTKNrLiSXautHywA3Bx42MQaKeKm7TNWncrHKQQ4wocZ1vgxR+7/aVD5PD
roSHXaHLz7fjEcpzjjObfeHF4Ry6/MjaAG200TreYd02ep2ruSl81GHFtB8h8uQvhdp3piXoJHKM
RLIBYhCRpqzkK6kUlLuSAC5YksgAI6xoTWiw8xF4iptrMhN7wiP2Nz3yENc8wIp52JJtiT+G6dEY
l7/4aK5NHZE+AFADDQ1kcN0CsmUHBR/KCOmTfe57h+Wl+jnHsejiF7LoUnAevIe4cix3K7uc99AX
6xAcozZqOYYwEfCrWXcEm2j8IZR12WysaOaxeZCEaZ8Zua3S95bSlvDwfNwgnu7KtwYGMuBEgJGh
8XuP5rDrFDGsrXk1nllkFEUFwC8bKkRk2uZftBlBxGoPRn0bGV1rD7/jOqL5GcS0F25Eaa8vSW7B
CZL/9LuwjY1qwECKIm0jr6/zWWkeCwMIKrk0ldeZBSpuJdWiLHn3rzVl+Ut1z3dt6Mz+abcMNTl4
BxvNJjU7k7DGLbdZg32vRjkZYdSrS+1CFuP+iS1i7sriA/QmC+/vIk9iBaZC2f3bFg46TVwWlDSp
3zY/2SIsB+68Ctg+uyJnDAc3jLbqknCxh2WvDz0ilehXo3LkIQLw7NHfiHlBI1d9Hn2T/CQ5bQwi
lQ6KzEQaRISVJDfKO0wp7YM0GskOhlD3XW23p6R8yEiMuMMXdRNiHG20R/qTLDbNs7RPOSxG8Tp4
vLiw16EuDw2JEu7xcnj9f7NMQTirAfMZwqvkPDBp4pUWGjcWFkyj0sw2nCRGMoZVQnDuoeY8hWEb
mXR6w0Kqguk0gV3oTXXtYM7qBQl9+3LPKaq2vKkDTEtN0WexHoxX8J2sqOcx164ef5WEeo2zVZdW
N1d4IunKWCJc6aQ90BlrDUff7XikgKXZHEoJR8bbUwUqXx6vTkwjwEp5W1Ekf5VUr6LQ56GnHrJ7
mkEOFiCF6kOZbTaBVR898fuiUSfGRjHgY4kY7OV0UP5tgjyyJxapbx4EDdxvjRWlgZRfKkV5VByL
kG0S6G/7IOx8nobKN3u/9cYlwl4k6nmRWi6t8mHEEj08xmMLA4LuaRTU2KDjeXW6BwPn1xTl2n7o
UilcCBIAi3gaixxBBmqas0EXYZWI1u59Fv0ZzbXuaAA59RIu2LvStlRhp2T3KBa3HNrN1M+FV+k8
RMVIqWETgv29UMkSLV1JKhx1eBS1AMPffRhunkqcFDQKpFwfF0pMb80IlpJmkH0/AAGCWSsj6Tt1
5W4aJ2IIrFIOGhcLYw6VzgQ0k/02uNOmU39T+axjFstumSTONFEjTR/OoXlnl+/O4Ilz7yqYtzjN
hjSZN/SA1EPonpGEOw/PrH7xl+QcwgO6ZKVXVI08V7S0TPXiRKiXsnfVY0ObgFh7SunCPkqEKtTk
/z+utFlx7IO3rZuwdDMEPuQjcYDCzuOVnhiS98gqefzCB+ScttfLIw4iUEI62Bsf9XAxrygtGYrV
+GS8K2+d0LUol0Rc3nkHPvsYH5g25vnqmjOH9eH05veXeENGE8dCG6BOQVqmyEBJjDwSS/d1ls3P
um9Xx0O2hEmhBBLqMIyrWEE6TE4jGRV95X5wMQrqn3vQ+fs99Fh4J0LVm2pmyjX2frkZ4Zardn20
NbFKfN4xmH02jvqFKJuv6fdOMGlIVI6JwH/YosWgfHnLa88zOXRQPsd5Gu35+pFW0GzSf3Bt+Too
cabVm1Nekne69rdD4AzW3p+Oi2EdZEHzR6yqDdKy7x3Ix8n8KBqQKSf2CRUmF3lPZgx3829LK0Jx
4pylhmM0W+T0OCdTyWkD5LQEcwLR3Gj4UZqcayeTT17Pn5fuqJSIhxJMgB3d5Bd0ndqAdPjue7Bs
7JYJf64H+RPgBUbK76OCNm9lso9/7VADQ3GyxA6bp0qSdArH24iC96EoA0UyVPFuxPeTFwRo0AlA
Fd5y0uG763I7rYVyLYNJNCkMdpmPEFpkNdGPFEgTHI5ynOtPP1mvIPBzZJr2DIXf8R3qJj8U5T8A
TXm1RiFdqSHtvntPeYA9xq+0HaHdeXDJXF4G82UMI3jTy+UNBq7proQB1xV/h/W8FCv77NkL/CuJ
XK1kODT6RV/S+2kOafuHXrreLJKVZ9v0sbgHsAa/ASaNUwnympxqIOSYEdr08L1AoC96BlJUSQzo
5OMIS9By/j45pVGg4CW3DaPe4PCcQc4GAFngGNEjam6XB0uobC7oyO0xgM8d++uA+Nc5GKlMRUri
MazbyaXmfit0sxpYD+rHLAZdFTpeQ7jKJFcGFHGyZwwaC42MCecYHhN0ap2yfH5dt+ki64vVIqy1
7Cvi85aN6/tC8jqSV+6X5PUbHjovSDOBvagJtKml1617LtTlPuR5BL75h+UdVu/aBz8M62SAVFEB
KLmAJ7cjSamAz7fyNCYkwjoEIkZTjjNefz2eHfCIZE1fSejalU1KcyahrJjVmC4iWOsv9Ui0gxk7
UhT0mVhmnUy+YqUGsiv+aIoOOfNWgGU3VJSN7+GgoYOx0umdjX3/YM2/k7VzSAwUZosJX3LSJplu
4T/vN6ycw169cd0yOigELqs80ejIph5LW7FpnQOS9xLVLPAV76zAaIkPRyBPMoDamDtzZMgOiXWa
/clfuTk8BguEd5H6t9oknlXOFvzOFR+EIJtJleXSb8mNozW1EwOu9MRCcJ3AUTG/2Vqme9g96U1V
VckovcKPF1dCxhZD/iikY+6MNtJ6l1Ycq2Fx4kk0Qqbn0HI47kzt6RS7npxK0HvzNbsRzVAJP/8/
R8S8zIwleJb0YjnTZXbrhjBijQcW7aec3eWpwzwoSAhKR4xXUcxxxSSc0m9i1mWoutzKKQrNkOmf
z1FlXOmOHrDEi8gGDtg1bSIJFUtIyAe4e6g6PXjd/7Nl4FpOLylxF9h9OHSOxXdLafRbUgbi9QmX
TMMi9+TATLJJYa7dnuEu4bx51fpzNsln8MWR0J+trrsehKgwTiVz15vV68+zBkYzbqQe/6yLbAn1
1yi68iI08yeFOOIsrXNO+4sG+KgETeAJMRSKPPu5gGJ08oY/P9uSbk8SZEqB0nVZZ2gxxFqV3vVU
XPpLGeEm3TL133TgzZJOAbneB4Fh6ymE7K2zQyin0BzjKXOfvdxGAAkU8enjwGYjzBiqeyF1fdyL
a5Q9ByYXfB8/58XvI+Sfs5SslNphrGLcbn+pg/MYwsx0qgYj/7/5G5GkltIxopkiek0nZdmTPwqs
IOKxivA1rt1n+u9RkOHJcl4eR2fJUOpdAyqPDSbLarKWFtaiY2Trw5ZuUyVlHwBu5Iha2/Be23XN
9qDZ0lNAEkFasJ+m/63se8fWOVIz6hqy6LucoEvwYbBwS8FNqOgi40skj0gm8KpIA3wUqnkcbwyt
c03SOsdsEWRd89TXBxhlyNrJ4hA6eWH+fWp/xYrMUIk3JiqI6GYOn1s1Ra0+8MXgpOM/IZUz/sh1
M5fk0aZJj8IeJCzimZUxsU9+bWyLH8MyoHFP7ENAOySMaRuMVSzQyVQ/YmwJkDvusFaffn1qQ7zN
dtt+RzBZ09lc1+IICu0oHAPvNfZ7dbxy0ZEllIHgspmTMUwJ+ZHQE3tHxtwfajkP8Ez8GDhE//oQ
06GudkQpT7O3G8n2Q0PrntA27/A2Ayl9ioZMtPawHv6FX1JeTvh1TPw0iRsBXqHkS7uy/9xok9sC
zJlauSv0Rhz8U1PlRihcotlBnWVpA1OljvYUb9pDBtBNb8pTzBp/3HBKQUM96omH2zXhbdgSOzGp
n2tiIactKtiYY4tw2rLjQjDLv8YM1iaceYXUaMYQsZ60VFtnsZ3VPdzUuJi6o/FROlOIbKfJeo+w
/8UPzk5LGtAxLq5oo5zkm8lBrZ9vHXyxx4FvThR2rAmYwwt7C5CF80A0o37uo/Gg1il+o5PQxPU2
5UsG5gZbf6ZN3HToP8eTqssvFDTmMnKzNY7fvvukE60g+TLPpIebnKrQah9azsd49JbfMH90SpRI
Jq5C/1MkUK+Glqpj4Lq30y0akZ82tO2xzmkOKvjkC6UsW5IgoPX4HIoOz4DwNwxOH6ZM+zr7vmwU
zoWahOMD/YkzvEtrN1R3Mnd3tq1QJwCd96BA/cuJkuLpM9HBPCn0yqqFa9X3XnRPrev98PULCIMw
ZeVCkGCvne6iGjsvkQd5kao+JzI2bAOvusOd6bl8rkmkLi+h13iePBBqzhN1Mbp91dRWotZIp4Sl
6S32c1cqtYZQiyoeodvnyzH8UaTeEp0xLG3sn8biBDX7x83WUcWQg4dBwzSYbUcBEpkdVfPho9wf
mBZsYYZdze/DQSD27RSZoc8ZkV9xLfLJq4V9vN91ABIVfthoL3GrxxR/OPkucjvIThY0xnPsEBVA
HOyKzmTtyEnEHCzs38ZcjAuqv02+JPu9otZl68KQnPdggQJ+k6RkC7P33HLkli93yai1KZCMiQiM
hHdT07eCmgmntupW0W9qUz1aN8a349YHIIlcDC5HgmGfyf7GSDiCZ9feBt6Ye/acPa7T5iuR/lpg
g0C+UtRlqCItSQTJySYz44j/GN/L2HewBiUp6zFAgVgVC+ItVGddnYH0zCzFJT4XSGUoKcmSBVsL
R1fvF4IkUR4gtLV0l1Ro1crwFdosmwkXad9iUf2v/Jne6BPdDaAWdNoYAazXJNnb504804H22uvO
QCSbsiZYV2vq2mFDExXy7pgciRbe7a/tdnAHnRpypa43fNmEurZcFe9pB4v+Cpeb3LVK1fif9DOn
sHq124v5V2dsAAnU26oZSAeCuTcFOfh+UQISbCgTmfBos9KQ82G+KHdhE/Hu8ctjmjGjPDXKw4EH
3bu3NA9UadvWxK98vLz2u0uqcUoYaf9lEst0i5bzRgCreEVh0kuLPILCmeWTURmvzia+PnTaR4v1
l4W7yyLGsInDlPewxDlknjWe1W4oVCTyuiAuYGpbI4TGpc2KmR7dkc7KnBuhytifbxDxuUYfrG0K
BvtbAYrgJZO/kAEbAJf50Lye58f5pldO+MwvXkBREZ8s9o4PrN8xaDqiLhBltIP9Rc4wYGhZ8kln
e1vU9cWdcaCu1kLRJPMv2BXo2QsaJSMhLKUiwHxUUptXerbSjNvbH809onj/BhsbQzOhAOKJ0dU2
IyP/UBYwFhgVLeEmvxICczewoVWXxNC18frGpGiIjspBgdV3FSnhukV3KCIMOnkauvdVg5CsI6OE
HhXRIHaj2POjm+4r/TAWApWVD8wc+Zh+jpxqCP7zRTNS2TP+eXOWovt2nYsC3GMlewzO79xEevoI
Bj2m/UTouQsqZU1vIf1wRqzwmjfbIR+pQxJuZDqTQIPVs68IM7qZmF+Jrqpbx+Smtg86YzcymDXa
VkXo1Zt5T3jxyMIH3P54o2UtU4rF62vaRBfu73xqCdxaSYL+OS2HsptTFiWSn6QMbEer3Rxk4kSU
iDN2qmwJ1kaAD9//4n5HDcf4mQjufoivcdZTugH16FWwI+94Zen1JfPkvp1ZY/bFWmTaOdZbPLa8
jPblJiSP0VGl0VEebyGdi6JomstN6Jitr1eyO0MhNtVHpVUbquClX16MGqfToYNmznENoNHUgo9F
KapcT/gvZFQf4Cr8zedR+iAWwO70fvMId9kXrkp9GjjSevAbTwx0ZCOhfyfX3o2+zZbuqBVGGOuR
oryUHQsGc8YJHWibRTHadcTW8OOXQ0lLzShMvZmIBJ1sDIgczYdFAqJQ/fpiOdLt/4JH9Kpc0TfB
Z6/RnkW7uN5kh4PH4pMCEu6TRsC9ZvgNcM5rkXvvBjmygOQKFWcclI+pAx3/xFAZhuYxRCHo3BZu
3bCqvWuCBvx3mLBKVri0mgBfU6eLaqdZYmYdVHpM/inXsUjuQDf3rOW7ki1fW93u6ZtuFCRylEc8
ftlCcbis7mRy1ti91lRU7E7+kVa4N6449vqjvKOMh5K9hL/QApRlskieGaZ9cpQoV+kNELL+oemO
uc8YlVE5RuLnElkX/SGiYNfn2YFbXq71a+pO7JKMYeMjCiudfi6YqhWAh0kxc5VbAGzNwMAALBhF
ileDr6eQpBuK9Gp5WwWWRitUBAAqIbFXFXnHv2TiIaNWTZwL9gSUk9rwXwn4cpxOxB3VKfeWoMMC
x+poa8c7Id1NqQxJbonEE14hT8hGYreuSBu/IlUzEMh4IEJfXAiJgFpLa0hSPH5cmlqlXvjqmPis
vFbErbTXU86XXF+C9sAFKJWQRks9HCLjG7192lSl834+XFi86ZY5uqyPcdkgGka+eW/1t+OHNtVK
/PkZh2Gw8qnrPS0/gjwohOaXlFYxA9nDCyfuNuvl0etjZTO/TjOWltx5Yjo74OT5t0gt5HmAlzbK
Vs8Tj7Itv3cnDDVvh7ukwOJnO5ghvWXFJO8+7bkFnYGJos0rjzbUREarxs/qnxRBAbcbqV7qWnTU
fvnpyrn4AWelZ7fdQpPmFzWv5MVyr1yxUhz8GVznn7ViPfeb7ptD76miREpJhN5tnRifuL11Ed1R
5cE4mbzyfVJF4+1r7sbOOvjtAy92cK+7uz8X25/o2/W6VoCuf0hnxZHPKyKCrXCQQ0lSFwSEmeBP
4QCi8Xp8ZsDzyLRu0SgETv+ijQLpyWo6B+yxqN+g84POa7zxBWWPT1sbaNgbpyWSm9TMTvzgqIuA
gVOAywf25ETl4QyzA8WPnmp4Rt+EUENF3xB+9b11z60cXmkFU/TahZZN3PR5cz3pfZghEjjQqxNg
Xv5PKQZF1NUAcH0XJTmzkezh7CJ97+pXxAwycvpGaOQ6Igs0IVHBruwpvePbuRir1z35itFMYcNB
uq12IPzXrqjrwutZ8CxFDFjpBwcso7+7nY12QzoHvrgB+9o+s5rZOHNtub3FyOd0ND+XuGK0TPI+
HvinfDMbdUxjQR4z4zuSXAYaKEPKihS9ozgK4FyeXmIGNcm7Ue/8d+wm5sVRtadxFfbXzyZY2g6O
fQupilGdOyK+54BGeobOjwA1r1+/of7J3GIAeEdh5kglojo7MhnabfZjd+80TS5ZkI3m2SRreDpv
BeHrMiufWSz8asZhxQKI+Lv+Ng9lwk8f+w/0HIgd8WLr0CUbo8wmQx6Ybs9TExPQ9SUYjEeDDwcK
Ytb7wIEQygHomrbpeGmFhbiLndYNUOn50DhYT0qEn+jxx4r3g0JQRAx+x+JbkE+qyZ97Zo1+GPJd
Xhw4ZLzDbcYlAip3Bvz2ahocZez3j0a5AgV1t78iEEhLk2iZSlX10vr47Bl729qyiUZznFDE0m+J
chkdOjLK5KlU7VfaFISjPUi8xsbGDFY4Ckv9noKjHgCUHtLQ6ehXO0INKFDA8MEgCI69gv8rOyX9
kzY2PXc2sieRFJgyoSfc15ZeCCxzKk3X0qB8Bxqlf9yogVIRpR53jcaXv9KLsZipCTFeCDPJktTo
cP4x1U+JZo/sg1csaHN8itqpbo4tln2hqedDEOKgqmQCrAVHIIhhPO1b7op6//LqE9THNBzMaupg
BgIz22laokl1g8d3MtvEV0Lnf9YgZie2Or8+vfWGIDSi6W/kKkU4i5AECN2CrXUgku6wgxLXFY0f
Ibvgj0MxuMQLLH890Ew/bqjFEkGFcXrRP8WuCTze4/AtYxvFO6fbjqH86wl4pzKLSbglIltNqaPG
OkCb45IsNGZbidQuJuwhkMg6c7bQeb8m2yhDt+1bfHb0uKl36+KYrpv36gUE74PVSwiPTL8H6VAd
0/86vO9/PG66TLyrM96Au5CnJfDAGsk5xUzPof5ltLpMgWDI46Au/hG5UeGs2hzBMLwumKVsnCzz
XUP/vlJ6FGnOrOqke7BTwHFqjUWFFExnCSvmjRlsrtxUYWRhGduL582T0f6UaAaTHqSo6Se1go1q
VEhTOI9W9u2ElCCHxhmm2a0Mo/N3dN60Fvtfz24uwxMBHWExafUvLX+NcUaTItpU5oLvDDJIPUae
e61bhxfiVzS3D2H+CoHT2MlbQ499E7LUXkhjaEu/mtQ0+fp3EeqPULKPhIHAXwZxrc5oixUFCO55
aES0p6VknQU9sDE51eL8we9yeXZR6NsCVlQT67mtP9zYA70/h79y0MBN7VplCephKXE4f8RTrtHE
JL00BNja+hfbBczOsW+ulGx7GNijknvOXehI9MB6hvCXIcacnYJrF+WvmwV16Yat4cFtdd1cQc3v
AXNbzaJ/3vg0FnKr3qjSiX+Nec+5ED90Sr25/qD2iCz8RLC8sS2CD9SYAfUwBhpfPCrdXlJPypE3
c8EulTBLo14yexgKDc82Tcnoh27lw8m3T5owN9P2ZNwGbegxxyoCl+BP+x0hA3A3eMDpHUf4yxc0
3EbnPl02yNHR9EsOU7n3EDWU8Wg7+D364TOphQ07f3Gzwb8CUk9Po2Sh6UiaB2v9fuzNOCBktgNP
1Wfgd2jEdyhfJSFd703lKGCYNV406+S3Q03ibU9TfO8mxzgu5ndj8bJKaccDLCBP3/cP4BM5GLni
pNizX/1wDfZtBkvORRNX8Ge/K5QBLqZWrwRZFIfqtcpMEyqXj4nSx3TcOtaITvqlPCkkVSAgi+Ue
5wJ3KApiN4GhVD7X0SmXxhrb9Z6QZWLyKpB4mxWB2MFvTAZbIXbSXa+BZFWGYU4+nnm3ZeTqgWQt
SnF4BC+mcRrGuQzSiRcw6Y2E604elfqFrJVgDnIzsDteP5p92rb8gkym6jStwUQ3J0L3n/Tmzois
qPzQWIOlv9yVJMeefdx53yYIs77IfceLuV9MXHER+zb5WUCOgNYrFeMxiZmOd84KgP/wOEeLo+tS
aSWRZuBbNYlrMkCTPr5xw0BGVQIU0KyoTFeC6PWgqSiAse0hqkTUbOWfTN6KhnWrBu/X2jhSs3rv
lO5vBoQ2nFLZPPaN5OfzRsizIjsXlxROiXmV4ve3koUDhRyZ5D40MoWgILdR6dsnE7+irfWAciGc
01vL22KpbUpbil2k9FL6vtsLL6tV3t8EPRE5Kbp45TQ4e5CMhHJY7zr6jNCNKXMbcF+s37HZhaKf
koAYrvyKkJGuPoLg59cdVBO9buPy6R91uzadEmImVhQXMCw9ocA0B4zeX/32IJEVz9sUFiVuwXW1
zqr4nQUmudC7GIwCfx7jefWewPDEK3YEjgTNVN0As/AWPko/Qw1IvN6mY0T2W+5QnYQpZP02w5LK
LetZFjtkWRy9OUwWRT1ea+FRzWjcDaAloHnUMqWH/y/tbOkfL3s9Fxxgf15mjSQU5X/Bgg2NSsDN
wPmZLcz/X0uCwcheE5oZGt78ycocC2eXcaGrCKsFYdvGI24e3NKcEXwZKYU3eWK2HuAb7RNwUghs
tCw/usxOqwnn2Cp2ujrpmGpjTr5U6nF9ckIaOBrK1aD83RXbCcEwWEbnHgaNAJ4SNqavt9S4AUC4
nJu6DU0tnbYt3R8cZFrTofUtv/C9XM8TyIA+CsmvhzUmnwZheokqyJbXVnyOxTMX4M5FzafHEqm7
Q2jMAcSW+bfr+/lsAxouko2e4sevXVUDrxujrxXqtb/1lZwh5Pk+nL1NnQ+Fu2gKGD+kYwUZAIZu
8vzRrFSdStAhH54GFOZccG+jJoQ0+jOQzel2gGLWI7rtxbHsUfRMOZcmT0C+AiHV7gFS4QboZTUs
kjO4mWoGF3oqTkPFfYMmsH0dyoqvFWK8ciTNlOEoih+VoS7Cu9lgU8l9DTl9DLTuY95SB25VZRQi
eZzWfWUx0lFZat2IZXgeLsV492FC9tm6n+4mlFU1Oj9Nvzf7a6E2QuO3AwRVTV1ia47EnnV0nonY
rY+BuQ/s9w5rLYehN4Kb+QKChQWrUGJU68iuABc3pUtr3GFmUZohhpayVMicD/uyQy5uE9i5cCPx
wll7y4p0tSF6IOqNUHTH+cao1RVyg6r1mGNAmUniVljA7XC6AnCydiIOwTYU5oMqgqxI4/VLy8Xg
jMOLaUq4hj4LiFxgXMnkkncCGmIt+U/RoObu1YAZrzh5ARVZ8NlmSEK23q6nHZ+pTa55WZ8ItRki
/SJqCVBNbeo7wABsLC7ZuDl+bgCBSIDQfwsic0/YJqJqYsRYR3kkqttp1zQeKtmV98FIBM6Lavke
WwFSwmgRb2D7k5VFTCrKA5zgiuMOoOxXKCFNzHd4yd1xbEM/WP7dQSigLlKX6tNsG82zxSciF8eD
AW4ObRGJ5/mBE6HdbdBUu1FK1rlrbqNK6fHLrlnV4ThBkuZi0W6emBCUTaXaVm2jChaRp5NcWE2e
vC5fLXE+ZGTcXlHPeDncQSAVkDbc/OmeZaAO8TvdzFlyorJlTU8JnXsNPSJKcENktoez9BVeLgIS
te8GS/wOuJxdjrgmdlPR+yCSURhhaNvysCHNBnegW3urv6eTKK5at70qWfiMe0XQWu1tDrmI1P5W
fTmmgF3x7XMijxYAUnFNthK6pj8s54QSH6Z0fYInhoWcCFUbTeWkYht104evlYndi8PIkr44Qa0A
yJe+DPGAqdnCkZjgCwJf1d/Dm8xD/i3wn8U25vu5aCNOTVzFeZ7EW1LN2A6zG9UcuykKuuitrAnX
AG3UT7dudxy8fnhNWybKAATK0JtaHUpp3fZitWjamKMlRRDm3+R9/Ky1RCvhADb0IBxMufAm/UVs
W86pJ//wl3rOzVfF9N+i7B5pEWR53guwkNzE8DaBVi/Fgbx3/kYkPh4s1umD2lr6xrRQOqXgqTl8
L9VzztNetQO/VnFdSDgli656o8AruzwiU+1GPwyyI1zNTaN8jzesQvWUPtw+20iEywrK+xMIUZwS
zW9iTgGn3BXYGePK6dmntNsp7Jl/wpma0JszgqQzodQeyygoiZKXCQsDmQz4NrnabTIWKJEL9zKY
h07VVBP7ppNV8Ta+AIcGZichuxqZ/BYbvRYpuBZtGK7BF81NXgnIIltmv2ddrwXEoKFcl0/lMaYa
rHe6LUSaAacjgWiUETc40SE8jz1/GdSZZeRdmO8PyLT7IkuZZBTKYiHnTjQfv23P3bTlc7i1nCMI
IjQIu8hkmm6VWrALIxbmszYZeBCRgUtX9Q6gEe2ZKBe6VV0uVryk8YYjdXEQQRm41OENMrK+ZZPI
o+2ha36hukTTgijj0lOfX/uJZaQ4ru8NJ6XV1nGgMz+yfHGFcRH0XOX4mg8sCALQpZPrBx5eK4+a
4D0NxX5UDB4Ea4Vkl0q/XabeyQv4Bu9CTS5WWUJ8qS0gOVIBWUDkqc0wrCHo0eLQus2fT/yt+teL
Mt1MJrwddsFji+rvmWF8Y0HPGt0zPN2kaWfUUqC61I2bF95QlsOoMA8qnbe22D0dBXK8Tk9nhRKE
gbTWn6HtkI5FxYBKrnVAVgP4/DaEcmkJfA1oFZfi3dRIvxWdU/ktgoDHNtQ49jprDiuNOPMfwBBt
wEMfpMtIRf8wif+6f4jKj1TSDbrkg0AOb8rxo4akU62ys6GPzELVYGkzukec9wVh5k4gi0SUQnLs
GJQL42XLy86CNcYTLk1SiVOtYY9uEYgAUOff9MZyWkyiZQuJ0M9Vt83IIlKLKrdOtb5ZsbcAA/zU
W2l2qwMEgGsDSPD9crpCIaZ7z8IHASWd6LTxWXRJVRAdm7X1jjnuS1Effo4yvsQrARP0ZJwXfTHB
ITq+ZjL3xS7y+mscUcWFbbWaTy68dn5/NcUCa7X9BV4TSMXsjEdwAG9DBAsGtEREtBl0F5Bfz9LK
Z0Bp/N4RNj6JXWmUNHA1TAXH8xIGv7Q0a4Rr2D7MrKPdT5dcFNrBGvvFd93sbcrkX+pTWwhgzF36
gwxStr25MFoxNu3MfueUm3YRVY5l8N+OIsd33qiU28k2YFNXcPYDTk43TgNhc34MzWst7uduNjj8
F3i2aVjjeavvgI11tbp42/1S1qHPpkV37Sl5pdvAcj4h5tiTmyL0E01r2Y+6Tiw4PpT9nMewUww/
So/TmP1HLYAZ6Ohc0sae0dKxECCyuGjXgrYnQ1L/YH1ZFvcwWDpzqtLZysrK/H2nJa3+BJY6Q505
+g+bk384epxDzmLQtaV7ZOzwJfRqNBFMDu4VrHkH1or9sCAI/yc6/onSx3CrzDseMNwtsoF8RZBu
f1a3z4y0oPDawYYHmBWeupN6jnyx1757bLNluvfaZAxDaYu+k+nbe0tdrk/IswAQQFDQNdZR5sYP
vWp+omer06RvK7RVSVyLlp1TJCuh+PhrAGLlAy4H0uAw0aKmYGvWR49krONVfmAke9TnVYwkrMUy
1tDC6dhkYdAPziHiE0PgrumFBrlSd/xASIp/P6e6O9FhHJmUvRGqpDyz2La93haTC+GQxs2aSsi+
PTAsswc0S9oUlBkQbgWjWdHbE7aujeGBavd4OvmLgH2NkOrxyIW3rwRrfkMWdvcAsqleG4QFov/v
gFXnGEzx0bCBWHd1+bLom4qILbVX6eePBnQmbUYt0+Q0Tyop4ivuW0zdoiOBy8MBV+m2L01WIlHv
1jAOBxTWJNvvrCRTC1dHfKh9ot574ep/ngdaY8A/2hlEMm/XNA99xuqiuEJyQAC2bsd2FzvzGDmm
bm1dfgFyc6fZrn8W2GKaks85J3BiK7UqzYJMkaCwHuADs9Ejmr5o7ySML3EutIhf4v0P8ZMW2PhP
AIWpn7OYWJaUn7xahiilVw545aIbvYap6TtBuZ4eGszyRgKyBC1XDT8ULvq8xTCQA/ELzRPtlSex
ZemDFbOzNCeFLSmVhN98w8BIdWRmqIvHKmddKBKrF5065XLYfiOazQtFRKgIibwqqY0VNB25w+LI
Xxg13ISQHHRRZ7gqrgS2VrWnPv1aj5y+Zpbo3aYFzEu5rWNaQu1ncWc2v9MyV4Qlg4fhsnRpjnHi
6hdJhS24Qda0jgphtqWE956LxtTNwXAoEIblC/wJNV2uYtYDX7VkNi2Tl+1Y0/uizpilauU8AaXi
rMHKtxfKntTzE1znYaRGl0zUeuBmwm2C0aWjIM/7vyn94eKERO+TyUvXHpVLGzSO+AYu4lM+j7Ll
598oHlip/g1J7rlli8jajAeZov5vbek/QBmuzegnCFpBM0iEatR2EW7ty+IBkjMWpyXLpmDCMdEN
wdC2kRl0n/SLLbbnNqjPN8O2QX+2YqwsXhzMP8kWO1oJu453A6toNxhugOqjs6iuObUtAsoPjg7V
j27zihqf0tAJoFmGQ/5GMZwRk1fC6wVS6KOqDD/AELQr6IY49IcXxp4016UDM9RwouzgMPPwejiy
xlfb3MrY3uF9F6ksVgaesiduphbcbaZHBP5OZNNSGgK0dni7IQRqrZwPO5C57at2yz471PkYOd1b
x85Kt1a4QMUEdZQD289AC1CjKHn5vMa5uqcOHnYWDL2mp/4K9mRohQ8XGo96lIgzAcdYTr9NnCga
avl3r50p3PMSMBJceYdbZCMg+ip5h6fi/4LhJOP6aA06FWpey5XKc5cSOyaw/mwKfaOy1bnAeIg9
3TpDMb8IB25KuIFjbIIDm1gz80Pq9mliSIdT2/11H0UvDtRUwPZWWIkKyGKUcehAYgUmY1T150tJ
40HNL6F8txSbTJLi8nngi/f0rziii3tUtigEKgPKce2Lpy7bcugRjqFO1iJxXdAphyt/Ug1JiWcb
4AGzn9wXIFZ0X7kOL9JRCI2Lr6VGPuSvL4qamlIP9nii20/Gl7+q4PvoUAeTaXfHleIenxmri0Gz
8SRlkzNi9WFnw0uPZ52E5PlAFuL7g34Q71HSXgTtmFBo9OGSUDW62As2yCGoITONdlV2KNi+34AT
XutWgfNgckY5zwxlCOvRYKg41RMrzw/LJrxXX9O3nlattOPc6TNRJIm/Jw7iWbzQJYCcmASlT3u1
PvlohNyJIrvE75D45alNnZvQEb0lhKg/e8eMFhTkhrev524KKDGmv8QqISgzcYXdc5f0UuTB2u+x
HxFPd/lh5xIStun5sfVRPqUKjY8Z4Akk5aIwnIEXJ8lMFlMykGuXhR7STtUON0VmcbBZn/kry4yV
PZ/L1d3DMUGAvLCpP6zVExZ7aQqc6/nDBQ+Qxa3kA4zZzGxoN8OXDvqDzEYJBQaVUkzE0QqRAL3h
qwXuFTAjsZcRt722y1xngtmZ42AUBoMq3VgiYslakpt1MePVnqPPDlxqg/dgh8FG3OYssFW4Oe64
lVlT74X97a0A/YRfzXJIuZbWO5GMLWr2JHwihD5je9DH8KjRbqSIKukA1QfYlVts9aI3MJJuflhR
2ymSE2Kb7SuDN9t7VD1AUwQaFEY9NkfHKxmKE3hLXdID8KAVj9cd9uJWfheI9gNfh+Nr2utlX2o1
6e8cwi6Sq05e3jas+yVkxX1xlvhfrq1OKtYtQrb3R0ndv+lMrN4QNVji+DZzLtGmD7nha3aNVYl/
A4wxywUH+vu/g5d8a0PazO1pYFwbPP2H4CDjK2zm383Bly81m5PKMeLw/zPTzSTV6wcKMzkC2L0P
9P4PUF7v5oKMys3eduTJxHzmVMa9bvHjk8J8E2BB97gJz+CSfBo1GIOKSxaz4NNbzZXE2GPn6A97
BXl2RurBWptW672GZXHqT4ZUzUVcWdimfVdm2Nefx8Lpy5Ytso0YASKQE5HZVNIdM0+1UlVis/CS
S0hnkl1fQyGnsfdIoOvdYt2X5LKt/5w/aqJbMm7LFhyWnA7Zcr6N9+5lu5r8e6DDqKT2IehLHXSf
c1gHOMwt1QUvTurrBBs6uLAiuhqLUzIjt8nwIh9QPSxnviz0yT+7WVrUaN8k04J3uo61L/U+9UtO
3UmYkSJ+fjcgb38Pe1wVoVuCQudIWjjY+dWUhEwfgrI4jyS7r/OKzX6uYwGu4ljKtiA75QPKqwye
qUoC2dAcxuzgPYp1mjbDP9G5b9xd53BKw/n2K5QhqYm7K9r9wKjSASNe7C5temf4osNiLl2kl6jQ
mX4Yd5+F05Cq8uI07L6r0RuLfaRuXqeTug7RmsxbfCLsi1+p5Q0FcIoUaJgCCm3OIjpPkli/gBiI
vNNsHmqthvBwAO7Y5disg3n4Y0NqQk2k7VbehPkceZis+ouPGb4YBqYqSy12XWni01xT/GTYifxl
AdzH5SdagwrjjWMJ4O/gncpr3ttqrb9X8vrzifk7bcIeaK7LFD609lWX9Ecvr+ViXPJnk1HukFVX
M7viXcUV0gi02T/2wyauvuLae+2gAcpCgaJMWdDa0vI3674W169SQU0QJ9xS1V//qLKglZTyY3uq
s8lkTGu8dLKaJ39Cs6d0qdvYQF+pFxcCOITx/GuheYjxeZT6wdPDNkP5XopmCAbMpmT/CyJLmy9a
IaqADh3V0c4xYgxH9gKlKqiqGDuQMd31cTMJo71xzBedLK2A32WZtoby0u3WM5SNZukvNM5JkMbB
J28rU9vjaKUc3fEDjCHAE7HoOZ6bs85lFqykSQsiJrnfr+sXlm3X8IGErXTuyR24oBV+1w7raN+Y
+j3mfvD/65Zs2JBW6bumlXU4uKbiWEQHSdwRp3ncpmyWbFpaoHwKft9S9ZlW/Ng3bAdBgOtcfjBq
qsjFmEc9nXMUSaGz3GTxqmQhl5b9WCl1ATI0QwD9dqENO3mdRw2HSsj7bf4JYRYQRcjT6lpWKx88
dsC5piuJqJcgdjuWm1Qm/GohkQiGA/1OGCOmcWbYiRd2wV4Q2l3NE8kWJcHKg8Q0rCXBq2VOQLSp
aKG6V1mlQYLHqWnVQCRLoS8CmzvFYHYoFh0TgiA/7lzwjLSxIna8GwWYJQVQldVhhCM9mLVWz65k
W8R1GKsdPbtiTIUhK+lEr9YDcVKLTE1J4MwXqqO8/2KRcjfjUPzVNgtvgUTzF42Lj9MgMldy/z6X
ObVkrZvcNJ7t2DH3dxEaIk07816hpnj6Gl5075ERmy7VGQSj52O7WqLIdLNQSoosgfVO/1vuRACm
6nHUc2fraKjmtfDWGjBOKW3lIhXQoyxi7lIyOADICKEWwnefyt751zHf3QkYRI+Rljiq8yi+7zCU
aAILdujMUmUxLt0CT0QCxcCZCy+YHZmHphzaP0pmklqbyuA/iycu8Wk48CVbkqLlAy3b4Qscjpq0
giUK+nppO5WFqRAgzqrC/fIaTI0DJH9w1BUyKcUxKzU6NQ5sxH2KMWjg2SA7Z7WCzuLo6iQjRE5Y
AhdtHFvfKNk5f5yW8UbIbQ0L8HRR2RLddop8NQWRWa0fPP86NrEUeMQc2knM/BHvq4BRhfu41Ag/
ifIdD9BGUKSG9Px5Gh+W0khJSQIkB+BraVjvvY19XerxgYpJAjP/yxRVOVe2VDZH2rfGlFUlQi6H
4uoGfISflu44itI61oFTkkdAkLxV/FfrQkhR3GmVM6iUAbp2NMJ1JhlAaYi573S3s8vih8hd9A8e
jerJMmzYADz6S5ApBD7hcSTqBomD7A39j3EqvD6RjjzkexvlxjucH2BR6Yju7INyM4HjjyxiWqSC
e6jMKxIHnEUgIPZ3dhNEpfT46abomgZokYby3KzT/A84PcBtm0g+0J4ceuPv/TYLRT8gwXb+s17y
2h+Gl2SKPKKQVQe43jG5WB24POydCzfc0QhmAVYpNZ79ys0Hn1Ml2dsbZebFu+JZM35IRxYhTEkG
f0QMoXIcxGM01HeaaSiS0s1FQ60WTul4VUIs+M6z/db8n+ZtcvNnZoAhU3I80qzzfBwl6X/1ChEl
t4LpYQ3/4LxT3RADupDtWZznEmC+UYMaO6JzpfMcQBDYzmjGZ4CBvae3I1EyFQjUB2w/6wCPlk4b
aLJaD22aoryXV6NlqohkTwAdOMXp7cjH2b5dEspPtPcSEh2s7VdFb3LfG6tUq04ZSsGOwABknxEH
7su3Qeh2BUPg//bnGH1WcM+HqH5k+iRHmILib5wNMgvY83fyeBl8pCwGxuKZD2DXbAoXltf6Z8bc
Au4iSoZFPeb6CCQNiw1piHbKLI4MuV9tDHUoFKiqeVha0vsJ5J1mD/Mt81+ZO/P/sAACJfKAgQD3
raIH6QTZT/s0eaadeIguF8hAQh6AIdm/1fxtlKSQE7i2Nnpb4i4f4pc4oJRzxHCJvHVp21g+kMNI
bqUuEk96TE1rCupK6auvZYqRKRuvpubT88XPtl6bFi05S9KMnfwF5dIItUkYLcKEhRCb8fPzPAcJ
krtaT/kDL4gZMqN8BPid43GU5Q3c1YRNY5SrlLB945y0ALft8gqbSSMVRQvdSW41G+vAUNMnlJsP
mTxfllljHe8jL+30gM0fQqtw2QMP3dv6wQTFZMOzPDJAWrQdguedgbQ7GHnZ5mTy6ndN8nxlWSll
Pr+1OlMpTPJ/5JB7B8hqtDMj3l/gpMaJB4XdetvcENUT/VWxFbCgrwRWOwMnU6ytISW0oCROjh/3
n+eL8o6bUDgE616iemEd0dB0/wQxaAPdZzS/uhztbWV971gFIxg1Iecjmvq1kyV7LNTFDYHxZGZ4
/rXm6pLlNethop50jP7k5j/zp87JbNoxlLIrg/5IcmyULN99g35vK0OzpPQtkhqq0Gax3RaFkRXH
eJn5t6G4W8hKfJD5+NGJtiLnRzvFFLELWX8Vf8JfUMUnFy0CSk1cv7clQEPP3FETmpuzpCd9NWxu
rm+zuq8xbim+hGea07b6/evYZt5JWC8YO5ZCEikC1O00IhcRAiLWV7GCTZan3x9/uX94V6plrdnG
Knw0aXh6oqsRINTi+MQu7SgDyusXEUSHG8qGToOzvXgbtxESbadX0KycYJaHxeDYaLQci1w/Vw6e
uFEFFEVblUQIumTV3GFtXfPn4t76QziVIFYi7mithztnWuOjeiodDVhR7IQb0hSmsMr/4jlu5Gcw
324XXmBRnNnIi5RnqYi6BDV/BqBh7cl8IF9w8Ko8iMbp1l2Ufom9+jSDDLJ9y77HG4wON+xnBMYL
0QAn6c1MGlrfsaCEsHSPyINhNCShprss5h8svWRVa3GA/bH+5bqgh+nTVTJdlmnIJSAGqECg5s8i
4LG68rQDGqQvDMCuuqLrAi+3qttca7z7wTD4eQgsxcyr9AXc/pHVMMMBGDxHGJjy6Oz4RDzjpm4B
WtkF30vy/g8Vrc/MhwO80Ad4GM3ftlxXr5j9OeMxU9QcnEYxEN8Cf4L3PB+fBg7UrmHs1yJOe4U9
s1p5POo0O/EYR8t+XOKeVudDR1hctOpkEdbl0zycpdoitbzM1r8mA0vPDp4iqLSZS7WqkZlzCDNP
6cEnNTsacz9lZhxhqlGGzsEzP7pL9iITVUshi74JvMR9dkCVIP3wTFjzaxl96CAdex3AwwybOVqO
KUzVtGoGhOJsb7YoH4Nbp+qcXb2BjrP4n1O7b7wo2JWaifF9Q3YazpGFxC5pGF8yKcHJmNZhiqLJ
fKeq5ZZKqCiy8kgickoRcomEVUNVRIPVRY/tB9iWoT/eIXDDbVeiJujwKuEXNFeKrmcSY7YzPBjq
i2xDA7gHzLVPLB57VoVkO2kTgFUQ3c6/YLoUEWjnlpF22KjGV59yfWi1CIV4otdNAx7Nkydnocxh
QMWh//JM/+sHQ8jNIHTYTpMwaAwEF6Cfz3hyE1YJrh0mpCx8JssB4+KumwqeZ6MDwZ1mDKSi9dBL
gsKv/ENNHQVCVhdFzwlWMhgPI083gDEGElzSr+UjNjeiI1dL+ZmnLLySbnThyEkdzaOWCmT05nKF
qPBOlKpb6AEwGFoCU76WjBPblJBW4qMxi7LB8yROObvODkq3KNssvVy4zNfGyMbNM+l+h42T+z0N
EOhuoCAHi/CX+fpPlkF9AdHPWfa154y8EGXUk0YgL7t5F6kwpmUmLFwpaNHQDTcH0qP4zHNyOSgz
yzxUMS3y2Ltjpjw/XxVN7sbodDhBoA00ltKmO98vfDavQaNjAhN0jbycSbNOV4iWXSYJvJJhlRnB
oXlgtuYpemkKFh4/8dwj2shu1OX/DmnPNDyt6fU6d91du9gjUz3LNPU1o1HCQbj5GGJhN2zrlsc9
5R6kBOcoblCQ2vXlk0UjMgul8tzI47CmF/7ajizr7YfxnkaKLWAN2tLxY5o+T5YXnci99ldIIzVR
zn9J6gnSB9YStNYVez1ST86aKWsL+JO1Kpwqlxi0GNxoqauHhwRsquUo7rNRMkqWoURweK9pmFxi
rpHCFQpQnXWZWnHiYKol/TzfIVHiMKiXJprYVka1oX96NkUz7ZaHrv9W1vInYkNtLnyz2y+PwwZM
IFrL7kr8ogcIVZxHnyY9nZQHGkHGxwKIZctbh0VkbX3vjLaV6DRjWAUkLb25uXH74bAdI8A/h3Th
lSSz1YWeFlLzYHvr8WSNgXv2yxLH09uG92kcXBJdQxSXDEduqRc2r5+4W+z2lqZlGFk7rhhW/9Sf
uEACbbbPHowhMtIOhbIKk8zHVi4OT/OapX0yj7jLcpeD5Ns4g1jYV3YwQHYS3SR/V/Zfsw/TopOT
SVtuV8+mifqw2QHWrDL/x+f+pv1/XOQWidtdB65GClGNpgGa0Qdyf5mwL7bUU1LuyF2YNsPg1SBw
aS4vMjaccmmE9okhVpM5/hXG4iHER1P3zPEEzCIQhvCBjSIRLn0JWE+QcIIFC/ntMkLZzrY1Ogez
7cko+q20J4TM2uVzJw0koyk9Umcy46UD21oPKliOSFXADnLsOU/+wy+CosMPu1XgDCyg8nZl9xdl
H99AZ0hb4w5o0ybfnA94ZFu0cXPC52DDHZEKwMcj7kRnAfmfdeVa3Sy7QH5ztdTKb1Vt6bNBO5R8
srLn4IEL+CfukVzGHhikn00C3U8FbkqhfTJHXGcVNlY65ml3Et9pR+BRyeBB/bVOAFR1NHsf+Jvk
PmhPOuusaPwnQpoGPkjS/LEbqQm1H6r0Gd78jgpg9D7bSd0nWZFd82JtOHBKyAXUu9EU3OvKJC6f
x9AOGE8zJtNSXZtccSL9v0onnXOm7BF3tZQ6QyZieP/RIMVY2c09pNqgXZtxGz07TAk7QtPCEpg2
Y0iLc3SMpUFTPHAxEwD00JDFRSZLWV2whGm1oMSZYC0pjVN16+gEQHb9Ao8C3Z+PiacbEQdW9QkU
xwEnZixsk/XPRmdpWb/+LMGMwvdj84gBXxkyUS7fSsRZJBecaoQV+24hTpfQYFJJ09CT3pU3FLYG
EwFz223yTA4aourQo/opMLFEyMWQrrVdoBbLCJEjed22gADoeHE1ziX45oRL0MeGYonluaJXMtOB
HahuvsEGjCZxbX/O984T9/BotqKVXswgfcJSd2OSQwwcjnBGiSEmBtdid3lmrtyYoBMI73zlRsnh
ob5uUR6iPxURTyEuzeUMAPHMSMz29RTVKgtUMTwu55GpSl7H0PBeQphvHDs10PPm/afHyHy6J2Ol
FC9OKkZ78/eDb0GWG9B9ox5uhwsGHQCpLwXfS/fIz0gUHyAwEh19LjDtmuex7V2ZDeYJWeD/CcAL
518gmeuAXQ15/NHfpVtupmosXqarWvE/F/NsfDuTyGMAby14qgoyTfHVNSg7UsXvsNsnX274Tud4
9dDHsv25NFmQsxZf3eTlM/qmNthg9VHwY4CkJxumLuSI8/y3hQp6VSvSgKt5ufVtKi6WGDF//px7
9ADPFseVUdBS9tib3UEQNBAnCmIc+TM1eo89wR/k1D51oadRWuzWc3vAFy/lGbxuV6yz9JswrHKO
jl39aVqhzxOeAI7Np737/Dfel2/nz6R3jLV46r2EUqKC5XPpnO6azT3FFLJFA4ZqNF2C8OBuqtF+
u4dFY/Q9Xl86kbK02DxP18Km2nFQWRnfJ+qXy+fEGEdmixVf+iIucVIYKwrbu/q7GUIB1uaU0aqf
pFV6IcjGZQn/5WZRAyTK/P2gxOOWi3+N0x3coLLuG6rt1YioU4/klAsAmW+DttetwhO6AsmY3c/x
7PMOXUnsP2My+dP2Lf4H5PNqWWtEBjCOwJW7hlcDZ1bgpoAoLJZ44WPjmXuKvI4kdYVWoEovZdTr
foM+ySbk2591+uVZZvpPemsHFPdXDo57kOotFNMyv5x9dEj6l33t0lQ0s4SkN5fJeGz2jPTbF+0J
cs08AvCLzEUJjRGaunYu/p0wZkCuo6c/kczC7XBCT/uVKjksYd2s+lhdD4ZdsiADbDWnS5VgV12x
RGbIF6JZPcLi3WwW7GKDCzQu80l39/IWhyev1u/M4j1h9e6B+wbg5siftrwh9dGmW3pSnWB6f7Ve
HLDJ3x2Db/o3pIrC+VDQ4+lpesY4at6CUuQtDjLlrJP12eXZJERAFgF0tmqsvvuc+GOULbRWM14o
2v7SEutNgvHaH0TTEdZIahCL++YzXh9o4UJZGI9Tmc4U6fkMqxPHc9MFcDj9NJAnNFcT0Er74bYK
gWGUnNULnUUPMQDH0YCacTVcOOa/PquABjXhE4TOsMgOpoWjs9A93KqSBnW8Iugt22Rr7Qi11d2k
pQ2TrF54AKjOjWsSpOqM4STqJHfEFP98SbTDYf1iRwpstJsVAXeC3Zt6WcDaGn+9n5q9lw74B+YU
ZzZ0EECDhqasa9Y/chS6BnFm7kpv1mpoTI5bpmP2g3K1mRBAkap4Hw/7bEiQbxV2XQu0mglnM27q
ZiqrP5MvADOz2gWmOb7Qx79ilS4yWdpDSyjTHAUn0/a51niHqHFRGQrdvqJA0Xqh6CvBjE4LFYAT
TQRMfROQTti2G0lI//vtCHi9rVm3FSUzU3PHmw1qT6HMqY66VQjA7IfduFaZUAv6SPrjIHjsjUMt
om13kr1/rEEaCzADyoNC1Uam9BUjFdOAqWJM5H3fZlr20MdYEVPMU0qasm94RFu3Ngr/oHP5XOoH
mqH1z0S5u9/cJzL92RVPD7ELYJZHUq0fmlDCLa/+7Yc2Cu4GqAdD5RzPbg+tMK8H3QhArVLDQy0D
yAldsjzh6w7iafONTfrwFYH270yEOfKzEGdPFK1nueOVBKTAv/YoE5kdNPTJZr79tp/ZzBpgsBaB
/oDJzmjbFUwZevzQLtxgOuQuy43n5POqU3sgl46fIcyr6knbR9X3AZMo7AQ3GswI76lbqGGsDNPd
G/nRt8O/X8VZ7TsI1TSPuSoqsvW2sW+C2d4YYs/XpxJPzS6BsjMQnZ0zVwZaPWt9/Aat70PrMRax
5MPudGl1OvtBaAK8LmG5aG5/en79kTtlGU3ZApVhNyX80sm7aIe4z3pCtk6xZHurEYVoBcINrhAk
FJtxWHp2qZ6k1H9sNDRIsOeVerutgbM4F3qH8a8sbkJte0+TZ2SE+wOAIPBVd6krgN7VQJwKws8T
XYYyt3cvutEYgUVu0CoOT5mnOom/t5DH3MGWgafhbtjWPmmDItA4teEREnBJA27kE8hNT5Bpohdj
kZ1QKbCNAIFtruurBqLyhfCE7VgKVMQV9Jz1mI46K+VOzkDVSRRoURwFnoMzfGHs3sH2b5fUlByB
Es5y0ZpQK9fWKBZgYJO7VGOALZZrBgiX6kHou8NAEDVIKvcq7AtsOtWLJeKRafyJp06UnYsAtqGB
vdZXOhc0blFzQHcghmZroBIP6kR7NOgVNyuhPw/ve+xyHdhUB7PxDy6e8d4uqsq/Bk9602y11boK
UR7f2+/6n4M+r3E5OunP8E70efxTgOKXu1mPp1cEIOiq7m+T0/R8P0HFfMMlRNSiL3YdIxhl6Mai
0IcVwPq7DSNZgZm6J2kuNg4GlSybOkhHRBMdpgtCQcIPV1ovqEgfPhBsJNOV1oomhdkXCWbpDUe+
GZNN2Kh1n5XsIFMdLohl+WUQRhu37K9V69CCfqYSOYSsaVOo3lUJ+PeaPfPf/dNSMphCmgPLTIPE
B1TdQzTqsFO6OXrvQ6dG7fVa25qzfSn7hIFukJ6m0Sr2YM5+I4tBrgKk7hXOO1yot4mZfntlQev9
++gF1yM0ysTpCspb5xl6G1FXn0KHl1DzDWmYxC0qBricMdmnwzd3W1KqO5avBDos7XRzQIYJKDg1
mILpaaLv5Wb9VA0jVAwygQ56wh+P44yEWCXVRZuEfgsr9FNg5X2qOPoRLTWt1UdQvK/S819fkJAE
suZ6IIfniMNay2r5o/7h8WdTzmJ5IrF94MlZzELfGU2x/CyK7e65hLXnBK6YXlvsIQnBpjFcuGwK
wABcJvtPXzyooFy6ClC5aBz7uGWua+ytVyqeSAz1T4LED2mJWDTGTer1z20XxJgkmUJ97ZVxwmdQ
YtOFM6rIsLlJMXGo6YuIWL6r3jLhXTU3cLcOtj/5BA+pwdRpX/cgBGIu7NhNBAJFq7M+xmMvvpBI
7ljE8IU5oiZA9n483HN7rjLqbB5ArG3lUlR6WMvO2pf69mU7rzw3rjm1oWNcbMhZNVH8p11sP0Ds
E2oiV7L4iu9AuHD/uYJNRsx631q+V1lrPV4S2t0AtnTUE8aJS8BzoJ3SC7qKF4vQEGrlwoh1/E5P
NHXDGCaSge667TmYzmDPOLf/JWGC91GnowdeOX7QGEpLfqpEKIYCyLZruOp7+yi7rIsLkyZnbxy5
Mh8RpuEhUEaUKtI+7WwsfzWnrcwVUTwPDQhVcUQ/hL5jIHr1sCjrTu6OaqplJFQQqQzC2qqxw19K
rzlLDc5eQ4yhpk3X7Lc0AiSCcFfKuTEO2QnVYQDlXaRsRRQea9DhH3HUHrt3pD6dE7Iu705xDKAq
do4EIKxCTMBEXI9AAU3lMIfgcfuFPvAKwRczz0AGkIrgqxyIchseQTUh3nD1QjDNYCP5vDvjgM+9
4ygGBar4qoqsUgvytccuFVemRyBT07Pi37dGb+/B8FTVP6L9OyVtBSJtZFwalaZvCDcVzbb2bUHm
nc+0Jgj75fhlW2bIi2t1lqYJieqaPPxIsNx5CGi8JhNXCMTmEXgHLlJApMxuJfIzHjCfb+FDVzDZ
Vnrb9watbhXikBvMraMf87k5JD3aJoqFuygXag4JKiv1RImE6TfuVo/qcyKmNniQ9I2F+ZeIkbL8
Wy9SjDOhDEVyRl/kBlKEKGOXPcFS0QgBbmmgXnSQ+WP4O84f6wp3KM/P4QhWjA/yzir7g/hRWPBt
1+nhaZEWujhtBdg+FaiN3xNNCTKpW+QGRqjT0v7pAvGL2+3pQ6ywLYvu6pnht3IHxDj217anMDd0
l60qwP/LzUU1nM470oKHh7foSJBEjXrItvZ4hMSC8N/UaMOV3WU8r1BfJwPwkJrYY+Shqy4+7Q6J
VDqhy0ba4IWMyEpCn1+7TDIws7qioaaDLYHRxL32Fe8PNMkHiR43XzIvNtp5rSp2SsLa1msy7McF
/E9WqH84yNPEa1CsdkzuSXu0LCHFBp95M6WCPDLekUAWxkFAWJuytAp05Gan4H6haYUVHGuYUfq5
7a5LGfQaWzHUhkWO+Nht4k6+qHAEUiCx73CLSgrZsY5bcnIBLe/cMUVZ8nIugefHaCpP0hvzPVy1
beWcBr+v2ZRZdV3JshKo8OaaVfHbBQV1B2/IeszRrbs8UAMWTUS7MabgvkiKsTGW9ZJuxukbR/gu
q2MZ/ugJ6rluGZ02leBLq7oVbreOn632ihE57Ogwd1/KyBFAGyd1A12aqpcKRsY27wCo2rt3cvQo
W/NkTrzAOC1ettZ2dR35/aTBzZANCQXw50etR0h8Px7QCZWGcBkuoVZ9y3/b/TiqIB0COMkZ0S2f
yDVSw5WhGiyzdYV5ZFq7m7NSmxBqiuHcPPU9sWoaDzJJa9cU8ojLWM1NqXFiaAi+4i2SNYRZ2KO3
ypGpuXW8kq+/wtsS4rVF1IRPal7Pvu0VcV37eKhek0+e+4zxbNd+Ikoa+ex6IsUpwvI3bUlngVD0
FMN6954Znl6Q4XAWFI6y1vqUkrjm5jFE16UhdORgdzh95lGkeWzLC8OW1QizpeibMCGtza2pZzKB
xIFI9gSJD/VzMQnweyRwAT6LLBxkdD4Kj8FRH9R3GUrSK1Ztfi9eu9wXP3Rum3fLAtDO4xkwOUZU
Rx2lRMtHjpxrzZtJarQnUCgjONh86lFPVl3Mg1A1PoCE8AJfKQBQ38nvb6tLzQEAkwD1z/5sa7jb
Q4phgpyiiigrw3kiZ6Xq0wTMCe27L2/T7bQI9UYVsCwFc3uTtj1ovGfmbPFqK46YxtenZVLmm6my
wZ0s9qCJHyArmT91/L7Dv7+qk/hBBBQau2zpCdYAHyAqjzLNoqTg8u8XH60/hSbgwExsq9EoCaH5
cxEl4hSk/1hYRwrETHicChZrLpRSICXTZTr874VDGlEb/kDwgO5ihiwdPCvu/QSvo3uBaxV+dnwK
EJ8m8dGmK+9KYAAh3gH8yC+sztOpOtInpfqKS4THk1or/J1DbqdfWAw6PyIs6wAFknJ5OBpYfaYW
96aWp4ui6K56MeRFY8IwGIXX00iH8ON/w0Ujkdb/846xAn/XpPYgbvq1uDDgYew1NCLrjRdBGn88
un44b/0MOzerMF0PeaiJGd+ME5Pf4B/wm167/it1kBwyWxPJE0t0DKl6tsMEK7t59tRVhEPfsVmZ
9+YSWcYGJ3eqda/4DNTe60J0OKgAdeZL7yiGocJb0DJrc6iUCRifR6A5j4bx98PZxZfEWLYR+tbB
Q3OfwdxOfN6F8fJ0D5BNZMvBQycF8MSTkfpmf1s9Pir55Hsj0aa04LLjHjiR0NS4DABIhNeKJ7a8
LJrdym+gEBx8ny60S3yNnW84M/rBLD9SeEO0+mTswcFBr84827OKRboOFgkS/Xi34orqYO8lbxWD
zEbTK0Uh9U25hsmKrbUstYHLZxwQPNSRljwZjc/SYn2N4bxmthhTCCN+cqSf3khFBVJvJ/b9KnV8
AdK/Sq/Me7X4Voc0vwwedpe/M+JdWaqdli0U1UgWV2Z1LpbacD5PjMPOY4pLmTMJX6qmIe0r5pWT
xkVsTm1KC6hL1XHZTJzMJXFrbipBDP++Lip1Jt8ksh8tUjJDauZGlXXjiann63R5Xf9nCdYEMeL5
4V8ULDoyq8ETKVmT/t2Gc6gBGB9EyjENJUMVBFZTwtEugqqJpWTbbtan+RubXPGTX90ToryDKr0z
wjCOMom2Nu42em+mcN/jCOm27pIwgOOtPLESROK9L80i42L5JT5lVI/XXhDb9arJGSgFXlvuKLhj
e8CuuYjnaIaGxSexQc5tCi4xjWe1a5ytAxMktqm4ti8Cmwm19tZISKM4493oAghpr8fz5i+R2TtK
kWYB5BNyoijNDWxvnAv2DRkVOfMN9gYa9PmwayvIEmI4xkbdgZD6pV6eEa2EWnQAA4hS7PxCtsLv
geIvrp9mb/Mq3V6ZkMVsmA1KIeXTyxswScIsQhqwwgiiNaos/e3XR0X2va+QmPbPJV9t2s4vPfGB
z2I0gLAQi0tUE5E+iMIfjY2zuR8esc7LyfdvfxjEVHPOJ5jm2vAsqd8Sjo2aaOmZTVg7Hp8JCrn+
peM15D2CDol7o0lCZdH9uDef4B2Zfa5t8Rs/lRCCjkwXPQF/Gs4fO6yzakeLkKMGeIUq/dMaArFQ
PQ8hu3URYSIxKxAniWCDwecFOFBLsk6exP3LrId/XYfiD5YnNrQCkEIoJVo671PfBZuSOHoiMf3T
sYDbY3CPBbv7JH0RZRXihuoyXYHtlK5+jmmaAf+nKZT/Ndb1Pndgyi6JTOJhb4BLheE1J3ealJID
umPxCEBVoIcfHS/71hKb7FHwPRC38fBHNyxv3bcQF1Q0ILHIL1MJ4g9QMTw+kPYkRHc6TFEWCmwX
F145j5Cicpu2UAzbhYJhRuac1hM1Tbob23H+MAQ9B11NXOeyFvuiMHGlMXAacIA3NFWQ7wLsZIai
qhe5YfP2kQvisEPhq4KbXRRCKU7u+2su1iN0djhGgXIlf6ZGuE3BmtItUEgI21yaINCcg/vppeNz
K+3eZN7tE/VZh52MiSu1baKlDobgJ5mQ9qGG8QJsduNNXUnQFGBX/fC03LlO8WOBIMZ7JwzcXPnE
Oo1Tp0//QPP9ANQX4wRDS4iNPuWvE8OjR7vmSL16PUmSGCrR5IRurf4zorxbCil9/j4FGJjPgqnO
45iU78hsC8q3OWRoDqYfrlSzEPl6v2rJEGE/7gAM7X52zsCBzV3UB/awPDKQQcyEo8QcGO/BIT/y
bkiFD5SF21GO3pNW/Ooj0PvU/m1IGh2Hr9aVDI/bWgUB1Gh2iOeBDfO/hX4G1gnKeCLQMw6M0AYG
oXFWYjKkYL9jrbw+KQvAYZ0SblnY/2M6BvErzU9gfyifS4dRCd8As0Il/SRjilbLn7dH/6DS4kd3
46ibDWfLjwjqJ/I1BVbRGRmZ/EFaRFPaQ+qDYGsVX3NZAmZ1lXYAhc8lLb9/Hemrhc8GzyyVtZkJ
TNrvlScoYcPCkrEBo+3BoEzcFJ0KCml0Q8a3bZsqHbWEPYyYrYZ8TWJ+fXZLJAclfdPsjRgp+Vyr
DhXXOcw6FZ+WwCX/csooXtsVxMTiQXDjjkz31LQTiMHhCiwYTlta7kFjaD6QJzZvUXlvREZlb7zY
eZi79645M0luYXkiOepndlfef+QJ92/o13g8XeDNLoyxQJeqwbSrTnDJSqN1nxylHRC2TwHMCdv0
fp4eI7nwC8Z8OrirkDAm4TPHmOlzoUPKtkRhr6qNogKUHiQugRrtYj8AHTJnamfD//JIIIBAfUyP
JIHocTIqbc4bIv0OrOY1HjAHH0NGKpYVnckAngfEMn+qMTQYq5CoFzYchhIkeFGOiNGJpVcONHYX
faPfH74GvhDlh01GkvFmxcMYgc6ezkjtw7qMo3+7fMzbVVeuLSa3zsc7nmlV7ck62o/fAiJdxf9t
HlHjgn2bSwnccz46ibORvDTlNWDIrOc34W+PtnFiK7eKL0dmqHG7H6rQGVSZwPYTAF7rCc4kAlPf
/u4TjbKkQj5o6LtftmO/1yV5O4yA5UGnrHqGd8KYxxxqaOHhl1Qyev+Pq7gahNBYIIZlMi49sv3c
ypt2O77xvE8eOs7buHSnIYKp1xIOcuLaFkcT3upLck6onP4q16bp6gRFiq774zQh3YJ8EwDHejvx
h1syIGZwlk0YY6TnntCj0QgmqWbx2GlFHn2ittAVlu2FPMphU3XnZICzwMYzVscKmaeDKBbbWJfB
uZuuPvohViEQ6gP41fZBm+ZLayvDMuTv1y1dCQkWI+tZIw8myWCHWAQOQyMkzbl/5ANmsCNk3BPC
2FtpDZgnSlTCQfIaHcXa19oqPpwj7zZTuNd/R8bwBZ+JRsywyDBHeZowC1Tz83ZQRN5eOjiJH9B0
RsasWCbsnUPsLilxMG094sF+QVWkHw/ODU0EBoy/PrmySj8QK+ilBR4vpkRhBU8Spg6cx8EPbLLN
lCoBpR4EKlWYfNMjxvfea76Jjx8MORWa6RWYrUNV3qXibMSPpAcGNDlUoFrBYQRrx0MgOZ7nHKoI
yRrU7/ulcH7BICL4LjXGYdQDK8UrLIygJZweH97+T1xAIcnlgCIcnen1ZJZJf0uGWzeI/AUbA2hi
RB937nBvT1nbx7iLTsrmTuOpNmUKEvgrly4KUAM33ulI7YQzlBFOzSxcIqkhmokemcrdz6vAomWb
4wPkwsW5BUcEotgDSeFj2apb9ePpGgdpKb8RAgr8TSDZbcpaSB/ym8Ph1SCo2YVUanAIeHwLo5E4
hTU+bsJlwCZv9rQFBDqtq7u5D6xKtj16uyaJ7W+fjUgZjQqmdcH/vaSxS42XOkm/N+p2oCqKJefr
x58h9YLn5JEsowT+u3Y3aP7inyv40sKwuhir8iuL8/np1TXu5tYnFNtArurp2vBpClII+Y+FfkOp
ZATlXc9Z4ULgmaVfDKOK8XL7XM60UdGQ+cTOqkKv9KTVJUhtJJQd1SAlVVktws3e0jIw2xmpx9Y/
2XO4qDkb5vPWNzbIgtv7k8XOBiy1DZ09CYnBfsA830Y2YPLIz0iPpO/GfroXJmleXevUqTv7+SKs
yfU8OIDjtcYtsDDFTMBLrMb+1U9JwDVnewTmUAVRBYUbUAuM4m2ewIL9XMb/TUXtr/FU9Y20cAJy
ks6kCGPEXOyJA39Pnl/JSEIlU+GHmv2xmXIRkXV0XfgMuegV/+h8FBtSwGTtp8tf9y0Xu/Fnl7lN
2Qyn1f5AbE8db4ZAmHBejKT0eql9XP4G7pMWUw4Oa2FK8zsjx7J8PUeR7RGqgW4FF5/NCdz+ubJn
EukVuM/ACi7u6qb1h5J4jVzTLVETrGOu0pxliVx/5H6P6OVyvar5E8DsgZpuSZlFjWfhjWP0/tqC
wz+80+BjJ9ibr8Ty+nlrrYAkAX5J0X98E2pMac5sISD+EJGCm/YIMmlGO8O73jnMzbzg78+MzQGl
FS6MaFDeW8ixu4OB0lQ3p4qpLWaJkXLfI9ggZOoqb8nEUcovHxc8i+keAqNaYmZ/lUyospyyv1pY
wLlx+xkAzfUcdBR+6undDdqgMsBNLyr6xjzK74sAoOhY6OHxdZnOoOng9CzTSgh+TKRZWkGEuQt/
1KJwRYty2dWFFicWSI2WBWMvZRKVdYnjiDwHBlspMhztPeJRld5g3nGR2V3smGPHiEsWTEHbS3O4
osy3oTnwX0KcPYbEcVe3OGgOUnSxwcLeNSRfT9Oju9IHlN6/XsiPFJD/rwlrBfMoaIRsMWJzbY4L
qnkAKLXX//TfoXF6o5dwRKtcMorosYXfBfTg/iLJFI3DtlM07dOCLWBdLYKMbfiFbK9t00AhaUpv
z/yziOC97xLhZvn9MjSLMMCG1Wf8uCZ54Ryq+c+HMXRfMeLYlhK+2yXa/n8Skbsr2VS4fa0rHhAs
wlxfkNtjLJ83qrBcGasDQzRAW4NODCWPE1T3JFz7+x0SB7FZM+BxfWWUA01mEdX/apcP6F/ZuJkI
ghIO1WMyVVEKtNhgZt/KzzrpfjIpeAUgqr5mx+wg9mP3tbuZc6pPmHo5PQIph6X3yHFfK8cVG6bD
Xr2341yBPhxttG7UuH32oyOB0BCdtjiDIDyjMsCrp2AS1oba8a+3GAvpmzmSh8N9nHU1BIqs+iYC
CnOg/Gl7LkmqQR7W4Q2fX7pcAip12wsiP4uX+ynlO0ZhnrVvgsJeUCyqs+dZJe5N2WDNQ47btym9
3feF7apRE1oxYf+VDwLpTPfU+UgEg1U2AWE+iOKFCAqsEG/EMlUA58bdODBwTKefbVReu0W7v7Yd
LCJjqawi4E3vBjJJpap1o4cgCS0TwptjgA1ykfQUS0s7S3hRkcPTs4ak8c2eS4opqwTCDSLErgvs
SNtLFdFRmsWvyr/Dkp/jeNwNJlfETIJONMsHhJZ6S7VzaU59HGPBeXfBEu1ENt/rPAIn+Xo7KzWv
HjW47yKdaqM00g0jfCuMAMpdnefpvfJmksMBgMEtFXPAGSk99RToC/smmr+2isAhUa455m5xxbNc
FGXmfiWtKq4XQ6SfZniWBjDbiZpXcnQ9Z/uTRwiODhq4fmXVwQZid4LWmHRguNNqY+heMT1BD4z7
YsZqaaF8N6FzVssVe+ofuZYRtyyJQUa35OgvPzm4T6zepl6svRtboFZ+AfEJoignBYNhdwwUtn4j
B31B/DofLiYF3SsqvUVpyOmzhe7llRiKFohtszvWPaJbl0OtcWCnarnc9FSMSH0kq3b1Qc9s9xds
z/Htm5q3oelRayUX4dS49cAV2Adn7wMahgLbe0fwyI9QQ9X/mD0SwvV8Djuwjbt7nRGL69H8Ial9
89T+BYUalYagJNFoRrcLJlzEhyCLLtREZPl9Uaeom3Vd3MLls2oxshK6Deq3zsLf0gaPstks+xk5
D4Bm2KTib36gSFhkr4FO8pvs2pVMrirf2+8B3QgDFUcw5QReQowEfGWkxrqYahOsj9dUzFeI3+kA
ce1GPb2cjE/uZSp05szOgEk/MzJLErwjr3ugP9Hox18IfUb/+TAxRK+wOqaZKOAeL60gsqxtwJbq
evofr6llI5BNKGTKp4NVBlXSytJDWZQBMy7y/N/LkUfXnWJiZ73+5MgvVlyICnD7oR7Ha4lpIIDP
0D3+3+EBOZgTUJbsPqbX/JLcO7IcMJH//OERvSuYeWoJsq3ih/dm7U/McZNkpilFpE2vfxeIHyN6
jCasP2MJK1JCoH3BaqNObQZmn8M1fN0ZJjieWmAA1xfLVyxveZvqEqo3iLV6DTGQOGW/AdsmMFOp
/zUJZVXV8DstG11Gle8WfXILFNlXShOWpTvOaOZgl3pYmM8Kmk87GKL9JZ5MxZr7r+kn14wd1lSg
7DhVzF2Tvx0zvnIv9McKn+t3Q1LsMpkZDkbiRtgy+C37qbtcd3Ev9b06LN6Ia2wFwtoOjJcgdI8a
epxoYdY/za6TsmmvBWSS7B3OQZrlHZWqcv0xMBEi2yQJXXhGFSVhM7uZ3kqNu8EshqIluxXqYwrn
rnztjllufP5eqw9XqOA6NQmig4+YTVfVZS+3s224vKiZbueUZ0VSdzFVwh2oher5TkwS99tjm4Jm
CTavDufK5E0HrnCxHdUgOnJfaUSf7xP87mLfYDhM5yQ/pZuwDcm0oEQh73zaWrjm6rM4Lbq4Z605
FWFWzbMVq236gO9lqQ+Dw7DB1BgB3IIGAx/N2nxjdx/Fu6MBoWBtf2ASAKVoUm7wa+4gJIf1g5A6
ruw7XEB2sxZ3aW+FoP2u5bYz+bX6QPjzK6qWnvVjYKXN0iAG22eDCT+Dnfe/+HGZxMxSF3gq3Ud8
E0pM7YnTgEUA+l9gin+8lftBsgwOuCzwgba5yH3chKfVhPtgh/bf9u+rPbrZ5C9XIUdq2SIIx1y+
wZyBJsQ/rLKXmZtDfu9neLCYMhjw5LQNd135UlSBF9PErm/prp1GoP66axUXtPa3SqFLYXE3DDTm
JUnz++Q6mZGcGl0RG88HXzKZ+0orcnxi4jU7WfDtZwbYS3koWFs6+ZDnkN5kUGexbGOuMFn65pzM
Myb654wwVaBtstkbcrDiTF3CXBj+UxSl6XkXx8q8yJh6KuTprdVNddOZz0oxRkKzNlde0t2GPBT3
QOkbgIL9Za5lQ6QrvqxeJUMAu53Q8lPwewXeXLX8CSQwC+ffqsANayBclOxOTipHfaHYhGs3hjRu
6SevLHAeAefFw43Y5SFLzMBC+aWLf4JLZGg//XDUqoLE9mtIGTgnol0ZOP6QoUGKASoEEGr/FAdd
opTXVxXEgP4mx1+vAT3WiXUQBi8pVEPt9RKL8gW/nH27p0Wl3RYBQVzDpUcEmf+NWJxM2L08QWhP
8lqD+F1j/5Vx0XLiRFmutIacJ1C+HmKJfCyEdM4O1CGLyNZQIqDWpmpF28AvLCGOzvrX8664yAXK
CTPQBKmJQTYfNuorDkZWyGh7ULS1SWMAvK1lFXo8ahk9YLBvUQ4133QnoUjTRvkiOreDMjnjvkYl
j8HltBT10rBj8aG+GmpBmoixmTcxyXVWE2349bmLe3MGXsdkAr4+mq8j9zthhHCUcGxGwr2VD+6+
cCwoyuRDY0u/f2aANkkLB+IJZWWarvurIamopPONxEGzXnQrRcpNjdSm/C2hfq/ezM4w6qL8QcBu
HPp0Ku23PenUeDWSodxmxuZmT320uREWo0lgneJF4qACwWnVi/sFn0sFFzkEbltHzWSohX8eHhzJ
R7MRym0x3+NGzIL9J6Wyw/BylWs1v5ZoQqMs2cbhNmWrigvxbbGsyC4f48YuCO7592bDDJW2TBdN
coEmX8AQ/lDstrpewntx5RkYmuOCrv1uY0AttRg2hEfkeu4NgdShgfIxuX2rc2+i834/zFPHxxFg
QB1fp3k/EaAV5B36TtpZMenCZHoyf9I8z+0zpAQtPyyLJzGi5CkYPuoKbnLzl/Qu74fhvqQmAf2J
H9zTvjp1hSwk0HOSkW/HMPTSJlNnQVaZZUHxu1UCLn5sntvWF6e2be72l18I5jnPPkJXd2KPRR8j
EeJtFSPLzgfcWMXhQ/Jyp7QexQJDrbfZtXGlAuTiTQyaICbRUTZ35pckgkolcuu9hy1PWvkYScMR
TOq9ody6j3DrQh9owuZ43lJOg5ib+Qm825XJ+u7nS7k4vKcs1yta4EwB74hsF2uhGE08l1zo6tK8
iXb21fPUNUS4u6FpNgrkXDaGigzj20sn9S31xBlBM4gyBoI9F21wGw/DvnNf/xegjNU5ygQ38SRe
n0ln2hoaHS0ctpv7GpLmApl2zBkPWTKp/erzTQg5Tdngy9qkz23H0Mg/hXWPk/u1WgwCY55mFKC0
42gqpPVRT8/DHoDzCXfpI+BpxjepReicxtb//ET9BmYsqpzmo9yVrJDJufgJT+8/b9/vVr5rhm58
3ZPYq1/xs0YjpnIDAtC5GW+gvPSuXKhQDlOz+pJp2odJ/VfcsXWWk73NmNx/fdymIxDOshKiQ3NJ
I0Oy3QE4EI+ucIA/z6Jso4zLpbCB/OluVDo4TDWPn+IMayraPIyiXU9qrAECOcM0giUhTjixOPqB
iQ4MEPLzux4TZ8+MxyhGuWZRnX9bfK1by3dyaRnoHOXlNfc0jEZEyq740TQXkivDOlzhzHFgreOg
1+m729uJQTkMm6vA8+RtrDHAWjQDP+elgSO3M6BXdT9F+Dx2q8S0foP2qW50sY1VPRxkV4wSBUGs
60clYcS+0L1VQ0tk9Ll+juWq9QwnED0uYciNDfpHURfqi9M8e7ODqPAVhIo4S+PGaUZtX6MCd9p3
eRMEsCW/7K9o61zbqpQDkXjg3fwxkrWfgjEPzrOaH030qhZSTIb1P4Shwq1+HLIb8LnYoc68QVND
Sf9UeaNpIMYiLcRyk8lBN5bnbaZMrRWjfDoiWegDadrpAASpVG3UKEaBSzLojBk784elGGJGV3Kb
5XAB9dwLEORhxAyQ4JWqCx/DoGpHKmq4jZw2LM2e0GFx0+OEv6ExmLWlBP2b0HzWFTePNv1B10AP
584izRDJMz0P3JEhnbyJO4Y60MI9L2+YGE/IQkI30blhCyJXqt6WLgBDWRx2RPiJoZq+X9jo0CKU
JN1lGLQ8S8E2JJGPOsfwOf/sxzQ1Q0aWpLfp3tdd+1r7MnlMqHG1jiu7c2SI1rsBdOz9Ih6rsbo/
FMQ7/C1QU9VfhkRNY8/qda1nP/t9r0/0PnZOfp52VjPShcaQzCqkJZ4QNI7hlzNWPXP1+TK91UMw
mYlzMhYSi9zDOM8h4YDfgP4j0jFFxvVakr0NPMKNaL3xqFJ6VcYJVS4FrxMtFMnCylBIVcDnS0Vh
CghiNTgPrsOjC49SR0u9elnvvDIcfMJ5EvBxxQ5s8Z68S4bezEr1GqQyn/mUlVtTlQ9LREGDxk3G
tT1gK59yGjho84VR0na36DuUmpret3XerVEG0FL7TH3ykjQlnA74mPTzrV/NNiZMyeAx/pMNT5Jn
BjBlUdqF1fTTSMOTwwfSQhI+SXY3pNYjeB5Oj724N39gFFYsAsMQg0rTuNtFAM4n5XJgJ7ZaVXTK
DLGBf5Q9Ub8kAmzlErroIPMMefJq3IRnFS7EqlzNcwPFGxOaHm+WOFgsiaBcvO1pjVwC0yJyZNwe
WxJ3k0K4La+MAczOw20GdYK/X7/DxdfjepiiednYfiZeZRR9++CJtQoxBrfWHdfe1++mCWcVx1Q7
lhZQDj4ygfggjmFHWVQjBim0GL+LiTXe7JcnO3VOIj3aPVbcVu9vVymvGYadsHPGkGjkWzURrt3K
D8UuZ6sI5AAg08QzE6Y1f9YhWhg3y87klejUKALHp9G/1zdC+tOqzp7zXb0qXsGjTwGeFpS7we2s
UIJ2tmb+dzcPhTX4VX3ye7ejDoCYhdogfHQzWEJpTRUz6e1DzhI3fzgd8b/5QRG3B0dpgmCyDNAC
iKybDlGGOvh62ayGNasFIIyrSo1FytLcw9mJyi8R/NYeW0gIsqfareM4GuBz1DO6sjd4z2lk2Rpa
xRUchFsc/0JqfvvMRKXtcczGvJvUv1BFAkvXV1CzezLpUhBQmGw7WdINXX7MID2OGUqUzRnKH+tC
KOju6ieA+yW/GrAGEGEkDJ5FhWyTsEx+7lwTisfcpu4KvYcNZVe9uW9j/L6XvhFb6uwQFTi27PIs
+JSRcFATgO9rYdW9TVehbNiOPjK03xm3PhiCcXSRJXFIKSl/jmP/zXdqC5XsJg64x3ggTRf3rew0
xT4M3oeEuAAEySwIDsjWQKYOTWmm9cYwR54m4N6ZT9dTAEC3rS/n+YtfQ4AYwGMTm0Ceo1YR/57q
vuw4g/1hPk2Qx8RjeVpwS9aWp3rX5nTYtpUOM8+j3qWg8+IG1gyvAg45kCLKczYJwqn7WtiV8241
K3RTahWOIHKUSiuO7z9tolNYQT3Ory9Mwa9Uq6gRe1CKKMelnVR34jsDkB3qjCLVqYjhKy48qyy2
QwceOR/jt8Tdi/EuU8XVYHNU6HO0O9vGmjN7YeMf/tdbxFSLRNaWJeg3XuDdyNYh5OU3amQO/knm
AuZuTsjApJldRRyuB+/3nPyXAfgssfr14j7P+L4AMO6tmDih1mhoSekQVBf02D7XUhH9msXL4/fu
6kB3QxFHitRu1LYR2JoRJdHI8yMSjqXapsRBh+po8ZwyvjArrWz5Ij7DsT2sP2hynkTwYpS6Zim9
8J6IoeTA0hgb35xdK4c7SwSSaegoucI05AWanodUwIHWAoee6RR5TJIuogZ1cVHNttz0LOwGjg83
ypj6YGBT18hsSxTjGygkZJaW9zJN4i/LV2fqCH4pzZnA/u6D4McAsLv4n1NEJbgJd9oKUcdN20yr
z3bCsgD8P/8IZ839JJnEA6qhJtvYcWnS8RsiAnG6bnl4XSwS8jFhg7pAhV01/roa7lilNAuYDG8f
JFeV28LgRfiCzeAcasfy6I45eYF3snAFFtl/qCj4tqpUYeiZWdbzuMpcQh/uOM7LsclxjpS1BMMG
qJLVZn3nGljMQVssvLBBQIcFK9hbDbVO+xj62zrXhL8Bm0EWbeDn6HJwU28DT8FAyJeLZKQiCuLK
qWRbsuYobyFnrpdD65T+KLUidd8lx4+620CsiecDGz/M9TBYkGx+NlFItuzPu3AjGCXSjC0T9ca4
oEXtmOyJwXfeXyeGqiH8bucjQ06zW7YDWpAM6lJTIxNLDoQXcXn+4E70jJMoM2gkPbJZ9dI5zRdY
wFK44s8h8W9FWdFklTlnM527rj3q+LxdCnhZBgmlxwWgdo6ZJYEH8MVLXeLXTWwUM/asGGqOK3jz
2QsD+GFJAOMM5Tnt7gNtTW7oBbQLbAW4+GPk16tKGjM7rjq00HNWRJAWCz0nBTbJ5vH9i1klkW47
qBQpmqaep2O68DPq+Fmm+tktQuG+BpgxUDdS2IOjWmbfjwV52ZcphQ4xlTcvBajCrXx73URZ4TVL
/HFKx0w0do7bWfktxK6xHukoJA/pBjSmZyjXgL/ReiIxkef8USujTuQjVurcMgAxcB39UIx8PTGb
3BKsmnAa0AXQndg5FmDXBe7P38RikdNvcY6jfkoNstb6gUstchcqsX4UXUGLm7IesczrFhE5dsed
W4OnwiuxwK78sl+BatSDZLRrx8FsF8bd4rpZ1uIvlFl8Fh8XtnhqUDgBSAqU9LMAuYCxVkoIbcYw
eofA1bPgD52SAM0sPWw+k/IliWG9I8tDr3lPoOfDkib3UtbkOBkZ6XgC/6Wf5o1tIeH6KewCdMtH
n0LvjvIY2b10NrI//V1go9IJ//npzCz8kEVyG+4UiiK9DsOwmDvLvsI216M8OV97iz3zQkW2+OYF
JW5yf+DJCHiqJKoUD3v02aQmSPXTHiP+WFKPyo227SlVw3HbqHQsZWwGVn3lXv+M1j9MmqYNYBDp
eqgFlH/iKhYwlM1L3f0QUNrx5sM35SVppQ36H/uqMCNCfdMmLxIcDICZivmGBujzwis4/uOzkbTE
NN9dS9yNFquxtr2ys1v3zu8IAEVpfPMbLALqQl5nHGOepbfoV6dDvhekx2MgrVvMO8VdT8mq384L
m2TzjuCtkZ1ok7JaHTl9lHOfq+pJ+azdYSWppnA0qd5CYOvT/KemAMqzbxKcPCZA/AxyDcqdeGwd
Izva6sjByX0ENZifJXaC27uSnI3W71MKUkW3Q5wpbivs7H+lFe74vk/EeE/e2tFt8erD9KYustif
xP6IB/q/psTjN9FH5uSkZKAAZAf8D2IRZggAt7BpNzWNZ19ISUDT+JYBOvREM1kb80Z8xwVhtXgU
a6JweS4ibD31GqTxgQqZQvFt/sXaT+YvNgAaLrehxIATbu37COvdS1PG4gJ8R1FLjZIzBHRklDMC
m0p2cXgzIpMCqOra3TcucPdmQMxrKL8Q8ghP92MHYWsre3q718bqP6e6BqWsr69AEsoct/K63bFK
GE4cBOkrnEqlp0hMLZ5fqktVfyP9kryhRpYx6/jNSUapf/O8XfSeqh8Tob8HbuCCzw7tEAC9JM1U
AD4H5D79E5EedcBSrNFTvNvE8FI+9CZkkEVITNi8pxVRX8iBBM7YqR9JEIg1Vq2rT4xO6vW7wvBo
G9J3jNdiRyuUlTD3rCO9aZgiUnuJbqrb50r32yhKy6m1argPdV7rkPbJbwr84jrzhEzia4Jsy37y
ZSItQfyEaujGFxcQb9r1zEPW/vmNOpf73fZhOGx81j0G1wOH0/gO/xQdFDcvrTSfw8NVsi2WpY6K
tYLaYfOFWbyUnAhiC6/yY55/8MVM7eCclFzNKHlBt8xBq9mnE2qMgH8YD6hzcVXtPZ8Xr2yh3Zi/
h535pcfVmAu93vNvR6NuYZO5ozhxOz6alnhN3QEuV9b3soCTiIFYAfeRmk/RvACtTULETaY9EBkk
mJDzWERRGFvluiLe+8EF6BQmWxuUZgd4uACLsj7S+HpJ+TTfwI6/S1h4FzKDSsaKVMy1AcufuELf
uP2FhYV4u6gM22CUMyIuIzQI17I+9YZv8O6/LIqiqntPMZFs+S+j91BMOZMFm1oO8zhgBmgwy3r7
PvN4G+BLQfpQOhtMLbsY4cj74FQY/16oP63WYcs8drc1IDhgcjogaeleNyBoNzLJDxR9qAPdbYSS
XQ+nC1KrFdIsMHcYovv+V0rwk4roEnV1SsEjuiOKDZU4vGnz97eZzQIYDmcugvAWoBzCYKSTDGMk
Ywj5M/I6citeHHbIRvuML3lNaFipGDHND0XaZbZ56dtgQ+RXVM1DYHYuHb2HWXeD93UMajAIr+3j
ATPaPZshJ+7myTzqoYotqGI1qSksIZwEMKqf3HrEWNFF2td4a5K0xm2YMDFLkUyLuTCg/kxot7jF
qrHJez5G/H21CjlXDGlyI+joAzY3wAb/SOHdnmN1Lmz9PD1+opvBYUJbUt/p8phq+2TzJqUq+/9L
dYyJDXN5pr9zti0RX+O6AVlW3wa3pQPeObyCNSmiShVYFsCRy8/v1W6ex9mrnoCdw7fd03z0o526
tK34eSY+YdDIEiMVEpT4B+rzHXYUTaWkKy7GQXGgYn9l3WEKHUdxErW1Msgy8SLjHtxcO/8Xemuh
uxEP65Xo6KwrMtySPVByYu8UG3Vf/aU6WpWRO3NZTgYaj68dT5ausTmHEcbowi6aUjJ7cW6XrhRW
3BOg99RWELBNj0egAnxI0vFJ+od9JXbXXTG2BHw7SF9UXtRar4eTYoX1RISQ9LYeQ6ShMFAfXKI4
VbMEclyPIeRSztImtZ3+AHNO+74StFl0wILpcgTCdeSVBr8u/KfVYbqnD2o4s0kvmPe8dBqbGzBz
lBxsUJtiaqA5F8t66pIOv62cY6LshfYwlrYRI6kPUkrPZtCEdKTrus5A3YN329EKFFlgYKqcHWbQ
4UBmN8AurK+Rn+LLXIWskF3jGPmg/Z0KCUnr0CfBs6Et7T4Osft4KR8/vmrxHRT/C091IxYBSXFY
j4RQZPu3N7yPWxmGlvYLYpcFXtFrheHreuVYDE3QCvEMOu2YLVHyoDHR1Da7lymtWKFZ5wECpz08
n8m/UBg/0nNndNwSrwYeGemwai4lxzbA/5v5WmkbLC+/EC0KDO3Uh8RefK+0s0kAQSqe+gUJ9w/c
vLtGUC1/V5OQhgCOsLWGeHdtm9O/Wv21qY0z7HS7yL7aqIl98ToM+TEfN4RYFHdZjj1Qx7X2pRPO
Yc2XEJLO15GcTCW/x+F+lsMrLjVirEYQ5gcunhN981C/YEIGxz38qszYsa2H6r59QWMH2rj4SUXX
osif0hSHymvRmDfaCbqoPjJwMDxW34HOzLuYAH8XOVqK7lagQFCBh7NynmZupGaU75fonD1r62lU
A43SEHGHdGVuQmaoB7tfeib9//j7WV+eCBwZBvDILPvYumVy1VvtPiG4u6uA4Ygm5Jo5AxxGjDGe
Xx1BzcqZ7HQ0SunNnXLMKFXquP4Nv3a0WUM7qcn8h5PaXhG8xwx5eUw1HWUQ87azmO/IPzBgL3Vh
qRjLL20HHt+0nwvjDl0pm8+IclbfbF0c3Y5OgF0vQCl7LnXGNvoSLsnVSsT9MUNDA8B/Ru+SZpLm
+dgLEc3DAV37XM6WcTYRy9k1RcIyOFIcnSMlch/Y3MHumgioE+6Hg5lCE4YGFyneToLirqfTO5pm
OP9f2Efjdx02UfBQRGKeI2YwWBjmpOLiPs8nmyEdSZ2vcr48FI8AyZUOgz9s4VY11/6rVvEg3RvJ
SUQb1Rg88Ck1KtgPHHyLVsFZp1aRPoIPYQKFI6rjBYEDUfkAxO78Zjc3D35mYkdvt7K/gls09wKr
nOM1w6fQGLSctwbPztiNiIcUOm2wzsHotDgRyYGC7LoNHQep22i9B3qdAjE97W0Gzn4N3aFsW+Zp
pXwpTy8VPQIvax5IKOub+IApnvrI+63sZPmAQiQhfjh4J5tOVJMrICOeDCoW7F4DiBPnP2byYUe/
GXCIItznOybwMWIAxyMXX9PXMTya7hAoIPwjFO6e3Zkbqw4W/h8H+MpwJnxfVK3GJF0yxeG/m0AE
pqSSkgyfvLEwo9JmspAAnib+KxYYggaDbIQHa1MU4lxo5VkgJr4pGWkupc4i9WA7MZmou7QUBzq7
ZganO8AqEO4T0RssGtxnGAcVhAzboi91tZ4lrKKSgGFMRVvRvE5tNcYQ90ElepNmN6HxTeODi1pv
4weVlIlLQMyLuay5WVttq8F7w575oMlV+m+sEtfG3cjYwrotblnhijV1izHUVxFOddxOaomCFHae
++GXvV/rDXBvPbjdbCht1l6v5jMCNDsEtgbHy0lty2WV1Rl4zqztD1kqsF30Fa25dPoelE49ssnk
qS4JYHk6JMd+bNKoah5V6nq1tdvyEaXgeYaCImOA/y4kt5Y0bGYQmynKWAUgk2Jde/DounoS89gy
y1lDSTU6Eb670e/b1OecIkVR5VD56jVv/pbw4g53WIHHCLz0MrmhDmxJzab14WfejXW4LXgwmTl9
OkyQOPRKajIOWOO/Xml/tCaFtneobztxkAT2Ii6lPxZoDS+dRJSH6Wd2Raf0mySDddtzPyYaqZQB
uUlXH6oLiztAnJq65TuQcnmbtwoaUykK8U19p7tJGdkxGgclz2rWw6W42fF5JBOpOQ437i2YFd+j
mKAffnifjW17QIyAvQVk02SL7+7PtPtS1IeSUcvu+tn08UP4kChaKpC+Nk3f9+2Oe/YOIzW+Itm2
67nXSx7bRkgnYVC6UPd8rDfHSXWOjt1VMXjUItQBB8EpL9cNF4wYO96IwrIJts1TpxhEhMy7r2xC
762NqA4UgQhhnzzQVsQkYJU4OoJaY3d5WPTgW7XBnxmuPFKiD3kUVDt2pjVCS8B+nfk6BWv0ivzP
OFzzgW0GVxyr2d0WQIesIa/u/cuRtS0l1PS/WnZtMs1kskFXjBJ8itzdyUgqmSbSl2QIQcJaNWqR
gaFCzBIqQg6mFv44iQH3DhFFW2vsya019g0Y06s+wo+e0RdG3CAbIYsuMYs50Tduqqv0/J7BI9Te
+pQxmUl0ZJmsrEYcALnyBVnhSsJnWKSYfSrUyB7wAf5FMkzpC11t2eBIHAxIlQx48ZiP7emQfF4V
A+NNk8B3yPjv6j2DkrMWHssuiZeVEE1J50h2PwKVyuhyzaBF4YLocEZ6Cchcp5k0FSI6MyEz5eiz
k8WFpY4wS/H5leaa9kbAWiL7Zz9wLZa11NRyMzAjsbdarD9IaGnvJaEzQDgZFs3PWaNvLmC7Dftl
YgJnnfOXT3e/FcGgnJ1ifuga0PIRJbGas42KSPWoKmPLJ3Y/nvj5v1Aj6zpKEq708gDgaOsIT65E
yb408zGsSJuJqeoTdJOz8wI8IMY/HDHjcJ63kiOEHQHtLW1EzLgVIddDNlWL/dcfKkmB0RCoA2hy
5g2KKNtIFOot8gJ7dz+BYBMAsfXiGRrpIQqAtv9pc83ahdpMMUSruqlbtr0yAxCoYkHXnG+CONuN
WPxSqSNJSai070rqEYqRKYhF17rcoJchF07026CbSiHm5NvbRVwSkAFQMnu3DzjcibIY46Jmq1lk
Ba/Wj/U3pPFgUQ8r1ec7iTeUxnwdbn0ze/I6miYRz48J5Zxdq9umgb+KQCIE8fNa3wO1RvwjR/8m
L9zZ5Ad0xwCXAETzrAAPEpKkE/w+JG7ROD7zjlyCdTXHttpXBfaWTrarHGstB+QrHVslulFAfvgs
g1Z2sDHBu4TphD7iDlUjlGVvLWLm32Cb2xrNcHm+2uXtp7ku4CzSAeq97V0XF/EA+DHkSD32XwXc
LdvgmDuCprCCb/o0tE+OsIMUCBk7i//tgKl4pmo4VAsUUDZzDr2wwUa1tZeSoPT9ByFzEU1Qe4DL
ccgFppQAMf9Vs4E/PmGOpIzsB1S0oe/+jZ0XaknGCBy6YpSTHIRx0U78W/T1/0D4+ZJED+k6t2Kw
Z85EfrlY6kH6faJFtlEwyFgZib9QbRYoEOmdP4kJMcWi2U/X2cTKoih/A2cLekIMfvboHVKgWa3Z
lp+8NWt16dfAbA1YdahKcIplb0D3C28px+AA+DFXENeg+Pwa8ARjvbcezBVEn3WQZrmB3V78d09A
KWA+Vkf3wPE9LwlPJHefIFV85oIHAQHsch4F9qkORvDrTvQmUGYoBqq9PK65EUy637wHASP605JX
GgHU0MGEWvEc2YemCy5aNqSvicELMO6BR3Od732G7xzsWYbMQCq0wzYg1xktdIHuNNRnPeSZwcpn
hZWpi23yHqhkNf1qowph58sm9Cbl5eYC/NMeGdZmDT6A6vMYA+tFMOOnIoWA2bMd4zD+8KO8JpH7
CBqxJgwJhri8Eyg4k+zYbOOfItd62qK+RxGcOyiWgTGO3bUpN4A6/FA4opPkPCOK7jyWsBD2TwMA
13LfUKcw0LpludeR0NXI4LAzyFjA40OyZ3n38dC9yxmmKY+bR2NaKFDEccvOK7t+rsPn7xx4NCGV
7WhkPExylYuJ5OeYkiCB9Pz4zF5BcwVPiciDZRVeo0toaMh4K11mGzIr2oKuB9WSylYuHJCQRUDw
5j9/mEvkA60SEup4ogb6IxiaCiUtcCZ5zFNbGeWGa4fkvt8T8JPz/QvV5onsvzxK98LecuWZ1cCz
FLTaYNELWVOuyuB12/1xAaj5Md0ehnOdcjAVfKFU+Vh/lt8LKXU/0xeqEkEFk2vG2rC2fERO4GFt
FNHNMhqFxhiSdzJuuYCGh2gVf6N4XbL0hAPz4+du5Yynp5tVhoJFic6mczpiIsvhcVuqpri437Ru
fRqD8CvsDeaCRfM45oomhLcR/gWUaFfxUC3WK5tyv+kKSJfW9z4gLaPqK+bivskgrQYOU3Q2QB7u
teKLR8xIJzHAQWXPx0NEUiQR3nYnGzpJy78zfbfATbA5CEHumSxfATHzOuKwdgODajAuNCijga5S
00f83ugQgUic0Bn/u88SCMDGWL14yg9vnSNa9YP7XuVQPzd90X/oUACgHpg7TS9TSpzvXZYcKHWO
RH4kmnFnb9zZjyYpsoIkjzaaSXGbrVb9tpXcQcJGhKI9/ceWjXZeBKP/sOOgaPeR72JnpaZGl815
+cDPCM8/UCoKZQL7DeWBDYOffqX93vVF0Hw6dHJcYppHgDxlbfwHDZIaojz/o/e18eDSjttzbQ9E
i7MeW/oXDrVdYWLQwFsQZ7d32vSWTFnw8CnOmGqNXiZCKb80BWQG4JC9fddj40A1levonubWxjTg
I7rxRNMTbpF+onthH6UkrVwpYjQFl+lLhMK5PpBSXWSdppOWcuDYlMSt6Oyh1kTEyVm6NcA7gGy/
IH/m3fc9cChAkEi3ZZlBGso7rYlWd6i690XWJ3oM0awkktKkRjpjc0Yuf6eZW/5lnXFkKnpr5Iui
lh/pZUUVxNJSSSkyEvfisc+M9AojiWlY4WLO5JwsUaXnRxXWEay8GM1lwuS8bPhjs8h6je9z67p/
JpNSDYzGZy7u+ZJNMTJMFkc7GosIq3Jp5Sp4NZVTwbxQNvu99laTZ+ZBAI7XXxlEM7hXcNpTnfUy
2lLQY96uBvPMtDVXejXiqrbzt2zQABlbblYXzppKVnv+sfVPVME6xPDAXJzy0Rs7QYE9PGymA5n1
ZEgr5pnOWVzwGxNfKYNsUjfr7un7wDOhLAHJOUOyWkQuWVUn8UgDU/I04GIrA8GPggaDYafGo/HP
lksU/MNoXXFRw0AL+us6YxdJlc/S3wh95ePvTzshKRLhoae7RXdC8WKrBw1pNx9YG64eUhDZCMkf
Pc8MIvs3dQurS5AJ1mST22nNgaZRPAYd9aFXOmUVLSO2/knxxLy+Cj4iBtwbl1rxv1Ovn0KqMHo/
Tx3+7nEOGAktGdDBxm/THe4NUgsdsXvZKgkukmbk4QkeWKfAnFdm0xXPAdP6ogWP//uUmk7mP5CO
qUf6rv2/z8ub+6wQzZ0UtJlkL+75NlvGkGYYOi2+54s2ZYsZ1PC6HgVi198Kfif8L4LHJLq15TNk
42Stt0+cKv6DPCBs4BBEHUd4wPt1K6oTr3Ytujiv2NMSVa38DQngpqmxa/UZY2HugQ8GFqVZRN3f
Ql615kXyhc8Nt85hZKwl6lY5fh+w4UyImLNDZqeCT/cGiqhKzxPTaI4nrXFBbgmzu42+hMrZP/9q
pQ6rRhXTalGSKMDQkyYPtr66pUmD6sh7HZ9Rq+8aTJIwfbmCAWUnntibeeRirO/xr5MnyvIMRi4c
g6eHyf3+1gdvt5oelFiXDxpaOt9WCY3TtnkX9gAklQeI/hg0HXAza2l8FZogErtq3KitCzkT79vn
LmV0HDB9B1nb5kpf7NWFCYYopCieSDip6r/Aoa0v9t615fSsIkOtZ4glyfxkD0+msyuAL3o9nija
aBxZTXj5EN/NsOUTe9uMiHjzvhR24JVHIHqnrB2wipsdCLHl8UYZS+x3e71O8VHziQeGdo3u54Er
ZT8c1iShD+WoJ/t5II4yCaqkRnj9jE1seLyCc9cJLofXifiDQGpazYfr+GRUqqY1gVcqbrYaCZN+
9qmJi8pNpGEhbFILrQl95pDfMlyt2TtvF1kudq5Yjg9le1jOLOKJMuQCFgDAGNLsTFAOUi2kbgKz
E2SZyorQUC6CMdGS7RI8KXRQa04DVWtggGInkm3Kre1svq/f6X6TZKf4gYtEUpKzy9eRgGwvU2pI
M1kq/eLaqfOAx8tVZZGA8T93pPJHnv8nYHk420AxBoL6GWdYuHckzyPZM02sot18gwhvnEnKpJNB
wDimH1vjjx7mkctAatJIcn15iAMQS5XjC06ocdSRia2yqc7kP2LUyj3mXINWF4tpa4Cx5s3wdfZC
ryuhmiHNJIKB67NkKuEVuotLCCzNVEuZ1I+ROXScjmiuYMzJ+yqRy6odNXV5I2EHJ83QW18y0/Kr
BoBTXUxuJ6PD2J/LUlqTE3IHE/3Zi0ncmJvD7kDGNrde+4fj/QPPg4PrjkP9Js5p/PtFGWdgPn28
+kgiGEFoG0TxyqjfilGYMitU9He4He/CjsfwcQu2eMTH8799QINhvsYxh3HNTF/LfDRmfZruJ5L4
hpn9x83mgSCrFdYDudEbYa3ZoQQ/scGUX7uDMnSM2lUvDJUPgn7Z7ANzMtLPtYxWwqJ6dO4YMJf4
bUY+QgEpaQqJVaOhdlV+zRRDYRPIzyaioO03HfiPvz5k7bKBm4vCOT5KzAjV+dk9dNnsmO8srVtZ
7FRd5qlicgxE3ggn6WY/2+AW5NRbGYdFT08AbU+v3S7oG5nS2bBECDn98D9430lit0e7ifPO63NZ
Hph+1jehtpNHoAu4hVppRPlKfmpbqvDyZSnteK3HYVogXBOBSxy1jUtIdBhp5kuD50OEBXrWzbyX
gREYl0VeimeVaIhjcwu0OppoL/+Y5I8FszrR/kNHDtHZUR4QqbgjXRSdYt3jVBsdTfQzY8JGW7u6
uTD4z5wFtCcpsD3IJfPS4n3cR72WZXDsjTBcuhpc2xE6040XXGGyEwJNI9Wy9KhENVJp6PbuFH94
8zbGo8MoK6fT6b8HtatcPoaAQzVvFaaGb1BMFA+5/lqpt3IdQoCNY67XBEEY/8BSJFhLraxxrTlY
S0v1xpSG4Bjj53aEH3pjLlVhnKyCfzPWtJYWjqg5ACV5vy+goKJoDMZg2SR8k0JFWRsKXMCI7EjL
SiuFqbAnbkvyZkC3lgw3i66WTROL32BrOB2AFR/mm6Iif/6rDYlwgUChpANmJ3vvAbhzzQtfXVkO
fbVA1mnd29Xn88Q3p6ZqI2ay6FhTRgDFH98t9xf923iKy3TfH9Z5WKbVv0G7Br/Ki1Fjc3K13zUm
54/sqfrVxFuJMNL1DMYDV1e26d0ng2PO0+l7rRgzrRaISBvZPwVldUjEgHd7dfuHEaqSkII2vYhS
wGXsuvaUDTevuNxseKN6clC23lZs/efa408R64vNQMMTBp78u99LLL6iD6mmpORvc6MFDHjg2VJX
jpvHFWirWsL34kP7Qka0W+cvh0MhSJ6RKQMw6Ve8SaVF9aEhuYFp5SMeFUKYp5+g8Db6ovt9xfwF
LT4BxOdjqr/817k3lbOtinhtOSkBrulZD5bbXbMmPwfk0x3l2q0EEURaD0jfIzyB2XQXIDS88tDC
SdGTSr7NFp47hQ+QMwzer4iwSgBrYH/Q4jEoZY5X9vkOM8zwVVXz0CgbLoG9nZt00NNjaBULVjJf
0JURbxwf2PAyrdqCcwLA3amd/etncZYEfKG4jUE4OZEcKGTnCCZX/pK8jsHNkAdfE//cgKGgB4KM
e9mI8ZVfgaxYqvLoM0YaIkV0fWcE3Hh5qYrdA/PRubJl06bB+mUtEfjF4a2p+4RmZ58AXeGmpsnr
O8x1H4buF4VflYeE57cPeNIrUqxchUdQbUUFKrb7yC8+BpQNL74mr56U7j9A0tUHJ0KpuJWeAHRB
7Ujy0F31HdF/DCO6bAk/OzCf8hk7dZrPqdTHHBLP7uL3oDRYyJdDjYmz/bCD0Bi/aj/nhqm0UGqK
rrqZZ9RhfZdyAd1g6mprQFYcWvl8+SM/Zzi2UmtN6XxsDDRh7mzy6NidoYIrlCzjIbfGNLqpf6o+
EZOoiYUvyRs2wQ9aOgF3ETBO6KHcqtjnZ1wBr8jx0y6MoqJ6Vpw93kZIh7c1X3V2m6RPuMqQQbrU
crM124tqlvc5fzr+zXbZQr2gj9UNzsHMIO5GWiSG1szrdWdUWGdbbQaPZ/Kj/428fU0YMvjfz9ob
DJ0pE78fobVur88ylBq1GSBtWVi7wxQLjoYbPQhTDFIZIRjl9nR3okhsPlvVoARWMl3aR1ERm4mk
eYNr+2y9OLejFl53/3GCkYmMvEiKggG2XM0c7tgIJHYHkTRdDrKiePhTr/794F3kt8GFOQHjqcbq
PvHlhe72BTeStlq33Ww0farLt9EQ4DXeO/o3cRcV0NRewH8lbE606ULxvb9FfjTqTI3BzJiK/tNq
stEeMxLRaP7FH3/hU5flZhPtGS/qOmxklqM9db6GaVDfCFRBvZxIZuxbdYC0oc9GxOwWyyts9pGB
G9ZUksMr8BZq6WFxb9a3E6NW8rz7Uu9w69+HI9Ih8QILi9p5oZfhv//VhcPHfx0sONUinxc+Brdj
qX3ykMACozGOjIDyJgs0MBlltPVWXaqT4tba3T9od5xYpge6zYm74HNmrAbFebyxPw55FK7+wugC
xRyX6zcwFxR8gImQYWol/E+pvExzU/n3X2Sj4oINtwAV5KlatOugBaZjzu7RolaLpxfq8MKw1LGi
tJU3zfu3zQacOLtes+CVbjgCfiynagitEddgrl9pSt3TF4tUKTbiFK3RToKLYNwgliU2bu+wSgAZ
Tit9mqVywgR1Z/50uMRHmtOd0kqiVp+9B2X6kr82b2eNMskgsOcw+ocbIn7JftL7LQq76VvdyXSp
FHXEqKQPtlouQ+ReOJYlfI6MYpZ824a+5qsjKqPUCHvwxnQrn5ZqUL8Y+yLZQ2BOI+D8/D/uzVDl
AfmivNU44aldFZWRu3ae+XN0PgFk3uieAA0X3DkYRqIvFTu8kTM+w85SkmX0H9VuMPEDWBS7Z0DB
RrjDVjcY8kM4mkUXOsPXiSXT+bIbsbaeTGQKgyuMQHdBgtAbqjUXJ8FSbddAbzhIMdylhSvlhGLY
0kKKNp98erwxPTKP+cW+wh7/t0kPnmJcZHbY1oSXwA3QlvqB5V1t0GAuGEDN03ebCI/8DAmL98oA
/sLfdnZ7hNcn4Tk/0A8GUoDQXv6wxGIcUyojpRuIr2q/oGpFYpXPEhNNBDNDosy6PR8NoCywsDRK
vxezwYlG6dX/2ehd/aQrfJJzeZWSt/QBtCfHYdZXDDHhCcSu0a6DJ0Mj/Xj1fifeZVbPBFdkubr3
dgruwBckEtnMeYn7hCNKkUg1bbeeDMDTLBMpgBmfV3+Fvl89aHQ/OjS34vjMzJtxgvinqh3fY7p/
WtFdTfOQ8PdxsZ3JhTlm85xe3fqku6E+ggX8fLKxvteaYj20kfd6ZA8nI1CQCuXNzL95Gy2sTEwD
bfVWLCm4NdXBDb/baOcPhZ4+rGBVaGayay2b+ORi+OKckDJnlOJnMdB5TlXHGXG6JP1invlld4oL
yuEuHUD/OJ0VLUZWdVb3YCIxJhM2/YmXqzIS3s/+MxKqtv6p8mxW2m6qLCI9byZAVQYUl6ZwsKE2
aEnwxX1noRHkFWhKHoSPjp6l3QgXC0Uv35fcTbh2LlKbjrGIwwi5CqKrExiU2F6r9rhs42Q7q2v8
U2gutjaweQD3qYG1oFWTPE+21mAxNCqfWGPoIWoJ3hGCw51LBdoOU4wqKGmZF3v2mh8rKiKgYTiG
wxfUYl7AZ496SEwEZNJHQbO7rleGjS+6sDF+qet20mqwqBAbNz7kNwQaWnfYlrE9ovDR+mEf1H/H
tTAQW4lgzCleI/RPo1ZtFckN0Zz2JPEJkRBI6kQh0qxFmdQJreuvSjH9X/+W4oa1CohVZfmq7ieO
nuWDJevprpDWxgwh74un1uEd4lCjPLpQH32DooN9NhrzNSwD5kaaODaXNR71ZlCHKuB2bV1pNkb7
gv6tr2X84krikAm/Z8oOzaAQQpLsRRvLlFU+a5YVraQaESVp/MwDpbYKVuk+Bwv2k0dUcDGUeeaf
ZPprJgNok3dD5FxJrRWA4RCqHgTwB0crlFRzl+mOp3qpOfnu3zdEQ/B6SqZQouD22DfbN2rVebzg
DdaQSo8PkAW60W8kck0GIW4goHvYFOzPjD3x66PT+SUhrNQ/7io69u/q2lkkjzJb1CBzv3J5XuXg
uKY1AhWNM8bK0sTYWd7+DQslyL6bh8ZThbpS0TCeXzYjK4f/ospQAw5siMQ83cTChfNI5I0PwnyB
CYhv34vUhwKSY0dwoW0HX3P0SK4zTDLyTqHMkEHo5CK/RN34RJRIHlcDrN/+Wz4/eZYvngVZepgp
0kRZ4NfgBORaDvDtn/G+FkKaPowGjQEuUcSdh2rcobJBahapg7HQpKS0N6uxQE18mUgb01h8ITQq
DppQzvYf2mjLyGVaOuTc4syttKaILJWPrSVxPKjT62FGYTI6T2waXwpnOrAmSOZYAaupR8py20iA
51K1FUVV4buF3awaWZPk0TZh6dIRN83t37N04qJkiw14UIdiNV4xaclOWgRIKu2ZcYbajSGu1Xf6
pwOxG0PWGy1I1S1sTlX2Hto/C9j4MOPV9HGbLzSMzYKzHHNxziYjFMwmvyVTKWMAa4qWP4ozdHmY
OOVkA5o2gQJwlmmZyT1auY0GZj64kjneAQdp27c5vyNQFpjXNIGhAjR4iPsCvqDCzHcUNSAXzzTD
NFHcA2IfIZ1nc8eiO/2DYTc/VjUP3ACt6OrtO4TseRIKzKTIO8Wr3giOrllLfgZZ/4jIvedQ1kFU
Y5shuM+vFelRJ/45Tv9k3gO16QYtZ95iD5M2qFcdjCxLCLfwiSOo/6cTwxoaumQwsLjCmDZXG51X
LmKFQpOHwnZQAJw5KtKS243j1GoXOtOPpJfdn8uHqyTx8MT1aM3utjTu1tUTAmmwfAB3gE7Vr95g
xp1XxE0mlHJzBHbM5t51r3nsCqPsGQhIcIqIaiXIFT9i4nL+YKNRz3ZlK5SAqkbIssmj5fLh/Pwj
TVySohVGFUtN9mrQMIlCWgmvG4natHAvvR1J8A9RO0EcInSLH09GnePxeXa5kRArLofl1GpnRjQl
4pN1AgUK2Q1LNn4lSDxn2Jezvb0TVprIgDVfEjcmjLu/TXEoVl/2utoK8KBXDX3eWThmnJmZYHTb
l9X2bkFEsWfujoIIvIFL3xv6oaOkS9UjmJusUq4O3GcwEEcKDXXKzo3OYc8KnCp7XIglfgcgm8pX
kIRMrTinuyk5YvFCgiWIlOuOM3HByL3D9MoIJRLTKhA9nciGYGEQKZSd3arHlg2Z9YB+gToCHViC
SNG1wOucb7vQpWESguadPTIc0rF1IehlodZlKELod1XH4zP/k/wSPziIyOTGgrJQqqyld+nU2cJZ
Pn5YKxy80raL5nV/cn5znvSx45lTk9wjyYQCwqVG2hgCx5QhNCJfW+BncMkfkRtSxGu7hNGs5Y/r
dd8EimULkJesM0RVUdINAfhVCp1yVFtbuozz2wy56iePsKmDG4suJTE3GE9YGHr8bxU5fgiaOuwU
vOxAERy3GOJMZNc4LypajQlCW8SpBHUBlGCtSKbZwsT7PUxwaY+EfkAtuN/+qUAhvOVvnTGKNiQ2
mfSUKpSq/RfjevA9vUzCwrqNIIBfN24bCNbNvg4CKCyDXPPzLyyg9Ggmw4y+obrrryAzOq0OxBUi
rku5M+J1ReEOIy78sY3nH3/8Y3hq91occECwXhBPYGTRRLpxOVl0xAUUUQWMKe1AgBktHd50OK3X
QbpPJD3PIvOdUtfWUQPIQFr5Dbn7woH3FfJNCoZuVFe7Z89FNnemU7X0mLYrg+u3TcRt+pDiZFjz
tprH9lxB6G4wxhV4LF1zKqzwd0Wj0YGtTasS/UQ3Yk0EqhIcR6GuLSVVD6PLSQHfVmc3TUsLxLbZ
IoIbCWjG8Tvzdoe9wjrFRGCcv4dQO7etDWSJLmBcSQmx9VljUMcKqJvhCy4VhW+FXe02jwM3nddd
tr0VIjYwZZ3GkbsVg+wZ60kBWqGxfKMmj4AH87nYSvmdYm9xlgzbgqIxYVvdgkZADVQlvByDaai7
E5XGbxFbn73rpiRKZMNucpm1CMR2Qup4tRyuwT7kl2hxZKqb4HoDY89IHPZzhneVaKmx81I3MBLb
wZd3/Rxj/K5EmMeyXe9h+ihv0iS0R4TNOkZAhAknkTUelYdWYU7O4xQyRGfNN0RrlnibRZPUj+Ct
GYbjXdy/dz/WQtyK5SBViXxnI/KDhpG+v9LdL9XKS8loWhmkdXbalNZ1M7EyDUZ02WNCNE3HBy1K
Gi1ALThzHLyA0ZbEGgKALKqhsKHqAzqrZNRx+U6N69xPC+gl3v+p5bMXvf5tR2euoBZmF7RJFnNP
+81BX/pgLxjp/4z2qlf50AhAUyNkDMmt1u+rymFnPlcCCYnG1I+zVM8ZCGGqelkLOwsqVvF+ZFxT
nnhG7B+pd7bSspzO3xYgQ3mRY7k881rXEwvGNPyT6/tr1ZmJN50tPIlsuXBuqNmVUARtkrFgxcwa
3dGvpacblREpQ8XiAiiH/Ja3ETqC45L4F94OPSLVK7/vrL4EeRZxCRe11vk1IyPhHI2AR+hdicv+
yvkN4b/04Y3BzLq3HgNKUfCrBAmmzSCGMqpBtkc/mosbGCEIzVJO1En/sPccSItczxPhY799BUJJ
qejtn/NaW6uiCIJ1Ux9HnwVzxdBlLtjTlKVdW7YGw5fRKvU1U8lJhJL3gVex7wHoryzGVmVC9oLN
uTHsdNXhqJckuDqt8Rmc7BLmQWJuJ51UU0Zv+rd9kBCF2muRjyStNQhnkG9Znu6Lfl/ZCXNA3ogr
y9GKp4lyX+dngkc129VnW6N+3QpsLy3r0dCVSwtI/hDdiTVPBqPfVGcEMwE8PBrWtusnmZLSL490
tcKU/un2cKB5qwRwn9JCLGJ9qbg/V7EG3PTdOVhyYBd8pWO01rsdIVLphs3y/zUSQ3vGl1W9w43V
faP9dLRoq+/owOHeGb01nXOLTNDTvrbzMzoC882dwRutTzFWAUPyU8DKDWM6ELHkROsxCy/BqQx4
LkH/ZoyAqSSZTJlK/veDJH8f03PvFSuXEkb2/rWNGAjIy8bK3Jx/WBXDQ0FgsU+9BqB8o0OtFBB9
ZhPpOgJwaqGsBlfa9K3u0DWvGWRrLHJzWqNHEl8+g2/xoi2WtUXq9jieN7Bx4/6843cjuXUTcwms
5EbH1gS7jDLkj7C81/C9DyEqx7+GrIkQeeXx133pHWdniplb8EtkY76VTYGDwJrcN1RjUF74ENOM
6kPsobXfXtno3m7ReBYHB4JVqNdF0g3e1ynbNQPLEN+5fr3U8Dz95DGodWhrvsiLj0wNqrmj/SvR
R+CVQGoPdsBk26+okxThatEIhjiSOFn6JewTPRC3XDpF9NJEMNvAowpAeCdN+FKzJjvzmHY8KCQS
NZLaO/9IBBK+aiKItySZ4w5bJcgcMNYDNRpGACFvhyDLZJe3OzdLxWPXetfU0fn2LZKbulKLS1u8
P+G8ky2rPQNWsaZ6N/ZtFsMRPCSyujnQsVfzGxnEANETqBnBcnuwrLO/MMPXNBBYDbUMgt1deuxT
/GSDDVWVjUY3qyyKPqIWE5BNJkTFLiSx++Y1Ypm+Lk6S4bjnXLwimzsezgci+9FiD3lYZDDOTU6W
Anjo7P1XtTKQR+wjhSs36eVq9sOiMwdtRXAtHeSKLf10/1pOoAdw8AVo4oCSdchqqP/6guQY82At
nUsITTdV+CkEx3FmplCImbYFdPB7P9u91SbVqWK2g5VcVm449qnfyr0oFdZZg0W168yR36gOw7oQ
S++MimQFKzaC6rySmkxjA1SDW4/rDEZiIeGPZGUmOXp7oA18hZBAUzmqxz656vnWaRqxUh2bkvqz
GVtZLi8Cj9JkrnFXz6/ieRQa5UMGW3PnCUCdQ/yryjWRyZdlJNeE1APmykjHZGGSir21VQqmgeQi
IflbVFeUqS0UJHMm6gCalGThIa51QYhlQHNm1V14oDAd61UdI4f0O2sX8BszbL64qsHnI7Ed1YLi
TEK7Mr9EDkivwI9b+F1mzifcDPxsZY/F/29CgNlyMM3NKbVL0XmSTqp8onsylm3KCxQHt+Qq4VQM
jvcCqp9ecmAGWncJ1OknW4s8VgdAFu8R27Y6knbp+tCdKe8DyJlSoNutNEYVoL1m2N2l7JZYFsKu
r5TKrywn5YSlAiGcnTW4fgXTlfSSRJzG7PJXSvY5WH29RQfVuvuQ/7/vnr0VjQcYZ/FhsB2/Pb7X
ZqW8ZzLdWL1243pkqj0ZetI64xEVFgHF/auBsnMvUFNzPLr6xHDMjsfaMk01zRVUpsFI5QslrNsF
Bf/aYyHH4IAeZ5Q9uC4xpYSRKAp1N5gw9qV6PpgfeTvGNAX4CjCJ2eFg0TZATUkU7Na4iO//c0t9
NVk/WIVWyjQWy2miwlEbKJdDYa2ilK3hD6R9bpEHrBq1WFl1nyaAwwLmYpgeWotSto6il4huhkgq
9Rm/dwOSeIZgFI9bXNED7bXKRwwFTwhKjxlZ56S8aiU9XuYwCUeooP1SJUfqiMwcUhPXW+Yz2++O
qzFGjJMx+2WYKHDuK3aXAVemw7WKX1geRCCJTr0HylZDti6yu133BIqVJJtz0sRmJ0iI2R9XwZky
Iulu6mXdunhKIHHVqkMQaqr0QBlzqHEoEDFuIaTLYY9NK/dryMSlT40zPp005boXNw5etl4QwnLL
5d4PA7m4NOBYlHfLgTaH0ofekaLBwY/NXV42cmhS7nK1bHcEbdfggJ1QM+7YN3F8mX/Vi9VRRnjs
v7ePH0WgFTWcnY3h9dK0nUCl0U1nb3ZI7MHA6pnw7urHttrzYY2OQhDoK36S9vQqOfX8i460oJeW
z3iVURoW/BNhog0aLxsOvS6ExXr2olDDUVPkfLIvu8+uH0RyuonVzxf5VPS/WdJOeeT5DaBZ00dB
9y4BiPWQjB4pahKt+vSDcz6jWBOUY/kXP0hjzB35SDE3UY9+QRE7LmckblKuTcqyl5e1ld5LiUmR
vHpiUmxghN5LCS2OcjwaQSZPE2js2yhHrEUOHYXrrWd5GtIAl2z01sk2zEYm3PcgENoat21o2cNJ
XdhYYT97LYEfM6TEaVdFu2CYaAnDIVni2lR3VMPMwyeF+HxOSwyRd7CZLrkcWeExkWkgJ/FihSJV
4u07g0sclY+ef6k7+ZSIPBfg+jYuZPMM0iuH61B93jeNcg8O1IVvP7IrBj5buW8UXcJ71B1xB1oC
/v1EIJYPXSrKaUn5veAgPygvWSvsNZnO5qzQ8Jc4J7F3oeZQQMQJbAHzOpjreiTVJ9ZXCBkXrhGi
8kpZJS5//ZW5wHvGX8wrjExUFvwvNiTDc1wsWJUZCxooBC7amb7hSI3LZh0N+OK8P9Xjebu4/Gbh
zeUx8aoPeSFY0s2eUb1uVxQCAiTXuSNoJ9lvx1Tst22tqO4y9Lu7L3IyoLKhErQRFRE8+2BxPt1R
P55IqxZdVNV/nBz3Ji3fl8DLV9k6N3aQkTpsBBy27IRIC9U1D6htgE623JsC1K15JxX3C1sAG6mG
ATvoyhyS85GC74eKcE0X22WGyVLootGN8nlHuaifKWcR6DaIMejwpRklhPjrKKY6K6AQns2bEVKS
WTSmxeCy5/XEMTLXygW7vSG2wnVAdgfpDTqJsUgB0fV2uOFiE3qeDffc9hiJ3lIiGt/D4DcHz57+
zDoDJMpZ8y+w2/RPGDBsZ2kdw09R5cTBGjNeTLKrma59FwvE2Kn9K1h+3X/CKXhAMRAsZYU9qajJ
deBnDgAHySGpkzKLrmt6x/pg3dtgPQlpxAskDeKmCpyd+jj5cZ6mnqeqGH5pmcA6q/G4fRa34EbP
pSd47sQjHECESeO1/uhjAAbKZKXHnTJzSD+Fr96nmLzvLrVRkJ52PG7TenVcJn4hIKgrVg3v4K/U
0sBQOnBo14K/x6S1NbtgyaMyDtvZhzjEMuxsxcRlY2otq4KUg3tMjmwMsLjbTi3JtAOViEpnDAmI
kHMV/P161aK3pqxjC7UhWJ4sO5zyPMjPe1k3Za1QDUyfQDoSayyhOe2haGvSOjskQgfwe5tldx3Y
WMZVf+XTXyi/KPuwf5Qw9O5V4UpMbnfit9CBqv/CvVxc+1FiW8BPo0aQhVM9Eb36ZzBAYhGKrOrR
hVo096+i9tska0sWbDU0koEVkk90X+KzEFBtu6+a2wmthuYgwvsz6k0rQvue2VdoJpi/aWsabYgs
MFeAC+7fNQk64m9LMPHl06Wrwkha6Y2Zbkf1WBwP/XhwGEumgEyrvB2ywA+rPgJez9RhVy5gJZMq
PwcCpoaMlgzDS5YWkJtIkiDxJQaTUICHe2mQlnipFYUl/wreOEuzqlWOHxIbyxQbx5PN5r8p9Ynw
r5YRpqq191k1cWh0TitLOqNUDlbP+Yuah6H/ewkYaXfZut2rkVp5dPShFTXHcjfPgQSTqH/FqpBJ
XVyEON91P7vobIkQEAjFas3zmEv4D0iDHCiz7EH2biF2OWPXvqz6X8kKqyHikMiUkNRzfWqTdnkS
eSAClyHe1er/+nlT6V6i9rA8vPzIYZY9HsqRDc2rEmxzpbYhr0wBAu1yjvm4ygdRv/M9DfN1hc6g
CcrQPLBgyXVJl2OLgD6hPuQF3PqMbYycCzhUWQ4ZG9rvZW/UVIHUSxRshjhExYr7IdlY3E3sTkKD
5hVw2HvUVi9EEtJx+r5dVJMRwB+AiCnryyQgbGSXVPmXeEjNDhcr95EAMp6iyvHJywkRu41p5k7A
6cdB3FTd6/Xp2kPmnaG6Gvk1fqPc+mPYw8hAOfMAbYDA9GWS3et1UzgopAEwwORBr59V2QLUzT63
Sbgj4F26Cfa47dSljdMDrQkNbutRRY7GyfIYEOddWfMDqUjLTntkH7oGD7cziU3qUzBKrsztRX5F
ZedWZ9uY0s/mKrCiBEKGIJDy6So8IONB9gTpLKK7hV9J6xxNtm/Eab2N04NJnUgvg85GcWclbwhw
xkYoN9VLDYY5cIJU/76MG/ytwG2RjTmXKgwFQZ66w+s3jICVChDUypUW4AJxzOSLMvEULWGWUyuZ
UcgNh9+7hG7V4A0wWQYKZtuxCLEdk/SpJvn75P5mo3Z+4H1sJcWXxH0d3XOP84eD3dho3olFIPkd
99auPUris2aMPYwhHT6YdZcH0x1/D9f0IWlAyeQKz6IZajspvMq86OZVjAkg/4paHhnNO2zoIbqM
ut6DL5i9NwOWy58Um8feutRvCjsOxtNRrNLTvH0hosZS/K2+fC7ccLjLz/mtZNuiIl8HiFm8Smiv
QCfrxk8QfbJl/KXOJj+yhHu4O6Fu1YfZ3+qDByraHobNEGe8fdm8qHRejIDUp7fY9di35TAq5qxm
Bsg4DUrhapPPWKO39wsFhaIW6TRqwcGWyVe4g4uGOABE45uGanLb0cwNPmLxS+iSW/UjJEwiDJLU
h0qhHh11xJUMHrVlfN78S7F1lH2ZZh+Va1vP9aGz9ZOvI0TC+nvtfyv7EZWm0mvn5xodf6KZzJrB
VqfF49htB1i/sDSNgABzMjpPnC4JOZnlI50PnfWKz+nF1j1d+VggxOQ0lHo9JI80jYLZLgo5tC2g
nvMSv2vA5GR5y+UG8+uEF0Fad5Xr8dNrV/Cdz3uHQIFUySKqt6tOMpzx/7R6pQg4j2VpLTyGQcQH
BNhxXrH2Ay3sEYgMS5Y0MAHU9AzhUNY3pJ+f1otmGjg1fyBamljeTRkzSFSGnNalDGHYkEEVVCFy
OFbjAD5QK/WzkAl6nk8RLQ23z8KMwiw//GSKn/DK8WcTYYRZb753MD1Ccn1QGNByeYyO0RA4nMYh
qlQHPHH5EeWJDfGPCgyt1u7pKGBiHZ/W3QiSWPpeIYRsCFAk5iW+5Wnti6zCZ3LICaUjd0bzI+H2
T/pBXDksCXiuRits8W79Qe0O8nXcRHOtixoDIc2jcpJLlDklGri4HMHhb64o47dHzQHhjmYwYU/K
9FxmCNJd+2Dz61XZKbDShi3x9fYOElHpxItZtS1bbfONYa/n7RYKrj6K0W7EBEquTxPTIcZxauN2
1FmbkK3YdiiVeGAdDTd7k2HEdVSEGZZr3OP5jQud0BSz4x3gfnBovANk8UrZ+9lbuDsZF7SERK0M
uflNu7DwtQKOxauelMHwNVrQzdJFEwJ1yJYd6innZ2qPNBP6lPKx/uKIY5g78mntMMNy4muWnSia
/b83Gamql9s8GHFZQ4H97sw7txEvSdRhHwSS8yJbjEeVMtopdcj2jQJernNsdYHDIzu6r4SdvnLd
MGbg5F6rB0jXuol1M5bnzBu26XeIqBjyj7iwCangf/vBf3XuUmj3A9m7fa9tMNQ0cARVQy7fwtVc
kxB3CwTj8CM+DcbjX8fiLVnjJk4lo2ZThjI15bIwxDjZhd8euGwchlOULMlqSrsH9wBmxEt0HIKC
pLOJ+ERRhXhWlw7yGHd5acItsINqHxmQHlPFjRbMp24uBJ7lHuRfIRZHxcHqveRtRqctC4NQvdm+
bLtH4Xhqq6FNcyToF4ZPGBiL+lUqjJ2YBunXMaJi5MZ8u5rerLZAI9oIySbV/EIkHyxXBns/+gvF
6PiLcP/SdonD5WJpKjzahbGbsZcoBPEDrutKctv/8wrjvDcgLZ6WEx3ZRr7Ey0RzvgFZZBykIQk+
uQghBfbK6nQqn9/ePmReCmwjBFr0WlSoLEtwsBsKxvjqFZsC+jM/SsPnA592WYiaMWOm5g+8/IxQ
XFm2Sm6sIVNcy7Iqn/tFRAvindkj+1dtfg21WLcBGDXi9OKlzekgBiE11xd2MGczNivFV7TWfA5B
VV2fwlH5q5j88d7Bx/Tq8ORnTmPoA5jzXoHr0nQ1F2nqqX/1TOkJ+4ua/SGVmKzqcx5Ow+1kVC60
GrKq2hRIrDs6ETwAXj5sGes4c6wcWK9PritkviNmCBlupJUdtbYxHsu8+6fBqvYWNDFStB2m3EhB
3ZBsOsBVGo3hFtgKKDF6PPzvfjpDyv9BA3GRfaTbfTD4jh6fODL1SLdIiX/bpHZ+P+epTGpo+Kos
8PKxUH6H97yP6wMcUHYX008mWwL9Q6QwBIYBEJboaP9fNTJBxLMAOFn2l/ETJH9OgQfESYKvPy4s
Y6x1tRVGVKk7I9SwmNLMMyWUOBB3zr/ERrAs85G2EbWEl0V3tsOpu/G9WaMmD6b0obkU+skVNSHw
iM3r6ZNSaqaKQByFOSIqOQ74seDZTeeUnlrW9o5MBF+mWOfXiW9rmaoG0Ydl+IKPWesTDU1sNbaN
fu1tFvLgcBUD3kGmi6W5AMJoyNKdjtCEju8GHofsn2fQL6JLY7+9n0bhvc/QhECdpCKjlnoDGBX1
YaSPEHcgRpPreZzJq0LhwMTQm3VRJ06nyGzw4cLBFUGIChCgvyQy4nAl+JgDxeX1AWVMCbnv9Mtu
reAhC4Aa143t2XX5uxt6IKjs+ylF/VsLQIcUs/bkAmfdaSrBNCiWY/R9TxzyW42f0cHLyVD3EWte
OaZseAHxRed0cpT6x7ZcgK7ynkIfmsBG1RFcPxegSaxOG6ER8Q39FPVUSHuO6YM65DTLhsE5goab
OFw+6KN7K7WoSc4AoS/TLHrNd06sbHbCqj6D+yocaMnmKT4OkLkjhN2kb85kQVxWN3/E4kyPcIgr
0xm1aJlNetyZsVhqSbn3q5iD1vMKfUh341ijfbgGYhv8x/VyXPGtzErDCqbjt2M00s4CKsrPjGse
LRcihRFTOULHvNJnGeIhFa1xdVc9y7FN33oi86fdxElo/RJrSpKiQz3d9X6rfSnC56MzTPWj4s99
K3iwuR5hAfiB0y+dFWfBVtKOZBKTobmWwhY3iC4NoNrmS1uILZSkwZcXopb3IUSvx7YIyRvIrTMo
cRqxlF1U0JsWAROB9X3+pOaysQTq8ugihvD9ITV6tPMS8SVTsrZ/fPWg71TLcA3NoxXUUQ3l1Ibt
s53K2J2DIT53yQSTUIcnjUFMWfVJ2zPzaWzIDpCMQrBNL51qL9MvI6olDJC1MWMZ82/ea2FxBHEE
eNe/xsXIzwbun4r049VZt9DpD8oZRIyNNmpsRsYTQE9DNqwsNj6lpnKSfUoNkdf8BS8xQX73dsat
LFUH1ZPPheefc7jdTX3pg9R00xcgEUCTTNafCJlCRusPty0Y7akxc0MZDfUBFLsu9wXOUZSg0mqy
uy2zZO5INMcyaR8pymrKZxiiTxVLvSiwspR8QX7+qaOUuRkc7JsGYriYBQdTDKP0/fnejEcw7Uw+
uCgYJvuBf15Vh91B8zwdpr76ehQ+6MgZAjVHS4iYz9ORXyfF+eh3EpNn18m51+1lGLC6OcW45YVT
hKxgbvVJMk5cCZP029b10v9mbDbIbMFkUNojbl09QQZ/iNAEuPltalGz/KjCt2yuOYFUycgS8MzL
4zVJsgQbm9FCpcW4dATEMl+xHPqLUFnJhOPMWNePyQiIMeq1A419yHKVCa2yIdowjz8Uy5yyWMSZ
411ZNGo4KXJnYppGWgPLMa2u89RojKJQg5NBs+JccyaVlnV1X5HuD7bINb0KjQq/NEIwza9OlDI7
l/7donpmqN7Fm/k4RIIcL4muF/bEHWHzjfEPQ7NRqE9Evn/rADhaiP5x3ySezP1nmziDkxMznXxf
Typ49m+ZtptTKfXRK+Uf3n+GmJ5L6xhzOeUbW4Q9C3Ww6+ykwf4Igtx1/JJm23y5c1zvpVKUFQ6q
1oH5YkB7xznLbm8f9ftM71tlWEukAfOtlQj8XqMMUn1N5l7+tp0wC0YHn/lYOQDTKkLWrLThM9Kn
cp4F2+3Vi0C5UTTD0edMcxIDXOAyaWOKPgVvHfqGNpINRTW3mMbYxPA0Jp2sDoOpq5FwJDELFgoD
/SHzfeS54VhEj4yHfx9H20yPel56h9FZaqi3dg6g65PZ48zIHb0grUdM20lg0TuKuhkWqfArN06G
Yaj3F9ZUQa0LvO8+brJVTZFpMEYWhV2dys+oeY9qUhxs/TWFeGUoENBN7meAwu1GVar9HqcWOY4s
Kznb0+m99ywCLrbKqOJMEL6N2p7A11Ke91ZGHXNyq/39/WwP5RfSWVZbL79qfaxcKtdJ/KorGnRA
Zt01V/Xk0cXx+hRFCRJ0lqEACtK1ZbqBr70hEkYNQIgKSkN8QeDxBA63nusCir3iVo8ybyiP17vg
TBNBrYoJAJVwICOv2Z2Kk7aSiNKr9rurrTgTJr+jLuKxrLWGwhDDNnGKYdWvi+y9tyexqrrieJ7l
+eMAcj5Q1nBrP2gAfE0U2w+l86wK9XBI0I5R+kIe2DZMMuAksGDYxHB+y8Bo5pZXsARcsw4+r2+6
lJqBL0QNroOGIfRrX7tPKqdR02THq+GgrEjFEN80wC+KDQPsapL6CMoZrqapFZVyzvvOk9Oy+1bt
VwFQg6mNeGnrpS6k/teE+6bLuxrSH4OXupA0gw+AG6aNJ9aKUTMMzhpwmfdsBmwSpLbwwZb6bm5J
o77rEfXwLUEjmyaSmC3WzGBR01pilGDaoQLXwhKtEUvj1GInzT25IgIj/9Wal9zEWUIcO+QTAQ6r
qvdFU4DkbusZ/8rfZbkOEvgq1n8oeu+m8e/A0dD4cjRBSe5MMxrw+ZsRgsQnzeUYqdmKIQiYGX0t
en43M+gMM8GyBJKkhJ8Wc4jU/Q8/VZLq12eL0PiLvNrHLXnKT7EkYUNFWM3lcG3ryzDLyo+BArR6
WU9d2D+Z6DxjxV9tVnmc/PS1HiWFQb+0Nsqa7TmkvLNZBqGRNbx30ASF5kIAPz8dSu6XQmwl0bhc
zdbSqFOQXtHfTjkxtxa193dsM5cyGMf4AERzxagGN3rBRn7KfAWsn4kBF6+XMg28AL86zMn+aUuS
ieL/XLwWazY2Wxy0pmaAn/Ew4jqoNn8zPD3ERS2yizvF1vW5f5F6OFJ0I4/Bqb12xzvZvtjTlcPG
ytQpV1+Ys0Z1i5ugGaK9NAQys17qLkx/5Ap3hz8xYswYBk3khs4rlzhRrbG97AQLb71RalIgFSU0
Zo6l/42kXyhhIWQEBwTVjtyQghXTRXlBOgC6X/tLpgcD/MRTOiWj+3G1xiedEEbxjMjO19MXsluk
Cgw7n40KiA9B89CZ6PEoj5U9wiFaZC5Kf5j0IyQ8kif0LtXyU0kEAWr1vsxTJQ8G6eE43SPwLUM3
C57QcnF5mjIQ8lVDBrKMPceQGuMTj+ZjshOjdyVDxpnOpVQArrFCRaQcgbzIzP+LwugK9qOUKcPl
V+q9UF9QOU+vQ6waUWSNAjdbc0C4sien1ZnSs9nKR/UdAJaqlRsVgabTcDzK+GYUtG3CKXe3S3f+
TSJot+2SuMSUafAkjgiFSi4xJWgfaFAnwXDAp9kYyNQSx9bNHcM6aa6Hct36/F404uxVeSDQ8tkg
gKRxSqss5Dmf0eP00WQWaORH+x/c0TW+7M6nHMZfMYQKqxxhYW+C1quUFEFVJmgke5wX6tD9fhXU
ijcL0oYW+z6uOh80VMDyxAMsiinuPcbguHWb4leD2Kr0+R4C5rCaUS3OviPVdVx5fK88MtvvZx1G
cfzxqUtKoOv9bZcMuuCqdCbttoEQnDs0DM/jJIcfgI79p6FMdIa92Am68ThjH20EDHZ2jClJND8r
Tt5VeZTXJmdcQkB+vqa2gI3mXPZKdsQFNnSZBXyeQyCzhE6zYAqD7ThlP0tYW7ruHnKQ7SbltbpF
WZ4mPiSaQcw1fEDk3h0c4Ozt2xzbNTcfgb2FEILa7I3yXiPeYEMjlWJBoGKlThZL9P4DXSkO10kn
qF7dtyKtXdMCXnBin021oWULp5DGyunr34nabOEv81UIZCEhEiXCQ5wLPw6cGBm8D90rKtEbHVNK
sqKVN6eIm47U7T5KXE6Shj5gqaSfbDKePF7k9Z/iTXs6KrTzcjvEEWwRsO/31WLq+uUsR9BOULID
pgfQgzhhcnVxxnyVj9tWwXJynYF2js9HpBVy2RcrsER8limPiRWj0F6ZQXAnY5yL7/2qKn+qqnsQ
eAX7DJbZQC2TRl6B1aYMeep5Z/1bXNHfwy85ICIYRJBUAjPmyag7H7L+M50d9vHZSenCthhCmxW+
XVERut9Nmd6iiNz/mY3WpebdhYCB6q81XGwbxptolOkwCC1QFexfQ5YfjliHW3Hzi7kylA5R9CCr
wiDQWGYmODrkU1jT/2alDiPUUIHg9C7ZVr9+SMeefIloH5GydnzkMGIgPdZFXWDTwxjJdEQ1xLIZ
srEP9NvcArt20nb6dcjZlifBNKk=
`pragma protect end_protected
