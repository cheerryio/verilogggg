`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 160960)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpIRtixhceot/hCKjnR0s499PVPxdmsqzJhYfJLqyo8Ol5N0Om6X6qC5pN
9Z1hTYlwGqc91BZgdeEaY9XIVYs8D4uKMaSW6mJwzZFg8jJwEhq92Jn7AwQLF8RTqssYwRvpwuGR
0/3llJBbg0lT/SGvxa6yNMu+14oh4j8NAluLue8cOgDkVC2X+vg8aGpx/XqBX9yYQp22Q4P3vTjm
Cwn8s1f1/IPn4Z8iiPjhOVdIS0I1B0mnd7C984jilGiskQONL3nnTk+TQCi8UJzeIN6yulA8qBRR
iOwiQxe6p3tnnkea5x7/ghCNuoM+7DS8sOTfO7TZUVvbS9R3XbkFmw/pc8wFuki5s+foUBMlE29C
6V4/7pUt/lRlNvwOPpXc6mn/+Qb2obh7Jc0kY8KL9z2iizaeiGz0Ijro5Pf1cVE77/wwWw+50e2X
2AwQ9l+W34yTjQ+IMWGUn2uXFwKw5/uVies3fY6cPv82lm7RGMsf4gosgapsFvrDuJBt+07mpcLb
h2OUkwjX6BMqT9NFtj506FEuav2V2e9oVyO7zWmkEMnfDpAv/OfSR5jCjSrd8HopGKXQnAZzFlHK
9wHJowXhoj63qdknsm6NwOaVNpqLm+PoXTib1WMIYiXbGtvnhR1nNT12/OAkt3OVm971h7bS1XTv
PAL1wpx6+/b8SP4q46b1yqSfc3qARmGxGK28ef6mXDCIkiO7i1SNcQVJTHraa6IxlER6s/Ekekvj
fHyepgU5NBuZIf81SupRQz3fVk4ixs5m6g5zKa4W8g9T42ARQQVd3O2OtXg5LJ3RdFVE4ME1OwtL
CD8rHG6vz3X2Z8ZySlUFeatSUJzpN8MHH9j5JjDCU4/rlFSIbpnZaWPkC6zmqQWPwFpcWxdNLfn3
wVCwOcKQX4MfXPiD1G7j1RviXFewcW3EAYsLqri3z2tiAoE3u3ab6Cchs57USFt2tsX7QPmTR/Nq
j4bRk4GvfIMVPw2I1eMoEmbtkUoqk9dWF9bUpDwfzQ2o2cWEK+r1FBZ71qAneJjmxc4kSRVx2YFX
8lnVVKWI6NH46z3GZ5Aa/beznl2kTo+6t6EUTLi6ibaKyQUZ4gKvgKcQf26xFkOK6O+YujyInmVu
l7eHuXfgdGmRw1qjygHhyqqVBGDsvnOVriAotxNR6kwGpT6tBhGq8o4mXsIWvOPtdq5S+Bj6MM2B
DCzCoU2JSGrulm7ePThgzyUwZWuCEXA4nr2wyTea19k69G5HP4WdmmQJHWV9SJ8fOs9Gwm3bAlGU
tsQ557l2Uj4T+R6b+hhaOA1C/4CNlAGkopr4jzB6yiZZ6ph7MiTsBF5lQZ2q+90t6w3gCuWhSygQ
ZRhj4VLDZ4nmXA4w7fe/rU0VFym7joVnAF9scwPPuHkf/LxQ0dkbWZRH1B1S9MVPeI+fLfTbrix8
AT2AgcoW07QXHB5jffCVm4e+Hj/qxnuNT206e4eeT5jYWVWtj6xJT8olhvr60xHjQoohiiKEPLOl
NKmN9dTxvOdum2n1WHiDwXX7Ln0RjsspYO5SdDP/P/P9JRoICkDs6bVv2esQmSp1i5lS3KusfqkK
81Zc8nfGteQeTs5JZYxhigBhE0zgw7LC8dYPxA9tcPHAOtbP2fzSJrdE0PfVUQ3RI/UkLo/GegNN
3zfrzOqh5Hc2TzfgpFM4sDBM1n2TYp0MsUv36wzbUx3NHhxDs11c0KOHUMkY5r2rqlecjDQST3qE
3C1aDEEb2xDa4tss4fYwJu+/BYMKLUL6NlOa4MHoqd6pHjZwKsInOT+ddeEc9tbQNfzWnyvl7fuW
A8PT6fQBVf2IbE3YjEMPyxwIFP5ureGU13BKzX8scb3O7pDfr0j8G7sYsUybFFbiPS7Z7jlaXwmL
lXuqDrLxANMxDG37NOHOydOKfj0dy/mIXwG/ETfWHB+PbojwGK4MwyEaD3RweBdzkzYhXN0oTt60
Ums35SMtFyg6879OloYXxLwOkpF5irlqOlIQKvXSBm9tfk2X4LnjHVo5TPfVn4o01tolQLB0Uh7i
ssw611XBaeMn4gkpPNqDYz2nGwt7hd/36E+quFfYKhLOh8LNZz0TOLnRvp39zcUS6HJeeTl80cqc
6sKoMcTMIodqJq0Cwz3r0CH2EdQTB2XgABbk9hGtusz5+RmPe8+scHeKFrXC0ycW5IRRcjPjw4rL
JODg+lnUGbrheQ4PHBkclYmK23npOGIkAPh/DzYyCdKH2TQjbvI2GJWiBByDUA1HTdrH37RjmJrv
t8/1enGLXi6D7TcwDNoMXVFsh254uqs0jXZ8acGElKeaDXmnkY17ERl0yfHYU/Jo6pquhBUuHf2j
mAnM/MLiiCM1VjEhkDXVbfI2wLmzZtoKoVFFTt3uLdoYyNU2D9mYif42JbvGTWoHO7awGVkYn9ln
FuaAyHeoNTL5Ug+zMKAdOikye/auPT6WNv0l2TFCCQ6tmkh3lrMTx3Xj4escMR8wdghiVszfgjtW
CmbE7hJuhH9te0qgGwdT5f1g5hKfVNjcwB2vcTgRdtLWk9eQnD41WxOLqwj4RgYUk3mUWPOQX2Lh
jOa27caFbjhsDMVu8xj5EL4mDR36jY001za0pYT8OEkqMRt8143QSQnER9t2Xl20HsDJQQ9/0pFM
gtACxCm3bXfEDsEdF1VFdhbWJUedMBhxXOkuwrfydYq4QY+eI66xaiKuOJDQHaAHIkwPfwH/bzjf
j6NAtvpZ7pAYlr5+MNbpRSyXxHSLYCXeR1eCCQaYJtbOo2LxJAMRgrkXpZf0sWZc9R63+P0qmG8x
DgieY9OZMC2+pZgMZKBRKOZyaSzKW3PactZxxk1Am9rG2l5Op2CFqnBybo8IZScPClgPlAXUMWWO
mJx6SJaxpNlMfP2QYb1/pURtDf0xSH8dTqtpCd9gXbLxc2yo0K4uHeVS1GG5vnO+yLJxRlBTSO7M
wL3vlTkG+Lhf/AeWa6pxafqVfzj9zmWANVUgiXcv9SMZk7b71Cr+j6japXAmOsDTmwGGtrKexE6o
KpZPd5vgprDvxem8PWII0LO8GdLXtI0SEyVwDSxsU6o0PBRm06HTRu23dc8V++UdvpfERu73fJWI
CBUKQ8A3SCHZOI/G3Xu7OT0o+02iFRTw+B4PLRt99v/obtTQgi6VgX4dt61k1fH3jwTprF1g50nA
7LjWOfEt0wUg2eMUq4PjA/k1JT1MwhRJRsmCgpwVrFjoUvZFKG6RNQE6B7xjS2YzwvUaN0ECxp4v
RzEGeEOggIP0aE5rDXRJiuetzfpac1TOM1FE0uonjgoOM2NBYNeB9PbvjvElFTqjANahUhuS9W1L
UJH7XmR6CxrmmEZtZR0l6D5+1jBrkdbvBcEdLBuk2yX5N5ltsxiSS15mRP2qHNIjvbbYlaqaDLdj
wreEGVVVZa975cpZSvhxwupjNOdg3je6FcnyYH1GBw+fE4xKLrz5GEOgn2X/mGkyJGnnQuP60Ud5
HPejP4KjOVY1KuuUgylhuG25CDX0yCAZ1r0uRtS+EaeHINMqGMpAG2bkitGLLfk8izM9iUhYZ4T0
jq37IwFfBMosucqvcWDPKA9XFcaA+lbAx/RJrV7T41ZUOshhyFow6UbBrQ5Z99KF+pDpvtUysAwB
m4jmqdtZQ4kKADgY8LRn4yq63LsgfcK8ZgqsUI6I4ussieqkovAUf/UsaUCgrzwQxa3Ah+jULBH5
wDjJqLxhndUpeXKdeW+gykkwhWjAjpcIUvl0uzj8bw5GGQvxM2cHfC8ecqhJ0Mis6wbSWzTCemYA
B0BNHXm4qgAXKThiTTi1Ppaj184rq0O06kQtBtWx3ntYfIVh+wgxkeztuPd60hdJAtrUkvWHDCwb
cMw5EHW/VvcnG9O2mqzroC+lyik3xB/bH3bc5PyY7wfuLrgjdOnTgrQelCNtdBMPFi3KqCbPULC4
oQgK5xJnBErIF5tr8OupiM78DPo9SrJj31woL95q6CKIWCbCkiyxYomrtHiQhPmGhZ0YAWTwnTUg
Lo48lmJc9yqErjPc6n3M1Th64XxThKWLWa7JxNX5TWYua294dA3deHmdcJms/v9d6F3zhD7WpeWb
cDZG3SXA/EGP98oDEewLQsY+10K6EkrJ445I2Q6IYUgvw51iM+fXRDJhwiIm5SgwUtJw7Eb3PFka
xBod1u/F0C4KUhcQLgKVr5R5Yyxr8Y+Ek8qpmCGQR8Av/tSjYetr6OxGabibyOIa+CR2qzBLwNQB
IpgcmIV6qr10hfA6rVhHtNhV7M1HKCIFhxjHS0jF5plgyTVn2hIfjaWaOqrrhuB5erB+uK9h573i
6NEvG0QPdvC5MQFROkakHU+vettky/ILdQQvXO1BdDURSAjsrWVxyOcqspUGvVb33JiS8suX1924
lQiBdYwsiEg5cu16tXeMv2O7Jyq3bQFc06doNn6Eu/NbErhND0mUY+1B/XxYrs+Twbr+3S+HV7eX
7B9YdyrVXIUqSwr3REOm31zH8pQSA2Fcw8dR6Y3Z1Zs5FHsaCKBVbR8MVw8PseN2Ab6TMDMS0hjm
UvfH7l2VRsMBLqDL2U3WNj3mRG7kLSpyCYq0C69+j9qcQgA4ajjsfdZw9ker5s5gcdj+EskRQlyh
m1jTG2xsJZPToveQbmEhThWevb+T7u/Qu27c2gRf5tJIcuSj83xYHD1Iu7CCbNYLdVESyi1c5RLK
g87CVVFR7vo6xqcqdhgbp8wOXsLsem6VTySVcPucTeM3IlNboHDhT4qqbtt1A/4Hg2xUjvYQAc8C
Mr2tKy3wQN/dq50q4YdufzY0rP++Uz4nX541OMQPHiCY1hZryWnIbdTX7UHj2nbZ9xYzmqYCyHIh
uJ4vc+tkakNTGdRusp7AgnwBLfmpUpk6Y1ttnpYce7mCoUFpC442ANZWjFTu42TbCuoAJ4UJYWNd
/pa/3e06X45qohAY9wCCTDtkDlsbRlEFjWENHhxw/tHYB69BcWsRYeBhRINCvpd3gS3IY8q4ikdF
Ih04i6uA8gd+QmW8wCwfkbqreaJzORrLM+Omd2xpwFtGoBxcodwPfmqjwvpEMIQKkJYsnQJ38UF6
3Tx1RnSRsg9sR13wR03CPf9VZlX55JILfDT+8OxLBYDAPz3X03mRXmqbjglhwLSNZIY6D0i1gUqq
609oK4sDgrlrbRQBoy1MELeJmeUWpAv1Nd2myVUlui4XvjIGyE9qMexy30/+XrgXYmeWxZ51jgTa
S+T9qF9NHJApR1lsEVCPmuCM/g0/aEyD369H3to8P4KtHTd0NOGfsqDssqxJZQAU04e2ETZWkOXN
sW2nVPV3iiijOs2p0UNBtl3ZuKnh/2ozKhtkfdQSmZSaA2tc4+PpcIEhTQrKB0UwnvFkxBogSf21
MojvPSdltOdG966jR1ZWv7WJpCHKMKdRiQllpkA1ZQHvkcPTwA0w3ElKszOa4IZr9+Pb8ugBoFCR
V1VNalrlwr/UdlVC6ZNf1dqrNaKOrNgW8xL/vPsmJn6Tv+i2k8N8yqFXl0pqtf6iDwDOwtjrLZFF
VTKICwJ4QdFhPgM5iN4YlE0xZ5hNEgh2OQa6HYz3DXzAKmda7GAvVqERL/4P6FgZc2gViGgKowXK
GLCjwk4U7EoPA8P+55mOxv/ryiRSUr1adosjc4//ccNBNJXilDC91cg4b1Jg6sfaik+hB64/Co1e
yHxr7MUfic68hFvzYmtU56mSZFYS2WJhxcwaH1UmNkQDyRwuzjhbvhz/VWH3WT59eBWEZOUzGQL6
DheLhOvLg6YZcSZooQZNSeqLXTtW1uuGNqOLjtoMkZkL319tvCcnnjdBitg81fh5bwJHfb7vEOYb
TFVafIR2ESg7Kmxyk+fbqZnv9qNfqhdeYF7FxnH+HvwbIVRX6wBULnYV3maMMyhZWTPDppjXSSdz
ounx9Lyd3qFeE5CyzxFLJG51ueyok+MpUoQXFfYxYjVO0cva8td0HDDpuUPRES4sAE4CVeh0chkI
RivsFtNZknHm/zxOaHUmv0OLwJLBhMCjXqDBaqVkndFlqqy0+AJCULWO8y/W2eXHXO0ycP9wAK66
Epw7OXc22XX762S6GOXML+Eo26PNl5TzTGabTz+1VZ8rbfrzfPr89kh+A3XhVqLrA2s5ikx2l4gw
SM1CsrI0SXJa5tFz6aLypvn2Zkp9SXmMjrsns47cSllaassJ6E2sF0x6CBg7yCS/xCg/nbjJyzyz
MBNwvXj6uTLuhIqqagw/tb1OyueXV3SUYyabTgV8Rqhmj59VwjZ5RNPCsFl1P80+4r4/9lX3huDs
1XE1W7Oau6UrYJ/vYpUZCXe+sGDEoR+FLULmjqkwLqutKddnp3vylb/g4PLb9BxbVC6FhO3XpHQo
ozPg0+EV6v9Q5Vks5j1iZsQg7OgzVYWb13aDZY2ML+EeL8bG3TEaCQGhp5jmmRW0h+fm4pt1BK5y
OPH3IqPW1KzqL7XvN284qB+ofFf7vVEoU+3NScOtnUmvOCbr7UKt7BWE/wxHzK5xZF+m2xqdTtQl
M0z4vPlVHvozTlkukS1BVOKukD/rWIXeAKSTSQ94b4yuhL/JmbpHadgEHf8WQznA6lyW1FdY0Git
luIpALQxky14crEoXVcuFTeCvBvDnu3P9W13am5149AKp7ix5ow80Jfb7j7CxqpMY8rj638ZOeNh
I1rPg/FBzHkzpJdnZNA1eiUU9VBb2RUmAmskmZ6q7fuFW/Ir4m9kIfzOEG6hxcpb2Z0luUXr1SiP
WDNt4mn8DN8d008EuLQXC8vfPM7yUHIkm0UOdexPTvE3P6tPT5LDj2RrEfCH90oaqBS65P5A77/2
JiXGLeHLuT5QrxlomC9cK6+gDRJ90xNkV+1REVtGv+5YBWHne+SjBok6WVXnRbl9VqOk+1OLMPH1
k5MZh2vQFxHpIaQpU7guBQ0OnJcVBvvphtA5Osk15NcNGnMtGygJgklUr8CvN2RGk+pQOLSpmYGL
ftSqyPi0nFqCYXy7A7SjwMqJwojlCgotJoaPqOk5mJyO47QT0wbmMj0NWXgU0acXf3c4cKJlWRFX
20PhEFqKIa424zt8kTniS9NX/INy5GWh+Fg9jXxPL0lDoqMJpa0rjrd+u51JfRS8io58FOe5YNX0
rEOqfe0DrQeX0tUJq45JLM74acrDrdKu1OvNSYishxjeN/5xhcID5msogmJRW+KYDO4QvggAVB3s
HAi+lwQlWqF1Hijq0bYgu/OkLQZql0DSWoQMEy0R9bjYQsHB77H82Z9FRoTB1NhHKlosqaEHAXRv
tYOr8s5GaVrn0u4x0gY2M96GMt+spl4o0p71Z6EJ64jhu3SUHnBBQKZqX+QWPbVm+oAnzruSLKBL
WXlE5FujNSOYTpb0gPSSucxu6dcTrlRje9XU3EUhwcXhLkXurrTnQzu8ccXea8bGkxDVh8HV5rQS
qaf/igpFfW8Bbp1pO5zq0lQlX3mn+rMFI3ucSqQTQI9bU7nJXHVEpgzcyuR1X4W59lmHepBsxQc3
nBuSCkh2nbVTp8L5uJTraxarN8ggUi2De5sPzq6Omo7cVZo+jQ3iufsI5OY9bauCtg1gdSYlVFYg
7uibs73NB8rscnqwZ8IlGzcq/fJQXYFePCEJcbZQ2WGmVK3sEvlrXQopVnrXtgieFev9+9hBcbbL
YyfXblR5WqmI0YyvWumf4UX9iZmV+mCJ2jcFfagHB7F429ebYFSRRlNDayUHOSyNDGB4Mv4r2I+y
qjOwjN4YtgxsYHsP8L5wi+E+ieOPSNXdBTaXU8WQrT9mxKZlU2w6RK24Owksocm08krEiKm0Aipx
bLa4zcXSwB9qWQoc7v68KUfWUrriQsmIwMgN6TjScNx/lE9rF03CqzuUq4X3t28mnhNaEc0Ornec
SKnQHoR6in2MGNHKNzgSCBZ4RA1iT9iHKHsqDAkDlwdF8AsdIG8OzmmeZHiAs2Qf2KLJn/miPwdW
QRmWj//oGxdQNYwht5keskr/CYGPskl97jjUMDPPqvqrVBWPjhDEAeRtGIT4i/pu4bIyEAYxdrX4
eyqeO4Zc2G+Eo+Yf1yTbLzlaQXEdbuY0J6bn4+OlE79RqgR3L7Sesm6cahtKX/Dt8qwuy1nU3Eem
BlCsZwhsBzWAU+IwPyzXJjemw1FrHtXo927+pu1/g2QkM5ULxmZLv73E9sZgEeB3Qgc715ZSUllC
a1v4iy4rahNZhchTyzbFro2xJh9SSB/PQs/urvMXJxdEWnmBbrtaxGbLrhrevhNjQD6JUIMIISUn
Mw7b2tMioMgc4RaMvCPeShyPvVV9ChxXE8vbohOUStfGGqTOQqrSXGUh63CVIWH5dDH/GxSATyHt
yakBY1H8XJIJnmbr7HPr6as1J1apIhBUfzuFAXhm2/oLgEc8JMbWG/D2Kf+K7e87omR1DTFLcU6K
aCcYldY4ezeHQ/j6jHQLmkQa4BHRt3Z2mrgvUGoO6HfYqiqzJ4iYNoUIXAAgZnGmZXQ1ZjuGSRVW
gRRVhjApK1b6L73vhosN+Z5lS2iOiHiz7WqxOeSJG8sSH1ATXiTB6G5XCSxHvmWe2Q+GZmhU89Dj
tt1VCNSKk4N7wSCPUtN+dDYSRTvLQgxlLO2FpksmH1h8gqkV353QveVp5MGKMdBs7FApYs1tITM7
huI+ufWh4D11EyWhBalAraZUtand9xjX9r0Zkk8BBqXUBaywt81aFRT0SHujcaa5NyIuWRENLRGh
q1cJYBiZ9YaCvkOZrWWaXb0nAvXNlBqOODiOcrDsJAnioB9yAH2qGMQtSdNmsgbgpsm37xDjCfg1
gG5TlFA/cw/l8cz26VelvRzS0tk37epn0xrI2Zw1SFwNUj7tUx8TloRGfM5a55A8IlvziMq4lm1U
66+YLAXBiUlXe/WTPX6TRk+qSp7ZQ4Uu9VBl4obeECvw0bTn55CF6DMunxupae8CBssOJtRbSOb8
8vrg2+ZklqeIWk3Ry13++f9zfc6KTMibpUa3fdSJb9azSm4Zc+9VkpehvxinHww5PDl9b5pH13un
PG2lJnKyYnfCX6zrRj0Elv4WtCC0M6pVH+gkxAXxR8BPz5Up0ur6QSGBSGq9zOc7MbCZlDAhcdIL
/BD2EAUBv1TMDaaGaJ3HwoKbmpUbfgQtS8d91j3Z2Pprjn9d98vHaawE8uTOxsFs2Ybcw1WNGwov
98hgUZUTwc4iFGBbaUKUXnM+sEa6ojviHQ1/0KlGa7bZ4MOeWy3HhAKipuKFXz+LN6117Xa6q8v/
4eTlhegngZmcR63iL7MCpOmQJHZtLYzydzmNvf/efiAsLhGPc1ep/vpV5Ac3MTaYaeNt4jU2Dp7f
yLMchRyES2Hb+sop1fGeekMleztEOym+yrrclXqc2+YdDIhn579mdrEp9k8cdNwxrkrwmo8vabOz
vBS5jrIdifl7nscu5+avbzv2rIjhp9I/mcHwJmbuAWBuwuzfbEv7zrPe5I0hr5Uenx3SZAxevsI0
M4cPIfUiqObt72mpMfmtoGDeFYl1JijtNQLtLuSQcUA4g6pzw80r9uFaEEQ9eLiMnLU1ZxVSJOdx
bRDI9vxAqZAaY0T8MBOTM1ptbHoBsIa6QglpQyHVqlKLHB7BLMlNcicxEog0Up+AlYfCakXLQh8Y
WVljkXHNfO0pYOv5e/wx6EYRdu8+sMla3jE2kyqB7JRe2pIKrbbpEM8BzfqogewNEwn31R9qKzNL
tkzB+HBKzEGmMOCz/drN4RdNlzz2RKpzZmNK7R/NTwdRSeyEDD8XPMQPOwYC//IUzWqNmgHLfhNB
OC16SUHH3Fo8AeAgZtezS2BOTKXuC2FyI1yX5C2MbxYr+LPZJQHlI+VRvwFLKnMnmuk+nEY7B3dI
XypZPPIL+RCctjql3tJRtvmXo/E5GpIpk28FxSmsmCvIigUQbC3JbcPWezDQBruBldiyTsuRLyW5
+ToyWy1pOIIwcf09GPr/eTLQ5Iv0ljjUolkiKIChKjBxoTbCdkhEQsVAmHIR91zw0XfP0YtuTrSc
hftqdLG/yMq9ze11hy71crstXBvlZDYK7d5YJI6R3RU/V/7pVjEB9rGDkZR61iCvRma9AArKVKCy
Zpg81HcGvVBalSdUgLZl/PZQupyKqP57qtNguTXl9Y90lUMFRK7/64bJXXb27ANSJw8RgQwvVn34
1bXzaU4Bg/DANWyJAFAisctOODurwk2S7k4Peorg0uCLj3rhDC6ivhcp3iM51DyIIvev+PMk+FFT
N+ue/sL4nh/CQaw6mLUk+WDwZLGwGLJELvkXEM563ss+iIN0AFrklPXh5o7HfpQz7zCi7SrGsRCW
jvnez8iDDBXTysgulMnYo8R5jAI6WRgk6+lJeVqNTrVVVD5IIHv5W46A89U37pY0pFsllACam2ND
nwm1zdSP5Z/ykO+P/VeaMCa8d+4tovMBYF/zlx2x0mWBw5mwM3yIns3T/GAPL7kQXV06A56r3iFi
P0tUPO8cS+Q+cOeDgC7JIj1ruiqW5nH9u76/14TRM5i6EgVUVXbLHCcUohDSRjhFB27Cd798SxJn
qs4NhPkhm3G8gNr3+rC/ltg+hMueAxQLPSw8U+BLl7YbGRKXsAGdZBUpbOJj5IbGaB6Ab+BWhe1Q
FRYIg7HWYkiImPdZxFXsQn10BegpN3+L/WM3DNDZqFITDHTrMYpFLv8U1s1m8ez3yVZw8e+PMyi+
rP+CtshNQWReYFERxgOv2lZaoIxDn/e599urtqqnL9V7CVSEicHXxLyxjcxHJp3MggZ3SVs2RWWY
DkExsGyqo6R11LDreUONzfgBQijEhUJX/RuEj5FoRSboJHB7fC+BiI8IpzaNJT1PTbTpfrfYMsm7
RjOOPkpcbN/IsCj6vkzQBzvrRpYzcPFBttT4ghwlKlJwYaTMWV8SVdgfHz+2jRzi48s1o0weYCbv
Rs6R+/Jzjmb9C/sXookeFFZDVpm+MccZxYBcghBKZm5xyh8Q0fPbU9+5yL0mj+kSBCySb1BuPUQv
39cpTxesE3rbujaG/iFwVSU4O/poYaLkCFXqYat16H0jFBetS4HAJVgNIena+rTRGX+mJwo9qQE7
NyZNKYL7H/fuW5zF9WApVivlaBEhJlgOG0bgysxAVJ04iota2cN4ZZ6+piWNxRdpCfwsOy5VvF/V
gOlOmzYXXZ7dw63biHuU4KuXuOucbBnDS7S7K97zUkAgequCW41x9zLxpUf5glojY4ey6RenOWrP
7k1NCalJiUyQlPAjvNbqztZKM8/RcsuPnrZzcA/ZNh/kxQIFQvTsttJScCx5NSQo/cM3716E1ava
sehnuzHLe5ljmQDgWs22YluVz7tjDT+toMnpeLJ8Bo/WtppYVfCnFzxtRZUU9rRXIusK36rWHhm4
kmvORWZjT5CrWavasPI55ZLy5rHN6J/Yt65IR9DvZpkRqbnvNKBrjkOsWP1rei7rdPRFOnw7ipEY
HmMewFcjnjaPAI+GRh8xwM0ik0H1B8zLNNgoyxLRf4l2mmn+Vt0neI7jyROkDLZzzuUqsvb2oEEo
Qc4YQPGzJGRiHlaE4orUlj/liMCcWhfUXQGLfMRBRmf442toeeqtFALxjiZP3Rz7nXrKT4cqOAaP
dXMK29FCsjKhpCJDIrg8Ng81pUZT2kcNiQ92Lb2SCZCfgdshoY0oY4MwIbuTQSIuMXmhL4m9rW+3
GvB6jvVQgOzgg9kaXk2PXbjLyte9AVke3SjqjwIboUKsBj2t/79f6gnf4WQpr/9ZMnxyeUS2zbg7
yVmpflbrLUxjPuGpUoRlu9XrKSumoRZ+e0jKA0X3+4Bv0taQEvpmxfU2cr+sTWoNxT0Vdr8JPpH4
gIdKoKravJR+4VSTx6nswnzQMXu71ZSgaQHGoumi6d9SmKVl80ICMXqd0YOTS8+TzmTkDcjkKWuL
4dMELAew0NEIxg/mfdnANAN0ak38rKh3KTt7YgWZel/vClqQgIxFyq1ImulKDS9VrUqc7T/Do57u
uzwWt4LJFmnGMHFjcE2tFW7+ochuZvzbI4TBYrWjC83uQ3cJK9akxQObTNiWgESDuJaZTXwofEjw
8vqbQYQmPgi7qeckk0KCSbIEL35SX6ghug0+9UJR2WBNcs2+dVO46Df+d6JdvGeNMNdh7YYXguJQ
fBuuiHz+RrO+vQUAsI+NONDJfnjvYBPYtScoJhbaPcz+IkfFqNkkRdOuW/87CXQajSSOGs2wK/mU
NOo8mNknANG/6ELAYdC9aY8p7HxpX4fn9WLtTuuxNEEtOYCY+PLBdeFd+Q8kiWT5oE2qGfcbYkee
WTtKQUulKcwNk9AEGajGRZPWz6Yo8HkKWYmE+Q2jQHCk1wIyScCIL7wCVVnvPaSDkf950hOKB+OW
np2O5tTwC+CeIYwikUd50bGhbRbYk2GYq0/eKkLf8nqPtLNuS8XCiiihcet5ebqtgFXdhTr5ZRDp
vLPrB0JCyQFgRIOcpGtDB+dSY4lz5yQTeugBzcCwNQbd0AGj6EsqrFfEV7EDoBPNSjf1g4pbU2EA
V8Tph6SqRq3yrGZQFmUaeOTqvcNCBNTapcPa9/6u9PouU2Jcnx9ht7pKWLWFIBc2BMJ/BNhz8a9s
He8yEumPt7fU2T4gKW1mi3leujyx1YVPKVoFHB2a+EsVXJq/gmsBlOA7NslFggUgvOeLi5U5Cmln
jXQqorx64dH6iXmIXFeuuEAIf0pemfvk9NCGzoAsIML7mNP1m3NX36zr7isabJdo8RN+y+ToaNzM
py6McqmKX+VdlIIgVYfEaVLVZfcB/aCMDHDlmZEb/aCsjrZsSY0JfRNsUfEen4Zh2/vNSmDvVUF+
sPg5s/MQyNbj0PR1qnLCcvbmoisVCLy2zAOFGHFBLi41FPtzBNRr3wSDxZrQrxHq8z2vAGfMyvyW
viq6TRx6ODGeoa92/B4rCdxHM0up8ryLE17sje7LxIBFAm1ozazm8DOZIQS1qZOPuLiWQcQ1+Qcs
2VKdn3zjFGDjzxwdzJ/sOhJL5UXBhHAS2rhNg77CG5e13EIQfNx3sDekIIqIFk37KHwhM92n3MVL
l7DY+zusiHzqGhnMo/c07MTMASDL5NRXbLpv4fHufFz0A/TfKlDP/Ad67AYJJ2O2FE++285n2QCq
Kw0JfRvvFYYWYfcbbiYEL/0DgSYkujQ6tK41of9itz6kobGsTNvIj7cnY3gCb28nccZLWcptbCuU
62U2BXOr9rXvUec3g4vvMj6T3oRdVqOo3b3EB9rbk1C4F/1pTmmKKXvY6TRc1TUHOSe9rcGBHOnT
3vYaUyRdELhwWU5NdW7GH1PpRAta9wOGvqZHs7D5jaFJQsdplssQ9SylSr0FhnhdzBwfgfpzK4iu
cvishDe/ebHSrU7SQoSYvysrkItfDtnChgOGfm+3JX1H/tt41/XaTBeW3HuWlw8LDvOXQhGhIt1O
/eP5b3cft/abWCpu+XJwo2DWKVznZJqJbh+54EgJcozQEUKkQIXGcojeMnmUZzAd/EYAZIgtELR4
Uy6aHaT4F2+Zstgug5KF/QlQD1uqyPI53/P52krNoj9ad5F3+t5L0W47gktUnDQhB4WDua10KMfG
e90Uly7Q8y4crMflSL3n6SLrTByU7FIGG7UrGrO6w+UBoYW7DKRQuSRTpP3auy3id8FCpxOke6+/
E6RucXkTdp2P2NFBsv8SWpfTFQStp90XIFOiUd87526cO9B+SvMOS+mfVYwHRhqWaDv0UZHOT8eg
FCB/JgQ8Vtlq/impolPmy87Rxl7LQY885WFGfy3c/EOXDuYKbtRdZgUSg0XRuDdAIp5xPVSLnYBA
5vVHCbWqXFKMNAsrKsFVPfulDMstE23uwKnoPf5/tyMZPgYuLzkpsvOGrraG890fBoJEYZX+ydRv
Yv1mPmwPTXlNpQbDI3Aqkf0ln1wURpNxGaAxwI7Qg5gKpXjxzcDOs+hZXsiA2KpWxoEV+N8JE8Zd
aLKKEI5iDPX617gEiDJ8n+UWBIB95OkH874+kyTRAN8FEfdo95QHWL9qHLRBl6u2+HkPG9uNQpNo
GTkhbkrq13TU8S+iyySYI57/znO5pkM81obQzl53/NICgX6O7gPQVaDw8cQBmwRiK7qz8bYiqueL
hvmlRFI9dfju+gi4iZmnvFA4F8T2+xfRoGcMa/Hgo8Vw8Ikq9QHsCqV47Zc9H4xgW03omBaQnoQ8
vity9mEcgfGIM1XEzYIXTj/EaUR6Dm0vUmfJKwAf9fZfHkpeGG3LBPZo7v+rUsRlljymJpDhIOez
cVal2MpfYsJ1MpkpZyNLWV6APbKS8L2BZKsayaCmV974mN1nPAH+FZDiWvAXM0jQAXsIAXIslqi6
nS281YLybVZLZzMuPCtjGgzOgGeabqpWQvsrCqI23Ak2WAk2P2y6AqSvICwdx44LrB5VaI+gHpx9
CKyBFodpDSxPhRZ8HO+J4/gXPum74pDInthQ5SFpMpZvuDRlnHTGtNEArqg1HGhfMxh+KccM+1Kk
/5f0ZgU2RZ2de9rn4dMqyQwb+EHghCA6L4ueXedBPcZaNowO2Ix8iT6viWbksLUPsDReCsoNhFAF
esRVEcgfEQT0quDfEYi2ZB/bosYWHa2XMePfHmVq6abqR0ME1n0uxrWWCb2Ls1lm1HSMYqZUYrJh
dULF75r0e1iZH+yaw8s48W1EhWtkSf20/w2HDO0hbJKg1G44/2AZc1It7UZntwSH52CEoUz7i9Ff
i0idtAWHBwVqhW+kpMiM06uabNnwZ1v5rmq/Y5C6qlfYPGAfHM/7mqFtNV26QOFsrFdnZLg0tpiQ
me7QsFDjJZbYxxJD8hjFdPsbArCEQYOdtWqR6kawA5D/QfJjBdr5g+OzKCGHnR4QzTlQsQ4sitR/
dBMiCYf4nzPULk/19OvKoWVWg7oJ1Y6yp3XN1vov299rPysfAuNqAMVv8fWIJCgmzMobJw7Silr4
QaARfk2QVgkwCCdNhnHSq7bLVI2tD95V5zsx74rsUBHfj83g1N4wH+mgvQy4KjFxJbtabfb1MZh6
gmeC15GuKsNJOmnTRw011maBryyMhFfWp8he6klN2uLO7K2Q0nI9qnwRnfkSjtOvf5OoBxjyleek
LoJYthFJCx/jK5v1BLtb64D84XBwSEFk6hX3H4+zflqgCnYUTH2uWbXapM0P04YsAmY4L7UvoRld
BpF7rWDayfo43aznpwvYcB73AOk4XO5pnZTVg95ukscME/Y6gKWHtx4VVAWl9sce4g9EtENvLXLo
QA9k454dXCkpHFOyiay7cmOToogcEDkRoYSxRT0F/Xa+N5WlB7iPpNrg2E/Vz+CzpdRF3+L205AH
p/rMk3ruOjJx4EdreOXLfvY8T64rp1Dz7qTgRHyhD+HhrmXvfBrF/dSxjw453Z6Qakzdly4UGYpX
MbV/WrUAhYJugF7jcnMAbMgqI2WPkeEYjw41viEJPyxaFhg7q14o5eeXLzn+Z7cIeNNSZ/DoB1/K
A6J6Y6838SgnflzfPDng1C9nSJkZlVhahwMAjMnOYFGTCuXRo5EN2rAmPudvVVdwOWjkf94/K8vc
ISCUuSKaRCKBR2OJyTZfKZL3IuhQvBkt0D6ShdIVqIqbPsftN6VgQJaSvhjg+XqLp4OS1SY0j2Jq
n9mD5P+6lZud36azblDjHX3aEg9jqfoM5vM9ZBk2EeNtI049bilajAT7DFQ+i/Ie0YecgGg09r5j
wuQfJqnFSmWZpVTeqXM+HgaVmc/GudBm7bOED2nyEIXgkzOEUEuYq6JzIpPJ6ZO5/8gEZap7e09h
+IgWjGbe7glkmE46JwZExdhA3bA36NGVtBKcyjBRyL4OnGQCUJTcimzzodijbcBhDpsVqGsf2W+4
luSWvHtTq5DI+N/TgnSTto0BC5ISvRZvJOZQCp5ufk/qnTBMKVeG3yWIBjiSONK5JoICFy6Sjn7C
yxAfc2q5AE5cNy5PJdZbdptT5Gai4jUUTuxcFe9j05/ASPprDz8T+7R2i8+KR3/j0a7NAys3bXNa
pLctoMTuyfwwLEnCxlvW2Y73FD07gee92MTBJlqoU5DFpeEqja/+aKiS8GV6RI/dFETcf2YmFopX
0zRLMS6gsAenjhsWAHdNbd3JNuiiLfKDi61bsVZaSn12RhEzfyfv6DWQk4NQLUDBKscfyUPHhwjW
wPwartJE6RP5TwRLsP5EzMe4Bgn3SiBDWl2tuE5HhuTTBCqnA7IMT/6/GUg2zwtEoLPk96U8jeEJ
06Lw5CpOG1cVwc16iscB/mc+24pN5yRkeB1rJ2117BilRW0t88dcl8tsiEW17Li8MahI4B+JrOyT
VC5XldYa9fHT9H/z+5382Ql7WXB5WYU1bPQByLmUNSoemD6MQVwfVaKyjgj3v1O8Bfwo5siKwjvP
iKomv+DxuHIrWoB5MTvQwuamfl+8am17c881Hl3Z2Mqxpkp6nPOJMwckJ/GBimtOJ0k1dz2V5O+W
B0IS3cNCKnT6D95OAJ+RDN5Y3SEoBbBf1qflmHoMUDpI8pJY2Efe8uf3VvyakBQG7pTj1el9zUjH
xPFxD7C4ZPTrCB0d1/M2SBA0OQTSdrCqt9updc//F94OU2gRzYhMatT49tuIHBZfEZWMZCZXtJh1
D9Bd4KYm/WHIVv6pkZ1kHx4ZKSUcEAi3zOx/4ah4Pp3jAdPc0cSbN/0Bl9iC5Pb30+TxZmpkXJQP
DL1n5Y2aeKvbHe15Q3qJjTR5ZCk1UP6VtL2PzH6P7VyqFZ/KgdUw9GLSj7bxFYbylh4roIGCpAzz
OyOLQoyddXGhln6V2CtrimUJVj3aCZQrLwR3ngQobR1evICwRfNpZt0D8uET46ttoJ+raEyUNFWS
+nzRx6bWrJD0F1I16xPrCUy334Fjjxc7q8GwgZEZcUW2kKGIBcrdS9cOPkWu7hYofqFb7cOwc0Xu
meOSfWNNfYquLe2b94v9zPd5f+LVrFQrQhGrGgaxy5PSOYYtZdYZjIvbAJyeoRW/Gl3uSoEdO6Rx
bEGX80h41sb6qMKU1EzGDjA/4Y8D6LQm2gDHpDKtI+K//beO7rhSCQp+3ViFsHnBq06cQ27kiC5N
+ilGbcCDzVDl+XxH9n5LFaV+4maD/mFgqyYoRkG8f5mu+meVpdpuqUg5ZQi3n0Ns2qxhp63QQ0o6
UntR6UsWZl9sYtF1FSsRIjge27TMuwJRsR5pBFOXFvLsO5XHRUuJxeC/qK+yy3/W/AMJd/i+HDf8
LzPbf+tmQHtKWL42AFm8X337695WZc1EicwplxYZVIYTnrWdoJ+IfxYcq5FnuNJK/puFxFRscw5f
xhVPC8NEbVrH5kJ+Of2zqGHq++s37s7w5Be6jO8NX3wJ6ekcoeDT14MgVNWjPmeh2q7HYnnyKSma
Cok4HICHFHTAyXYejCx/Lmgneclk7c2Q9SW9vRMSPuOcXf2RYxqYfJh+DF+nGCHDG9Bnpjgff6e8
kukuz3KVOpId10NQXd1vgji68LdtZ+noJCnd58ZD86+ixXZ2xIjwI4sAEgMnlGO3KCeEffqFmOnv
bbta3PvbUungOm9LqRFKaO9E6sZeQItkT1133PwjZ5MVXyOHa1lrVQELpbFqW4Rr5Xtpyqd4HDcY
+J0NV13PO5eCZOKKAekCCqWAP+hZsyet33fE5/hC/c8IzLrno3y3p0sb1OG/NLoWFJWa5crFhJFq
GuQ3X9JAZ6tCIrYiBQhG6WXvyb7GM8uYNN7COWdu+vKg88nB/wr6stvo+KM5nnF6V23W7/W7bsc2
bmKNvWzQYJBeOaQovu77sYj1qeTXwBbzEZR/ZGJM+GkTPUZEGUj/lWwDokJxbHCh4DezaVnJn4Os
e6+B3sFuYVudOJd4XHARKIto7GeQFQg5vrexurShXWXxleifrY9+2umyeG6icIoBGZeZubspk024
gxR5ZFgwTQdRq4koOxoPhmVpS9tpw+EHIOf51/sZOlzrBj4LAaZQmJYOl05eohm7WQfd0GsQgHgu
B8h58qn3aSDGJpJDTEmEp5IwjoVIIbt7GmC76P/MMKUCHbuUR62e2bW1bp5GB4rsUwZTJkSdOO3j
RR+y8yXbGZMUKzbgRNzW1TBc54itPvSaVPvONt60aMyWhLKV98IOvSGx76RtSsvDfgJ+oCtOB6li
IMf+hBBPycl0q34yfxaSaEEW8BlyuDIU/gGtY/Ydy29eDZ3aNms7r+TOwe0GI9U/DYyLKzMHe+LU
TIHz+r/+w8LTahopkx+H3pwDUSP6N9Dfonc/fhchNSvGP38Qj/zmEmHcU09P/prccvfu4E6z42lv
pNkj0/HmhUe8nctVKyNO10rC0x6JpvAjtoC3Pnb8xcaJm6T8OAjVX62yOiLwZmzztNQrFLJhGRz+
zVllpJNOw+/zOYfAfndHLqlC6tN8ttjk/dQ5As5NAbW2Ei9QGW6sQ8n3hM+BVLkGoGU2Df//lzwo
GbWn89ruIclCeo/jydtADdA+2UQgFKynCM/ngmbdb1CoTksr1OjaHGZHmltkNmVr/VO4pMCDXQAw
ZJiNKL0SxXS4cG8f5HGzX6uF5HApRku6Q6Nn2svF805l8ABk5kWCuZ59ydD8PUvvPqSHlnOJ6P3g
uCXqLOtrS7eE3INCmwBwsBd68JOLmkRajyi7RqExTm62bq8KdqOUA36OtJrflPRD1b5GNhB3rRyg
C2N4p9WNJ3mvyIRISE1dcFXfEfv/jN5UKAWTAD4NhxPXtaWX3zcMRYk8FW/Kicq98NxEKqnLmgL1
/IU7ui3UrhDl/VbJTw3pmEd4ua7rtIHAhdOp4fJUhoz7NyZ6BpTqsYLM/Pyo75AF3dwhsrND6Zu0
+AXv6CNVj9PqosaVBhD2ekRB/2vURR5bW34H6SuSD8CttUc+50n1bCL/yp5BIiDCiBCMZIlNT9Hx
eAOfSf6DFfYJzWLLJLDjVhhS7wRGX9fkA+SMIdkm66OIJj2//9xxZ+3V22NQSGTMWDLOjajpsVGU
axE2mTdWppj46B0x2x4bV7+8bON2vqk0EIh5FnO/AT9+2Y/HLzLjQ8XvRTKozAOkVtkEFwfQ/8/t
MjOUP4paElpU+uuhdU4tP5UqudHExuYEFxdJ+zBdirNSU+1hdAaV7mvkUhEcaPZVKm/V+KswmJLy
kdekII/C9kB8m8u1muW715TXfPkAXOpfvi0QBIq+BoCtkDduk61ZhUKshMuuCpGiCd3uOrsqz9bj
hkGfplS7y/rM+6X1seOWTfLs3SjdC1z18ubTEKr9cAUr9jihoYnhEsyIMnqTOv7sNbfGRuc1r/hv
RdFDqBiFCSJBhG+6xjqyu2hy+nIbMJD8oKfhk2rOxQRamd0C8jSwboFUZ7yD9mJBAezskoz3Hcr1
WGScOaM+IquFxH2K8jpkrLB2ug6q75mwspfZJCiCfPR5g75AuNg3FzUE7y9MKZGIwcqqpsohcVMU
L5gGTUFGtqgyF8o6Cd5fzKfIgNkbq74OaXcJPbrDQaYAZrq5nf30z+vNX3fTGALflxrpdsZTP/Kh
lmRwxoz7gQtP0LWdjWXAsxTcBU3pBTxF1Q+hP4rCE0CrrVSJit4j7QZqzhEx6gknUnAiInUiVd1/
U8obo29P4zqIGWZ+7T/j0gCuC4smIb8c7YL/XcPZbmcPkWP2HvY7mxCkAX/7kplFRt8fcKaewTnL
tJOGFJsCKSY8KPRw7JqT2QSsOIXNzFGOAAwe//8TMnYmszA6ywkBGTjIqhY9QFoyTrfrCx9fpO3F
JdzWZXsqvNwRh8N26Sm6uoWIhWABC94AtTAdgdgrU7+xqLUAM/cZr5RtKCQu+sdN/h3Ff4Us9634
7zKouPxsClQ7sg2uTQXqpwBjhaSx4Ew9jJWoHUzWoSD7G1GEUhcs8XIFHXcx5gAtPNq6IKVhabQW
KcRZ0RoOnN2AhSLVXXY1XjLhpZhZXg30K5PmJ4CFaTdKPbe52kbK3wQ5nn6M1JveznSTe3S4H6s+
CSD3vl8J0b9kDcRR+a0p3VCWtghXJXUjcQjgY0RIpW8ExyfwvvPkiiNtogWcOJPapasssNEwHvPF
kDaP+yAGJtG9pS2vbvLsy5T3mwHWUYHj6rtOEDNFX2hwlo84aqhQKsLKcfpeVl4fTCnIWKf9bTLJ
aSrpd9o0guMvPtq8uuNR08J5iejw6IIKvUSmDHWYlMY+QlYJum9CxDeAlpOV2QtUyLdGgQqWfEKR
R307z2wicoBiEUNESIDHSAX5MM7jMJPKKH6ef6kSMW4dYhZMqPXPOmgUQrAA+DOfB/wdeuWtYfyG
2TUerudPJmGnPEccQoObUKnJMsEA3BN4x9YsgnObJi4bELXyeMqKOhUfyWPNWQ0EaBSXLn8gKtiG
j0hYIYOqZSsSNcD6IECZfK4jkZWJCBcKcuKKxiRv5feIJcwibljPerEUj/f5dYpsRrshAR63cjjQ
8WpzRs/wgxctKsWwFwdOyl9PoM8SqCc+d6deWhfuEI+PtGS9rJvIUbJ9Ui+Q/Qz+oSmDRRDvBs/w
G0FYV7RruMihAwkKZigqAmG+tCZUMpAyepYnOuy8Vq2tX3kEEgiaT3wmBxZM1Wpgz45wFCRiOpqX
4+wVEpfGPQ/bouJePNG/nRPE6MXts0oBTNsuWxZ7kFa7W6IRbhIvMZO9EhBoHggFIe3YAxmupUxE
nEnnIA4xZ82oK2HyPUrsX7cbt5x+sq3FN9gsAAEVD08YAwgDQoWjLS6iL8bjSBYFo4+0gWgQwWax
rpjepgylMexbc3/M20LJENKGRAObKrEcP0jlpGhdS+IriLQumCIXuNU3RZYB1Jo4RbS6G8vL9RKW
Yla28KVBem5A1wu9zBS0ZgQkGFDWQfC69EyChYQvo77P0YPfChWl3TwTqv85uC6sIiLvIW/tiHTY
vBhAimhvTfkE67QPd43ylKBOByjUuyGj6+7Ae6dRP/9Kk/HnA3SweAQbK2Khk9CO2UpU1F6CYLTz
NHVivpqPLemXLtUZYMV2f3QaMZrIBhNCs8XCSFUpmBi4MuAjbBqJUQ5bVDVn5b0A682ajSAuwciF
oT68Xq2Zl8Qmq3rxBZ3OLazF5PXbO/XXB22gN4yJJyAYvj8Hpp1cNz/Tl8k3dV/kwRH2i8uEqfmw
uJbuCvVgg8XtVqXznUVYFphVT70qqlvpKw2ZO14Hf1QPEOzGdmWaO2Mw3UsNPmAkr8dupnGjrisw
5YrtJ2XEDO3SLRDm2x66H+egVSfYUR8axS1V9PotW+ddKZuqAoTy52xTBJePOoDWnBHkzDQAFc3Q
9cx3ov6FUpHM6rXo1+XYHquFNt0+JFqkLfIv9BvjYtKmpLpDF1u/p0BFjLwdjnvQghfrrE22yGDw
XnCZqcAihX5NsrC58FX0nWhb+ONlo+pRWCr1t+jyUn7Lpix96GdfEgpFO0Rif6I+Ht8jmHhR1epD
N+wkRMg+YEHma7On1DDgAnh0xFh5aFz+Zw8sufJAiw48e9W2ybHTFp55tnJUEXEHpNe5nor7SsrN
yfBFc1tPSU7bbleGuHj9dL7CnPhzvUNnYGI5s+t3DvDh94tNCZpyOGr8z5PPOj+5xs/kBJEJM+zT
/cwELJC2CBRnKp0D16MtcdxSXlj7iJDFoPlvhkadhnkSE0GRTkSKFbf+vNVgSNPnA+cBM6aiGMIK
wnoBrpAa0oS0ghmHPAYft88hj3Y5A5WZPElPyVywCOS67nXwWe/6jSwZoDX02oK2eiMuOkrqnW2p
vJ73is4nLJWQHzip2ElmU2Lz/L5IpbBbt4pxRU4imLe17VkBo8NqIEf6RQfv60ZI9FRiK2Zv+mkp
YfcHpP8clk+Qx6m9WAyFlWk+4DVGbePTBVQCpt3kRo1GWg5KQNi/vw6pB/zDsTOULC3W1ZT/dMe5
kwQLpQtZYTEVGVfMACpCr8ILRyBIL4nRS9Fh0VTU9YbHobo6chfMUogClTwbBJA/IQpS86idghRL
Enxko2aje3KoNP+jfHJNUiuV78cVHrS+BRBLsCEXsE8aTnO7h2XxAPsW4ZoJR2Spn0wjItvqaFa0
CcjoTIPoViCCk2FVrryUNWZp3SQGxmro92v+P1OIJC+YLGxX2Vy21JbWp6CLj2ix2Ei8xE5Zkg5K
CmOLvFjLAv/3xK0+mcQJ6v/QGs2l/sdKU/kXSolt+3NhnUu9ujpm0T0xROjHX++TGdYxcBCJQCkO
soWTbiRuhRaSmzNVIAkbz7ilAMPWUoG26PSrmvpCYAUlx90YNYnuO+SFEOh9oVwROPWjwFUXztv8
cZs1+xAiW5iSojjGm7I//568k5hxVJZnFtVQB3fzPnXFHBJ4K0EeaUgep5Nk+FcxTQFZq7oBhn4z
AO94yN24U/eQlX9iM7lGCMgtKOgrTUtS+/op36in7qY4soJE0osUSwKUyduuA3wruJpunxRDKbFk
QNfInHEDeRQcSY/MUt6Tfddfp3jL4fA8ZC6RmVpeb02vhEOn6D/9bksXI/XSF1k1AaBBWUc+PM6I
dFZsGfMh+i/niWetU4grvrJbGo+HJwi3/kuuGKvZFETzvhLXT54iApFlWXhmRmhy3AHDuUd/qT+o
1//k3XqiEfhUfDpIUlTiyoerpb80uzscXFIgQfaY+1mbdinYnaDA9ZSQr5T2RCC66Y8fwEjDAjc6
G1npCH323AkDdUl4pZr5Gb6t486Gwew7tVFtsgMMEwb9ZRDvgd3EW8dD9WuDVbrF2pon4U1cDLfo
re2DB7O0CAUSyEdJFUEM7l/lkbOnNrqRgKGfQowVinGlCzpNcdKHScSrGI0yEcU0Ob99fN70X6+I
sk9VG+mu1VNwGS6/bT3U5UFrhsnPct+/IZ3KpVan6/KI0LVjkCO+HDiQcTCXWzr4Q2xamIuW7rq3
UgTWjzm27LCd6j9NcQvbgonK0F2ketsotqg3QKwiol3ApB3pF4aT8Xwr5hgD0l0JqZxwRO7OWCNP
CkeD1qNjFQPgX8xv5BgFMdjTfL7fHt151tok5ffRBYbTNpGq7GG227n9h78267UoqcRIPRXZJ+rS
NdEp8R6rz+dNSnZxRXfi+H/Lo0V8un86p0n3GkDs1jty5wrdInNiUmtc7iiSImcuxujQel432PWr
9c0zYLqPl0Nk5FDCMEBGUHpvC5tY0bpznfA1dxfN7lakH/tAzzd057CT7g2DCskHZWHDGev6i+MK
j4RGGauiIdcFwg4wV5N9dKTELge7yug8q3zPi9mgeD1917PrTevb8UimR3wXxC8vS0uYiGKutUhM
BXxUDKf+R7CkTTYnweuErp8OKDJzJGKbfHeakJ+51Ar93lLuw2JU9hqg/LRSuB2cktBAJXwJ5xB/
MV3lxVqlMirlqZhC88fa5GLn488K4A337WK+dXAKzFVztM9fcJBCS4PhatNQH/kbzz5JzJL3Q4SX
sRlPJB2CpUKTXnnAciZHLM8vk5GSxyFy5t6Gewziiy/Cag7O1aJD3ZQZM/Zm1/+8mjQzjq7kVSyO
HdBsIvnVQwPar7EB5sud6tpjqayyo81QNzyWGiLy6szev2s6ahbMMM3CJh6o5FRIUZSsJPany76l
/DE31F29OrcHmZ4/WPuxzltM5xDkLbgf6TmWuWx4t2Aq8mTy3dLOkIFXNDFPc0MLLdCwvKrBNoax
FVzlYUinB+W173MrxiHocpLxqjmShd0wOdrW7qc4KI8qo9Y9jowQqx2Frx++jSmZPEqThg3I5c/R
RgcUOAnJW7HDr7FBSYjMlSUQIcOpw+ug7+Y6bSAmpJc4KQ91SUwjdlBkdrAhlw9LZCAuTxvs0448
GYt7252cT21r3PfDPPSWooV4ukX+iwBcpxMNOqFO8Qorac9MDr+cT+Z6MWhR4v0wBk4kEWtdC9x/
y41O53ACrB5M2Xvy0JZdE9wZc1uQD3dTFfnpLaDiilOGSr6Qg8DqawrbHUoImqjchCCLF7k77nQh
Lo+rNmLnuLfe8Eb5VPtn7//vpS0Oe26heyrHT7c+T2ocJIPkY3jOHvfvw1J77hB1XFco3cI1W6TN
XQm6ZtwET6iaVjDqIKHQYt4huc3dv/yqOpI2jXHT3qjFCl/hd55NiDRFyASTr6ohCSYRUtmkkACo
OboNjECybNcypf4KYraleag0eZyYh8b+Y7QaD7Lxy6V5ok6J+yR1wE1fvgELTXMZqs1L8W5sO2Pa
LtDvmt7yj1bpJRgMl3gB1X54uPrOmJt5HSyF7plt4z+WgNiTGo02z4xonwDX3FcTzywvCvf6uA6W
7KCQyb6sYFkmFykoIyZZSxirMEnD1uEQtq78YfL04RTuNUfHuspnO3tIiVHIsoEJ6+GEmjuWcCBV
RmA0BS+ndOGvMlHVAb1BLeuY2uljkukmpU06K2Te+sXJ2ruOzulr0g7ynQEda+tVnlqDMvpWkLGo
9vgF9S7S1HskZtUesOfx7smHgfhonJ7IaAnNIrxAP6wpMmnC0QtAR1aSjj6FrwRcHRNFTc7r5Ho0
yS3xvTHiFZ/w2KwsuqPRQ82k9n/r7Phb6HyUlk/qFC1mvpj5qm43lZRzlEq1a+OLVCOzxQ2CuC8x
cY7iG89y9zf8fFnSXH2lh8X973mDeVitJLre4ciulfBaV1z8qn16uhvjScXwpd6WGAKh3jKnMBeq
kFgJMbTGflX3HBCBad9flLh0jfWJWXoGj8pNOWJlttH4gZaaOnm44bBr4IISHmJKBwDJ3W8YJxqM
daxDzdtHva1IatrXXQHcuw1VMS6WC9TyFM13aEaQSkiW/Ssq6gFUmSNsNTCTZB3DO7TNCpPeAzNi
1607dD7jC2SsoLoQ2fjsnwlfZD0rGZP8QqDtU6Nl4W270bnFPyvRfqRLk4tbjr8LMVxlTsc0QdaA
Cdpjb5NulMBhHUBgZDrzUps9S97Pcqnoo6YT2glnQ/QjEx1BMumZdeddCBA2aG6cis8at/wSabbJ
aQPKO6dfGtcZuQWcfqAq/35JOw07T3/N4LtltlLwcGAkrY+Jcde7e0tu/4zAv3mxfmxpWR8UiYsN
y2WQdYrjoAeioDJWL6vdDJxKGfBMkRZGIZCVTcuY+YgKWLhhfx/vrTgqKrl3Pies5ceeVHL6d+0p
xr5NA0gd1lmUPSrhPuRcLKpTewj8oXRnrcdGlFHbet9GtYJDdqvFFMGt22X+73jZG6QVKUexQH49
tCh14cJ84Lsl/g7aVYoWPyH0mVD3W42PT9ZyHTsLazOOgT8Rj+W321TyJN5G7LQo0cQtk6tJmnAu
05TsCu/yekFodSjlXOdOnNiu9yduiiFQNLrmzWkcqxxFZvyhXPfCwIKWczMfDPMCyAPi3Luy6Y6S
W7oRbOP2OMHwFYbvai1FQ5ogWm7LEAKKcL5eBbTsw0Tfb77y0TwD5Yj4S5+S+KnfNJ55uiexrosB
MViAjGO2HZl8LKIcV1cZBLMo/RhlNRluei9YOdqIbIM8KEf06+37bsgT2MjhhRDUv8p7bva5qpq4
MfGQgtoe/4j8Ps64hJIl0Bju20LlZpE5HAnmqI4DJNljIEglnk0JwQr6100JLpqgIvzhfU+XUvKM
N7IDZ97ZNo7y91AwU88jxoV8mEv7594Qnst+9QWz7nV7Jbq4r0e8KngWazICibrX6oFwchRdKUbe
2IKFFc+r4ZLZRxuN/3TcU5fNWgCb8ENnsg6GWajqAxQtSHnLERQU54NE5Qz7lgdDQFbAFDWIwJZ4
7IzlfDSJyiH214ZwCk5essg6qTA7NN9tUwwMBHmj5YOQs4Flni3yFM441Q0PpFBG0p2/9XFfu8ZG
lgiyf5WivbHU94PKG1ILd7LOM2CZ+W9Fp62T0TL1KdoqGKip9JsmwEl/jZvvxxgiIVzQGU6d1p36
LjJw45hylOR7aZuo6FLaeQvWYOmcw1r+ewkS6uU9vDQOJ96KBXabSfAeGms1WfAElU+ZF4PZcqH0
flPmsv61L8YNYY6ds0OaHT2C8VQBRi28HyWWFOFO3ZV2eHEQPEmbsC8wkAk+6LfCY4xJPvOoH7g/
1vtvI5sDm35i2QjBPgZ1vUwaSZ2dpWmEWnBwliVxjod4JFyup2kcG16i7zqFDfpGOHsJZIe1pkMV
C2wC22EARQzNrRSt80boo114aFKBOd/QIESl7ihKUDVUs/Fr88H3FdYoxg5JPJWT+EJRt7Lm+aAg
mrh+RctsjVg5FzQC8ADL+i6Z/GclyS9sirmWBrxA82CIMtIKSbWLI2TrGSAM13vWDTaPnrYmLuKT
LjPI4Mak7no1564FIk2HoiOp1aOpH6oJ7X8no2ArL44E0Y7AdPjtTT3G0EcgLgsSAh4UxBwi2Puj
ASK//7OMvWhJ6af7yPN/8b2r+NeFbQqKoj5sEnPIiqko5XjjMJPpUMGNz5gCBTBRaluO4SxO2R06
AboXpgOCVG33N6d1G3gfxI+hy0yRXJVJGO8SCotMeGifSp+AseawGytE56Pr42/YvVFr7AwpCpnH
VqgzV0i5LzbPlgxQHon5ns1mpqxQ6hyc7Fvxl4Yhww+w+1F5DKGDPPxEid++WGbMLs1WTNNC3nRW
A1ODQVbX3OzXKRW+29d19HJk2rHZ5SBk+xPnN/mqTXnjEp0nK7RCT0oa0JwBl+Q7Q8MnjaET54UT
/z6UXSYIYwbX8l6XtD4mAPMp5dpXjDw2Ard4QhMvnT+TNbA+e9NX8CKmB1Kol0Aj4MmpFvaITgUZ
RFd/tOz1+bYL5pKf/F6vWWFZMgcSjNGryA1T/+YM6Pw47SA8YQBNV+o9xX+KKWBCaRToU/kb/d9X
Qn3xNBE5kY8qCgss+XGc/rRgimovnEheluRXEk9JfhK8E2bIdMHKsJmNjRAveLddFIat5dqwGcV5
pRmkngTYeu9ngLMt7PBlXhCXzwIPqqhgKN2EfsHAKMvcPsAYFIZvZTs/NyvgKLB99bT5/VZnh0OY
pUkc32qlcu3XqW/h9yjcT5+Xnd2jLtNY6QOzyTSeGbiCnGkV3u4ya6wASq9A92PZ4w2Dcv0D7/4J
HYdP5ypvQIvuglIkAfwg/JdfgWPqO2rBbac3Cl1b7UeZ0TLFI2QOUyn1rpWQwRUQH96bW9wAx7mG
CDkKjRW3x6LIEWFJ28krubWks34oaTaZOC9QvERFiz7oWYVXP2I4P5c1Bl5mG70rvcPQcG/vxL8u
uM9NjoWyPnNG7jDgVrhN/mHj6qZuwzUZ3wFIDa1EBEt5KbnC2gey5ZWcRP578FcCK3zI1pIl0iih
8afNgGrsdiXCeUMUK0wfcY52kEnCHh/ucp7QbdfLiW8CdaZONXjWaanxPDiDw7hQCLsQCDW+dah5
cyYvmqN4j/aQosKLRWlAgC++0XKo35C2/y9hiHKaUCgsYWNk32NYv7lzJaejrKm/AtRMqRvzrYrD
uMleHPdkxC02ci4zsa3cycZK2UClTj1aizzUlY86zzpYe8SBA4EgZTt9h3d5ErGVTdGtRV+21oB4
1Ew0clUO8UnT+IMdK100Tb6dYQKkhr2gPtY8DsrWA6Z5vBGKXEl9wmYcXhDcnQ29jJxmiNUoop1G
v3Oi8LDAvD4OOTYc69dTRpVGtmh4Uk5Tag12NzCuFkqYPvK4rT3zx0EdUOWABZ7fuxoOPbC1nWao
zJlyc9FFvPyXQU56pRlu1Ij0gq1TpQePS7m6RrO/50Vuf1/c7Xhmhh9jpZGHX+WJ9PRI3qEeM25A
I+SZB7Voyb3XZ654WpcewrytIP4iHqxMmIvR6Lu6+6f4Kgfo1VIyMcgQ2EgalHmFHhbVxW2wiOwr
brv5wcjUFWOf5mXuEOUM0gCfvi7r1NepoEPdMAibvH8lZn9cVVhcWzbzKLmswWSLGahG8xZVRUhe
RceiKbwdypdZJNQuaJt24jfMvTix9jPX2pRPjDoYQfNfq72cxlm8pKuv6snB1+Uj1grPkJPFhEA0
4YZEkGbr5QdunaUeHNvCS0gA7OE2fTqpUIKTuQAknVn01vDJsx6VkCiIAL+4qmFTsLPriAs8uWGA
lDF5gvUJgJWQ4oy7jR1ofGg3Jt74SMDLRETxHHiOYu0arfDrViVxpSEknpbBLDe7R4eGvUYBKNaL
8h9vYwlzA/yH0V/Ce3AILuX17C/vgSyT47Pl6bDeLGeV5+8X4BubkxHDDl++wPpx15lvgMHc8BB0
0rjEmycS5yek1Nab9g2KtauYTYO0OPnH+cjRx4BNhWRzJWbmvCJdSQlkPWZS5vj7d9AQrRaFOHrr
ofZbmIF95Gzpr2PdSLCx4KysAIss9IxD9h/n7Bpkcdhs+W5xykD/Hpx7lrgxiKELbsimCDYz7bwM
m9S2hwDCh53v1R3wnn58vzAP59ZKN87gN3YlkQGE5AEBzn9R1q77dn5SuQwpnvKgSmUzsczSlI8n
dQBrPveExQB0rl4pLikuqJrtQCirMS/NyD+j4Am/t2crc40nFMHKNzgdzjsj9PURm80rGdYXleJj
it4ZvcsHCQFcnuuSBVAbx/dB0hG6kGTvQqBRJD7icRnmlBSShsxRc+5/WAUd3TaC1h18vN7uB5M2
qnrV+tdirqPvG8PqUpoEr7Jy1ApCGLqkAA2lEKOn2jqDlOJrOwnFexlurkVeF+KnJzWo05rLsuIz
YrPtscUn4/m4bRg0aWBDraHpShQKPyUnln7/O4jfViI2++pn45LOabBdz2y2S/4ZW5eb5BK8661c
+DP0bkzhB1V9sf0lLI2w6+kr/9+7b4/t1uYYVxBcRyyNV9FrBG3DYFrmtaZmuCL7Xxx3ykvEP59o
OnJK8PMOa3JV5pvMvdHTUj7vV4KM3qa7s8Tg0AhcSw2u9laTxE/eGmqnUHzCikQK997be76Q4uOi
vEBWWqBQmy6RSXe4HJ45nUCGBH7CK6VDL8rFg1OOGr1al/X2UYrkxk46Ci8WHTAx1E93UqGkKhMN
DnpUbQllswaQ+SsFJPu/coreJ2OrB3IDWiJ3B3DzxP/Q3yI+pAzTDlC3Zt0hXGbWOFmmzN2J4D1l
3plgtDN9Bj7S6QxD85PDoZWeWtM68u9Ndiusakpn6ajzbWfI24HKahOTIKA9aQIyqPoRe8lq9fiK
K3CiwAqrRRSpJtICml67QlXvfUS7R1mpvNA517rhKysAveGpMtVyKl6Asw3FiQjVh+V/A3iQQFD+
18lSBysqd3Lo2fIinV0JGuGoOOzoF3ssmTaTpFag/I+VeOoh/WE7eIXcapACcAvGU6GyD8FWx1dR
PPtAZHLIMIAMV/BIPs3ORRBXczoByZp3zsQIT92L1b6mXVucNraws5uqCVceZuZErJBGawARHX8b
9QS4SaJOFFbDSRjo8SCbJqjdjN0qOKlI+1ddoo3eZsgkH8UocXOgIk6qyaI7NNKCAdYu1hO2+XuO
Y5vMTKgKNXIxW7KhVThDjiCK0433pLq+Riamg0Qc1MT9vayRUDEENbKdA0GVp0U8JttY3KbTFdkK
K0pEWyzn3rE7zIoVkiso/imOGnZUgJC6eSiaTUYdxcZHKR5y4b3zxsNFFbKZA8me1TSjgWDU59eo
RIFLO5mae6vTVEqdVjYQodIbtAaYK7zbbC4efD0jP63gCIuhOwEC1AKUPpLztJX+ImUbcuXz+SbL
b1Omo76qr938pYk3e8a+ziYRG1eSCl6WmliYM5ObvmjHEKGSpp4zwoibgRhiAt3Re12kCK0vrZJb
tx/Orhn1vnlNOkuUHl+xOHIXeTwSJc7PatWt8zj7WD38mHwJP+KmyJoz5ijf9ZA8g7TsD4qFZUYL
A0BLLJdsPDC50W5pxdvzdeCZypWhc6d7IOuyrPzFIzLIC2F5eL0Sn9PY8hXhV4fc7pQXqMDVFnub
TTGlO5qPJ5Sy7sKsJH4sPPle5gLWKAKrh4RUGwe1C2b+k0oo/bxNyvw5oVamuVtkMqNxrxIhyAnT
yXS9Cq+nQk7KRtWEEq+f1moE9Ri3FzkJ+bKTTWKJxDo2cpRzk4rZ8qIVwCXI9cfr/Y8V6wzQBy6t
Jzg0dYsr57/Mtm1JxZhUlRrbsklVyej3CUaYycPFeRQYvxd2iUOzUdAtt/VduxlWMUyV+HQ6VRvr
AhxDygiVizv0nsbf2qhb6ny5t3iZhB4NkOK4Sh5XpYgwxUcPkl8YFlCYEp8k/yaJ75LEGUraZqAI
rG/Hbjrlacuwp7BKDHaMai7DiMZt7If0DWCAXn2tTswW4wS+syUkbr9apbYWGxs6ffDV7n7Eiflk
fBm3v0eSYvHJ2Pgn882OuKUUPjS88MLH4cmX23MJIu9GTOFQ30si83NlGUhsFCNWdbY53x18r7mW
OsdOYRppwNPkVGU4KPBcZyXuAhaBg4ibXQWxZYhb0iVIpNtlKrAdgWBL0TiO02j5+yQMzEmoM0P7
lVkjCOZf2Ou14X38GVuCqWAAHADx+fitk5PT9r0mg/aCxUTDXErGzhsN2LUOBn4JqG4xUUuQA5k4
64btnYQ5CmygHzMHhUsmmx/SH0k0xES1S4MxxNhI3gZaWV6zLx1oFeDx/o6cJ09NK1gT3GUWewcT
TL3xtJMq/y5icorBNRh72pbxnkihsYFxBzRqvwBD3XZaQ6PXGFUdVXz/8qBR6MYgG95rzSVu6bKH
6EQ7oiUHcXxCRkC3vn2tlzQXHC3EY7twCvDKJWGiTYXX8QnK7lUPykN8Hs4U3tAloPkimPuGw5jH
t0GbP3GdXOJo3oZdg9M/dpJ2GSVGxnDOPHO144bBAwMEMqodnTOJYZbirP+ed0S7RNjsgow+OZQC
lDth3QvjNDtO/hoU15aKkdLlpuIhZVw+F881ZGqAoYt//8iNJm3IbyuQTbb2L40VR9EBXtmKcrn5
1EgY34/8iwlAm4HPtiDB49+O8+McgTRoIiACG+efPC7bYI6rNN2RUBRfy25CFtj7WafXHX0jv1dA
F4RIBu3XiHUxNm7b0wLf7qbFpGyR6Jxlj5RH0rbplDyNfaOu6tJumEcUofOQ1ReyGXpDVv+qSWgG
LnOq8DhCH844/mg8DLdGyZne1BJJUwaLhPD8yQEABuWBls/1c5D0LTHgJMPQN2TvdqIr05l0sHI7
a9Q5QqlsKSwuWyNgAv+X71+tEof6OekTIyfn7HKIlYsUxH3zrFHHOSFEp+3vDlIzNpl3Y/hvP6vm
9burv6eHOih+sP2Hmn+M1/LUbDqcQroHbVeJJ9VEP36T+rDdKKVKyA+SsC6n8VGAAV4K7u5sW30m
aoteNI9JHfRIR+Rfp7E5sEGRy6tVO1XY2tp+dA7XJ3zM35K6bcWaVdOFj5zl2qTOyrc041JxyVcF
9Xph/AxWrY2P2TR21ZxUzbjaDbVBLBnqQRu4nETVjJ7cQxJ/8+H1UYR5T+FZbZkfQ83tfmS4gUu1
E9HJ6dDMuk9FTE0Yrf2zfkSsTNqUaLkKpk3VCmZJNj6eY+LxmIBvrBsBT45s8vbWZbsBZq3e17wT
91xFFXkX+v6ynaNGFBBbju1qsjhGa23GX6ek0rPPA2Qbdfo3FTth/P4/E74WK+bA3Ga3yUZVLiqe
wRnRYk+OqK9J+l+P5HRYrxHE2rnhgIDYr5ZKeHBlaIbmkulwvJnjsRdzKBWDjBrYDexkbetw2J0u
1Bu2ls7SSA+JmMzP3MfwZL7rGHTvz2TnzxbdnXuVowmdy7R2u8ZqhtmCIoppZFq3qeeZLcxgE/ii
Y7hV2rAhFl+IO3NNoU8bWcDLyxWf3pk53fvgY0xCkw02Nt+Yc0Knf+pSaw2EIV0cLY9BBmd66u1S
g8254fEEj3XlHdPVTe33T8HCa8B3vARhF6HdqnvE5Vbah3ZlxoqZWty+nUAxUhdgQHD970+akS5U
ZPpFilw/exYuU5pA6dM3nT4KlJD8cKHDuEJlQbZs2W/LxbIZyfHwX6c4QM+UJUjSgP4mkg9nTQRH
SryDabIozJ09iaG6OydIyHT05tVH5FFXVS7Jvm4pJnPxDqaa7EvVUfmWcS/8chv0Q74PBwsyEWMx
DzW48DwMJsfQbkTuA8CCHj/Xo8KL4iq6IA0WBbkWIXVusJRHGYmZzX57SuSrWZQOcjiMxC7Sb2aG
3qKeiL3ysvNn9z4gmBFTSqNhFMoMUNNmadFyG/EZTmZXP17AyV33iIe1P9CIL/djM9PAMe5hEhXU
FISy0XcaW4dHc7i0UfDm7DwIhuj+RvZuM3MQjXn96u44MqSnq3qfFr0lVfUmHEy/WGsq0Tr7fMAl
n/Hj2JOuJ/W/Q20YtJc0y2AMFx/4T+QpOk4/KDRe9HpP2WLOcIIcDqi+eKv2lAs8OicuwAPZPjz6
uNbb/mOSg95T1bomzOrqkR60VN5RIOaDXQMR7bPzMeTu6VAs20EiVqnKVOLoC8HoTHiV7iZfInOi
Nyb3P1wjetRYswh+JSs/XhY9phKGXPnO03MP4VEXa3c/5qKkEHxMfPj+edTGoANMPlsU3qUpiPHs
Yb9bt/QThx7Q5HSD+SYkmxEjOlgpCQZby+EO8bPuXDIBGy093/LksZ0828JtdNQsy2biXS3vpHp1
L3YusvZyEbfb1v2fgPZBp1YgI6+Khn+gS34gh8PmcK5x5C6QkPk1u1m+fC/L3sJg8bRJfko2krE8
8XYpVy86niub14byDqCbzBGD88AyDD37P3QMPJtqR4tFQczsnXx3LwWUARoj9Y4LnToLlRur0Pp2
PI6Ba3UeaHV/STLedJDJldyvREg15CbY1q7+rP6ERkWfqqkUv6KiLG9G7I3uZi6Y8vBYin58eTRk
PEwq3etINlsYaqXUlrMstiNteWUrzumV+smOuth7nktFCk1w8XIOjOzf0VBESwIdJ0AjzxOHNUlt
ku0fMeEWG6BUCguJRHvImRYwf/9rmLItvZqjnG4B2yjYjlSXCwaf63s2rkDBRe2rIZILDgBEXvu+
Fm4s5ATKCq68kgiZs6HTk8xR9f2hz3aLvQtHQTsf8sfKs40LTgorsqhkVp2n1VLNu7f24J8awVZs
kBOxxo2d7/sks1alAjMyldCfJWvFeohwNV4K+5QeJxxQiDFupnQXv+Qc7B6KKDXODWW4P9MdOdYF
y22NPGIpq28qsCHCjk9tg6uuEjMGqoVykWM+BdciYzDlB6k/SMuN9HKX8J0Of49W5uVj1Wy74/cf
hNPgRiepRN8b3El+FYRoBb3TdFxnvtwhl97M3cJ8Z6MySfPPwTLNl6R7sGVsLGX4zY2Gv4rkFdx8
oc8qfn9viT13g5GfKHknJQ32nINxkxSo/4s/WDy/MJzQuMHQjw5feCzqQVnq4G+cNfTfPTLZXNct
Tf36SQumOaFnwPclsh3HwGKujD9FgF3Iw6oNItVWH/LWu60SjAXiXb0D/gIg9B/l/AvE1tKV0qcm
EtFaCpUcsehF4fEsssMRZiiIDvWsw88KUw3lK7W2q5ThLaagAnPKd0dEZL+f4le+QDVVG4o2QtG6
0Gvc9hZ32BW/TFiE5u3l3YSQKXc9RK1Y0c7/vn/Bc+z+PDKyyGKrdt+Fvi7+RxlF5D3rhyP7YWlz
zyigipjBQYwDgNJw0sZePMQ3RnIYe5Di1Nwdci9futlHjqvmD29ndHLUiibSoEGVylwjSW9XPFTX
A5ArALC91Ah12HPaIfEva6ltP4zwXKV24DCtaHPQo5CD3uOc0Yoy7czbtlSTu2ZcNHmcNZRLsLsq
elHFAHFOm3/NGYvszl7fNxeF5ELS3iYQ7B03la1UPYsQKqXFuKBFkVipqeunJgvMNm21acH8kEtH
URtGARsSw54k/rlQpkzpeebwgMIl9Bx9NuDIt503cjERMcOQT5BGn+HaEFKN/a9E1EDdgyEAz5sy
BDN584Q+LmhOw5bmVfyf0XCVlWx50t6M7N9YlNYywabAV2ICTNcvgEQaBVX/KVWSTy3ClM08/szI
YazfcDgM7M6pGp4Dzm3B/uQmMNBmWxsG6iTt8sc1ha4Dwt5BDSRpKl7kd7N1STPNAQFQRvB8bRZf
mgw4Gf0SGOlvQrPLg2kCEf4uz7WkUNkflSezL+n8XZ8V4XblZsCfyr2+/4H3XWPVc5KsyCMp7rr9
K5OiYHPPHh5eC6v3UitTKnwtc5sZ5Hv1ASLNSjoc45rS5HPLS2t6gacfOLZP41moynltWRp6OZVt
6cY/jJ9DhfjzdRMqb5H61sGfxnZC0h32euQdd10bXCb6REh2Z7fA+Sv9VJyHzVU48yDHxRV4ZkjQ
+dPzbnaZtgrNV7pEWyH6liEQQI5qC0N0i65yXftCZRPXA7HU+SMH9hhzlQU1EKHi0bHjy+24Hg3i
0V7xGlB6ujZ72vXoxkd+YdKEBkmS0Xr4kEgpyPockwjeguzkrn/SnTHth3UV0eiAzAPkTUEe4/fQ
qbLoGuVlAsbrHDFwZbcT9ygnFOAd+jQZCn3LLGuqmiOQ4eE1tXH6KZOA221LuEa85D2lV3xWVIye
Xpg1pBDQBUJRhT1Qec04yUkc6TCYrtXsU2NRXDuWv6zcK7yGNpS0Q8d3kiDfV61qJXJirkiZU9cy
GUQCcR6YSf3LUvYw9hShbhawjZpVCj2wPA6TXLRghM0REf9sToWb9nAZOz+pwvz9c6rWujJSR+pd
UM8SxbdAho4ADOxpYmM98z5MmDHuaHBUUOPrO2HdCDFbEAkxp7qB7fUCC0yKIyqLeyTDF/Unaq59
/Fi8FvWF+ymjpEtigEe/ZKZuw6t2z8prLpN7yASXPoJUjT+ButHCHuRL1BSoUI+dzTz4c+rcc7E+
iqjAp973zUy/UQN1phyowxDXyGFCErSSkvg56Oiz+5VPcOj9GsxfGjoIkRrphD8FnM+sL0GTyIkD
FJwYqPdXUJ5lzuVBVpIMHolPu/zHwdnfcYgyTqfQY3/Lb95T+P+FgUsqIJRepUqr1R/FkqzPnLs1
RAnhc85SGwGVvdkss14NG0Sj/4UgVGVmC1CApO2dlQ+JejeWqhU6kzmEzEXXGoU10vrp6KtWDkOM
oYPPQ5H9F3Ywl/C1hW13W8QpPG4ZPnKSQhRJXcMg0srSxpnyBMeySAoJ9GtsA0R1oVK6bWIj7v1P
mMxUaBQrzL2QhueQLk5CHUVdSMPARvK4doH2rV47KaXncdMFWDHtpbDlgiWoJkN1AvyBwf1Khbqi
JfJJ8ZcWDF1EEjcfgk69bdAa52/DzWEVgitZer2zun2kijIsz71xcjMK+r+GRIs9IboWQ1bUGx7Z
10kriObHSzZ+OjWx7wwOfCj4FpV0mtlY6TMcPPP809UEHa4GrYmBW1kt387q8TZfB+XQgPHm3h10
FSM1GOSyd2VOQQqH0tUwon0DiMBP/5794EZItoqO/zpfyErAsRp0ibtd9K+o+7D5HxN/BhhUXI4U
ieddFABqYU0EqLLvo2SZK/frBES/AOPnppsyzCyycShl/LOXOuK+jhbI+N+Y5m8Y4v8qWNkEKuqS
S3m+xmZM3jZ8r7CVideYYXZ+nQCovihniRbrmcbkRa7jYFvy+9Mxkl0C4g5QmQIRGYoJWOAd9x4r
HnHufbptLEmnx3qro9RDOh5zZoqaCHL9o8blSHskbWXaWYyhmWrcEKhKhhIQ9iENH9WASVeDR9/0
GRhYwEKFJPO9fu9NwAAm8GOnAUQEIVptwElHDJuk7jz9f3KAueaC5Da8+iC2wgdjNBwpFAbyL5XW
tJ8hL9Q0+UiT8r9J3mlue/oNptHYWv7a2jo5OJt2IBAgRjeQODS6WW1SEyZ7VVHiaj9mFP0yrT+D
5AfJUp3xHYBM9pbB8XcgAzDQuKJvL5jKGNd3y+Od1wqB273uQeGkPQuh264PYkBxI1KuDb3n8jAT
EtmR7UhEgh7xa9PVj1LTGw0OFjqlyJZ7dckN6o9f2T6+AW3+7S6ga8EewIiorMikf2GB7vvIx2eq
MeOfCxPtpanArpjNuzwuzCTYGRT1RLX+jECK1i5akh8IS82KPETNWZnm9sedqIhF9pVomVvHbB8f
zUDRoLDjDJoi28s6QFannFwJ4CS36SSt6D2mqrGo4go5erSDBSUWPqphInqCG8JWPQJLHAVgSCDW
2IBcGjQU6D5+4znHYehEHf/25IBMWh0Tx3TlsxpZv3T5j/WBOdQGhIGUXGtFKy1Q78arghY1eJ7z
sZLm/F55BhA5bXvsE08QGwwtg3n/JBo4PhpJSMOx2lMOFhHpq+38VWE0yx8xyrnzIgfl9Emgaq5P
gCwFHHMaoIHqA5wlrUrSTYzIz2EkIJtyk9Q6DvGABEUPq7enN7QJQPCGQ4+J1wIB1n2TZYR4NPcu
JCehvjYeRUavwmkucVOAfKMy+lZs0F/x8PxATynmJjRYnOmMODpvQLPKSpV5FXf09Uz55bbIlvMZ
pmwj/75ZSDUX2LlBK6vufXpG5ysmoPUfW4I5WaX+j1FmhbPa8P3BKiNWczMTtbKZjtv4Mn8siqvO
xWK0DV/A96jqKIXynYkN3kK/Q5JlGHNab7FTmoDN3kAqxeA57Nav0XNBZzpucbzyVg0YI6DZ/2b9
vYyggtO7/q3+tGEOKgjn1hLCzoDTpM+9FLbOt0SZgYU5lrO5ejhdFDNm2lmRLYmLhVFJ3q4276B8
ylPmPSDotLvQHVof/gyq9/z3Y+mMhQDIjKkCcOHVjH6kw3uXQvg6rTQfu1bnHatHMac/H/DpBhkB
jUELHFQnPd8b/am/y3HDOBucPzRbjgU/PJQeHeMTr+AIcpBOzrT4I7a8fG9GBwT9Is16hJD6q5DJ
GFb5+oBSha1XT3bbCsc+sllx4K/C7kIUpERuvzJyq6lXClBbMctZtzn3gGT3xZw4fSmx1IZj1rs8
mH7hZCA3kOG0uYZjZaCMmhxCBfcKjeHnrW4h1Mdtw0h6p/A+QLekIdmaMXYP7oG+jMXXGYnMriR0
MC9g5sPs6K94reX03XunRrxItQBJNk/nl00n7sFXFrbJWbjS4WUT2UIkOJWVte/SIimv+HQbn09Z
9XlCcfenCvAwM0IvjPig6PaXwDps7pteINFmJx+9e1QhlmxGzXsGW1PE+BmXcl7AAIavW3uWkA8z
WZuVv80YqwkqcDqJXNhtsCubF0gUozRn8ljUybTXHMhOfzm0ARarCclvZMUDDz9hc4jukG1Ptx3J
TVh7Zn3gNETRuBJEDFTCZWddnvZZNHR0tueAZIgKqUA4Ryd9Hc7HWRbrJ7gDsTKEysa08KSE1/KL
nMJIJ6tHY8BUXuTnd6b77GPF1mkTqwj49q0e5G954/zd+NMqxuX/nl2wzsPhutq+/n/mPqEJx0Bv
JY1uhRtxd+Ydya0XHUHb7kWDIsGuG8AwyRHe33zVg5Jf7NkVsr7GDYqY88JziCm6Q8eQ4RsPbFQt
xCJ6ewaCvUBy9UReIfyRki0nPDxxP0WNuplxp6ZXNDi8Ur+Ql9eUt6cwBYVs9YgxSijM2faJMXtD
ai6cvL+/XJ4/IvZB+bAOyAoHUADKMkxHX/ND6X9UPV9bqHt0O29EA0WkSwCPwBVSNEl2ULsQDUcl
/hClr0hV78L/Ok0z6TujfOuyqShh0TOT8jo+4upUv7CU8kg5AUst3Y6WAt0ssZxiU3LIb8DKfxsJ
WpA6YA2h7ZY8kH8p43bxOeGj4QyqiSUyTTDB2lWEiDL6kguq3+dCXf+jSh1FjTRXeugz4bJxkLYW
2AKdqaj9bnYJcLPtd8a4fbIr3qQQG8SuAFqluD79X4GISl9MnriM4hGCvB7MlnVncEkqsQrUi+SF
frVpm+d3dQEvfZy8s7P4qU1oWinuJPLuI/8vzk5wb9rdsh9GmGBI/DTM6909+Fv1IH2UNjpMGIBb
3c/pObpYITlhua8zk4Bgj+AwMQF7lj07IN+HDeFbXf6a6VcCxj0tmROYakesZ1tdj1LfHk64pLzB
4nxIQwifdpwsHHIUipaHegaQblt7lFU6J+6z0CqSNOi/be1MAe8AyczsnQIZCFB29qnuAlCLt55s
QPVj694SzFnYS92FoC/QrDNu0mlO8HK89z4hm0hPiQVA11gP/MPpxmF/H7nmzq+LUFEJyNSjqvBp
RwLS5bJOPlNBMNQYi2C1KMAg7YKjYQXbTJ6hp0GI1jooXQCrCzR8/MCCGze45x1myCl10FOhGhbd
4+xSv1xOJUyjJPftz01coqKO7U70IGoCwmW8Nj3pjPOF00KTQF7VL1Jd/qqsc5hNrBe9dfgeaAGe
ay6U8TG/HmZzrozRyyNz/Dw7piwJ0a0bqBzwftUd0Awt7n9Sg8SVba3OZQmG8bhjoM824Ghq7qzO
yFs1BQVX5Q+w1HXS2HPslhwW71pJpVW7X1CRebV4c7jqL+D65kpVsLSIT+Z3MM1VKcyyXZZujhOH
g7JDZKMJxY2uaPsqngbRtejSHNUIuryqg9lDYrQxDQ51zoG4P65l1OOc4BY/d50+x8W+Eu01w+p2
sYRvimTfs89ALrocHq0MIWLsox4ftwxLNud1jBIeJ4YnuOID+LZY6iCNJ3cEgWSdcM5GKA/qOjJ1
D1Cb1msGVr3M9OG2d6P4BFeYsQjw4kzuNl1fuoDRAAQfciDN5YAwm8Rm72//RL8jbABt0oAx05gT
uv9E4ikMm1D8sshkOrNbSnsPz+65PyX6xf0i+tIp9+MZEe5qeafWDF/o8AICZyYHoOBPF91AvObc
RhROxf44VNVNjl/+SypiGicZLHU/kdwp3p5b/NfGzUgt2KmiHRjBkaPodf8K3yy13T/Y2PzIC7kw
yp/zpdl65vNqajvzJzUCIGa/98wy0iCddURsyoenYq8TaHsP1E1Q0GB1037fr5qD9WKdrhRJ4Ffg
d8H7Po+sRf8YuFrAkc/fBexT1RfFquiDumOQL7oUWsNF/r3xJ0NbSy+NHnUwe2rutfvoHSKB0iSa
1LpsFSm/bVkFBORWnVewow3Oq9oZGKoUdtWAAUlc2LBN0wM5bwTalJu8LLNG9YRQmdJwVYPGvZ7R
JeiNjFK8fsQGUbA9XUvNpTpnuP4qZfB4r1BAnsNmZxpTdh/njrB8e1SqsdxcqtfAOzDzNZxUonFp
P/p4EeAAwl/nox+Eishcz1FTiyH3C+0BrYksqyPFRvWf9OB3Fc6BRJWYsfNUeLEmeRoHpCIzBHZZ
ZnIfiVPvVAUpWoA+UoHHnntiYvvwjEYYDorXcyDFNmHPtX3tRaKlaZZ9iykCNtMUBmQn/7Ia4TB4
HO4rXHFN5X6QadQvrT4hpe19qChwAbQrvlHc//i/HOf3pcPhHvoCpOQ2K/xhgdHIYEzW79dWz9OZ
Ei4lV/PQzZJVAUqQpFh4Daki/xs2hTmHJmS5OwdwwzEegFx+WM3YHVGcLqo+PkqM9THubpUUy0dT
e72zS0lR2RAzWy14Q+2ngW+G+xILl9f7nL/WnnchjNLC8Zb8CyA6mTCee8oEAuFGYu/epVWq1OR9
MtqxSBq+0RPPk8BnFo9CS5leQYiwPOIoKJtyYhSDZ5ab1BDNiJa4cHqGg8q6+FBfUzWb6/aUOe8T
mYcQzhtwwnlc+vBroURimqdqkhmqPgdUmnCUFGvLrar1Yzs4zMlJ6JVip4aDIp0ZN36d2pgBHC45
KVMy70lwdpz/3YEFMixHqa1ggw28fhP41ncP6e35CIFSS55xBTvRecu/MXukrteh+CSVUWydpbVQ
r3QK2YKbP9DqLXjqWrbkEsq47DiRKeqhCl+kJYRvZ7jjxJ8dxfNyNEPtKufHkQYFLfx5VGOTkJ2w
gDFJXZ2Y05UMn6GEvXiFpxGgFl1i17Xs/p9SgAJN8Lj6k8z/1/mBiGPekBtPSyfSmU19OzPACuwG
BrSU6frnmWJNX7PsmAFJOhvD3gKaHENRQ6jdWztAd5ODHx+ShuMKv1WUgizDbRSifcANcCnCtzeN
oPIdSC3kmU80StYynGhrbhYONUXWh5MzMfwWDcP4SOupeLpqJBNqMPvLyU+HLA0k4uvqLR2kgKyz
17UxgxSY9itP7LX3s868kPXrO3SMAKUoHodGTZGjhNeqZV8Bj7iTK+g0dwpbzMiFT0OnEyw7JiG/
o2AZWNserWm9rVIVVxHjfypc5tiX7UYqqigPc+xLwfQ1feURu6pyuw2wHJRJl6VupsBLmCFAREkU
CLimvzwnb9eFBs14lgA6XJKTVOILw+N+nCAdepFtcAmnmmK8rVsdL+slXaayJ0IBCXrXeVjGQwgd
/HCtC9zxYXy1krstS9wkqFxjPKkZBR7UlyJnvwubYjzKy4go+i8gC9Q5A+I8vV0zttvOYnj2Otgp
2dowhUDahYoCg0yz8W847diJ7eYbcqNobAiLcyXOp5LMWFfpJXmNXcELRlPE0mNs/Z09yQuPxPT4
2MN/j4GjmLPgkK+EAnyKCRePtKsK1A4+vhT3uzJUvGyIgMUIgeO1zYBbVH5S8M1iqfVWVhEh1//a
82Z7eQbBjMATTdz2Uv7DNB9eyYvtJrcUeJqcbydK34WpXXr5anfJQsSdwXxysoxRnC5XBajTqIEI
eJL1kGQsmQFgN0p51qsIfxyGXJ7945BCZnWNJgDKfL4XWaIULBdre0BjJld0U1mVjfWxGb5QjBcV
sq/5814hYd4ucjGYbfFKjgADmhGEdde2oMGKJ6T/tarwKU3jtWvBtfIh4/iHECxCwao3o780zd2N
L1d9mfIMzs2AbTPI0si4LqO+JSUajWtI66r3y1+7xL+vc8LSvLjsoANmR51Ge+aToNhVPlf1KAzH
cJIDo25A/ru318xj3wkIwJdvkR3324sG/JUOILGS0nmUM7dk9MXWWwMg6ScrThWD6sEu+w8Xye9X
KTCvGhNSr1Uo6ABiMMGIU1lSE3cVq1VJ6MxeHky891/B0Biz2s4sNWFNAnChN+zESADlSKTD6Cr6
H/UUqQRdFtBQWHXg69oyKG80Y8lrsYD0iu6OWMEcFcDRnBYvRoUUwUZ3/8MYgxpessMcnZe0Oo1A
yYCqpZ3ZK/sCKLK1hmwwkq0n+MUyrgNibdasXD5XHLIShYYFV9hnUorcbzeNarNRRD79+vdYc83s
XmLCDuq2NgHATpwIjrjf5bR71p6pzD1/Sg6oXBkGnnm8KI0qouCkrF3hgd2DZpNWcwdCc/vzZ4UB
tVqCkRiTXzcUVtd60FAaDOWCJeZOGo4TBZn8fShj6b6rv6Aj8TaqullRJlnN+iAFlWcN80WowjxF
ZP868sLSsnwGU3PX0WWiPMbPW3yZ/em4deroOp0eQvXtm7RmBfIA6zNVHYESkSsDDfwbdrNxK0Oq
WkOUwsGdV8gQD6WU+6PezPSLWY+r5l8Jg1TS/+rGBOMfJKOQwvyycsZldSXkYg4844+qUj9WLoGr
2UO/JGURmsA5Erb4OiMK3yV+HBfqoDLPWZTE3ls2PdiwwkK3T6XoTKB4EuocWO5PuKQgOk23HOCy
y0uGYMkyHYRpOvdZCgdF94tIMBD/WlDO/M+q0m3jvAwKdoYL4ZQbPvylxQMMSWOlrtlK3sVKMwT5
yWDcVqkANspGEVo4Ju80GroX1eJLQCRgt5OHfFQktfHY2Tgfz04jrRQqyYydjd1bQPD8YyGKvSMR
ou1V1+VFlCfZ9IZfA5sw/BNkta6W1IaASPweVt9nqv/yg2mYBrUXAXdbCUwX40MB+cAcvksS2+Xo
d6hl9PNrnboAIPMuaa5bb6iT3Xtms1nfUT+2emI2t8rlyS4HQDxLY/MEDxunaRRxtWWaYiGcuCIk
YNvBDdSUcbb1KNfLjwXwrr9uk9HHoNU0NosrLyxNJCOwqt4UTcF0sVO7Mteoerus2FTE+KBXQQX9
B6ofinVUCUDyISYisRigfOX1sKRetOW6FicbqnmawQ8RnVR0bZfUfJlyvz3st9f5a8/X45YjaTRc
rRkPSmotjirYMmGEJ+XV59xZ3PxMKWel3UsVro0NtN1dZ+zHWnx/BdxA36/4YlT3lXwYGUam2WET
LzibgL7PBQtT9AgWKKR2kSoIJyWB6G1PBYvDAq7vD6hBNf0wTnJjtAoHtrfj200xdx+WzEpXs/Z1
DoDIyUI127NBbV2+LTA0qnzSqEp5ZhtS4BDwvUOMBO9iL3K64/NRLUhrQ7ijUZdo/KmJ+6bDkrA1
8o1R9fkwAKLzahLTtEvlBYA5m0qkNyDzwu8TBQ8uZsLyhChwX/h5Qts1uS/cPsDO5LMXYOke3qFe
W/Zk82pKMkmEOS/cLQsDiLsUrR6mT4FhSghm5HnmdnTsnsnia1GkwJZ2L8ZsipiOkyn/clmEieAI
MaJDgQzbQWoaFVZDPfQ/gvXlDbbOlBk9FJJT8K7rHhCV2uXUnnLcO0IdzDKa8rfOTVF2oSuf6/Jp
VRpdWtW962WB6y+1cMCXXfp/DsGw++DVg0P6xWwJMZnclLlMeqWYSoEXq6V1nWKnXfY1Khu0Z//P
k6OuY9z2GN4QFQsbu7vnkL2PkkbzPcucwtcFimVZfQoxa9ZjPFP9fbflTMiMYqRN5LJO1r+yWA3w
5kBpc7M0d6fSsWojjOkgQ6S43c9Xz9MObYEcCQGX7Nb38kh22LWghLIEdZHaPe6aaL2aRxf4ChMy
xEqwjXIZS47W9kZeRLJYp3bZO3Pz75PLN8OlpPM6LztyfKq3dUc87Dq7L0gAM/GslyCyHrwLtvoy
qWcHj51Qen8jKoHvHn302HvMfqCy6/87Y3kIEmL047sqBuSYO6JHNSo/64sGZeCKtmvHsy05Pv/N
VBPFjzcCsDraA/1hk4J/Ug12tsJwFRKCLOBB28kp9jefAQ7gDm9nRGvejsq2L9PwS5VAtSijUXej
tnVr+x2DapQDOJ9HK9oWFvS5U0TZhrzf1zmac5oynGfP8O8x4bbtJ/uO3eqZAHvwCjhRJrgWPNUK
pJ4AbB16PixP34z6R7nV2A206JAwf3rvH67wHoG94i6SHV27EzOm2C1niBRgBVnCdHY8geteBUEW
4HpxYCtJwLRYMlbKPT7wqCIwRK+20QAXfWBbo9L6cVN+ftVCL+ugaXLEeJe5cr0TT7jAe5PMm5Zh
KhK842te1MZWlkncx45mtazjQuYWUgveVbkrEaDWluWl/995e+nw3qsfHirBhgKYUuvQSx2w+uO+
2GnB5ByDNlW1ykzd5BOg0mcQ807PAjbZ9t2Ab5SHHN3BPTLetFUn1P1NxtTAvx320fMEQmkGP9N8
z96gEvE+LibFWhtgkQxEzTON+zGwq7DcEW2QJzIjx6R3rAUEsF4BcT3x0CMbBusNlB0UZ5MtKE/W
cCsdGrXr+2KVnkjoIWwANMdNzSTtshIDYZHAk6v11F3iN+80AvlgJH1OPQrJIQX6Tg4Zj8ahe8uW
JHpnq8qKg7Wuilerxv9ZFOp2yF0fmo8z+lAO9QgHbenI/pHbAqRd7FkiGmbMbn4Jwv12HKGn3963
P5/xpoN5shIYzdYlboWnKbS162inUy+oZAUgR3otk23sUQoAvi/SVj/F30iAnx0dcjnrpuRrKFKs
rKQogQl8plLKV4EoxcMJLfbcJCyOTaZtn3KKC1SBiWuLGwMugLTWiXLZFXF38g4LReYbUdZrk5Vd
epU+rO7qZoA5bb5NP1KtCbR7O0I5zTz1nTDRSXHRNYiNQLdEn5IJTOyJ2d6DnuX1UcyyLX9uFwSg
EtIOfIgWG3cUlcnSLBtHVaTOcx92DoKgoHk8KpCEwmlb7tUW6QOIR93HljSIEY9PYMqU2o8xrO2D
sFGSBmPMY5Z4S777NuABHhphHxISPbq4+J3d55FIQ2fVwV2eau06NZ0RB8GjhU8QhnZ7DBxFNgf7
Hyych6n1mtARfOIZ3YBQBh/3VLWzjX9XNILW1ZBX09IzHTEJi0Q4cZCeVV1u7kDa8dlP6+4KSjqJ
1256n6KZmaoyE6saRcAC+DNhexXoX047I3fXKT9I2RKhXiOPokIUD4JZB/Fj6QnanUJN5dfGNkoS
n4EadQ6KU8vDWeMZ6rEAmlD/aqHSfzt8L2xCL+0G4cUrVLmjl60Qf4tzCqQjyOLPnJQeEwhxMZ4i
gifOE0d4iLet1QFtj4YrvF2+w+UY3GIbD3+IFN9gxcBoddufvLoPiawv1WHXycRqDz0rhO/kxE3h
UdR1h5C2NjbtEuIjMFD79a+lvsgLYdrB1XIFfFiq2BPrs6K78HNL0bTez+MFJJrRf5BZ5M69u7G7
aw1DOfK32hNKQWeNUkQDzYQHt0Jo5n91K/nazabhws+dKAPJtb46I2rUQ/VUYqtEnZ23+zxsinG0
W1e6X9JZjmTNG/+VZ5hRkhSX3lipfV2fJ3kNVQEAMzeHPD7w55ERZn+DrkTu1OBImw3zaxF/jvxm
GOOuVri/UI75YLU8Z6HjEpwT4cOcaCS2FLwgE5+KeUvodLMKxgHmeOdYQx6nii5cUIaaFHgyY8H0
c5dSfCVKfkTSTFOwKtgxWzUZLoAHAwlFSjaPEgsIUOrvcOxb+WZKAFfshcXR24hwVuC3w2cr0qHb
4oGYfEL2MZzU4a7xiEefmalqK6SL4Z+/8pJWtI9JutcgRG3qAZCMwo/77DqdlwJdi8A8zPZtmi8l
VmgWwBLwk4UJ4bLVsSinzyX1Kpe/qZ9SHtGGB9HFh4LUdLZQHsjWTbbc5OvxviLCSAxlJX1afAbf
T+LUmFdskr1Idv+/jTpu653o7KU/TNbP5NwE4i7F15Z9gsoGdK4JXtfdr1jTowCVEvmmrXvNtEz5
YcmgGjCrd/jhWM2u51E+KXIY7DNMef12smJF98H98tMRSOt+KGNOdZ/SUsmwobM+txy9HyydlyAL
jafpdWMthF0sJOz0wf/2khQli5FnZGSB3ztDf+06bgmB7q6iPP/aeYjpe515s+hBQDIjEXQuqBMK
zXE5Mc8pW+QHvO+Q69set6+vjgsW8P9xao7SwHkr8Rt7ZKWITi4tCvn+8Uqg0otXUjHrTdMvXTO8
8YN8hEOZS5Kb2ev5MEJuZsjZwTv3GTfnRRq4h0FBMqPBmf6nClbWweJ3Izig58nRZ04SSaqz+qKK
lyeyzDwIinOuf6C4x/R6CjAu7V5iM2LY7Go55fasTMpPH9L/V0Lu8PFd+aK+L04zYXFDPRkz4ngp
SKgZyMTo1TPkVq4Cje/xJK0oyk0vL27YAQ4hboHTTXFG0mzW/aI2HNbLq2dajYa1iF8dFhBZgoHu
r3EgWi73oMwwq3WPqXJgBoMZqEvCPw7DM88qkov8OT8SKtATn9a15zRDaCzzNqfTEwmj6wMb4I/1
caEquhxJ8KLGJf9lbxcHPv9+m7JGv/aT3iMxoD/gBNB5EbZwBQmwI5RYfcB21hVC6N06aK6CH2si
W9MXhgSm1l9UOXkEDVdeUTqp/vOyf+QaLexKDnW9nGQF9rDCgh2adQDLV0nxwfkkzYyaZZ1qyx44
6DfedEB6uxGXKNeUlR9OCGp4vTiqrvO6tHtJNYdTj8j/7z/exebBDDcb/zg4Er4XL4uFUMgyhDdV
0LjhLemdORjRmm+n25Lrjt1JEHl3noZPNoR4BhJ/oIrYMbVoCp0pWHhxI0yVCLRzrVwOTvXYJAzC
sn7k1GFZuFv2hVv2SOjaJ9kWbIOsuRYPO2AcL78vi1liGtzIdKSUZsCLOTfhHq4nDZXTQ6vrJVXG
g5yCCoEBjO/Lct3BbpvUXiL8fCuGhXtDn3O79FC29GKWHqkEkNjNp5d1c+5kJUOAD33zc/Q5j7WO
aLvD4+nsfHIyMHYtBE/gw1IKp3PR4M4B9uz2RLVELcaelSbynakbfpeysbVfhW2RQwdeyIk3Yxaw
4yLdLlpjhKDJxIn6H6vFKTPwzPyICZNItyAGY4XuWDNcjQGhXyre4gCsvIGLWMl7wLKBJV6yMVNw
TUUEXuBcjXmps/hHBke7ZFkn+dd+8bOPtAvcTSYGlrFSY1naVGg3HfzYhmwkeuCH3MoUFdoevFZB
toQvGEmPohAi6U/w5EtolaXGeiLZqEZF48sQwt5REFnhacYyKI43TB4O8w6HhM/PoEx7YI13UQ4O
WXcYw8VGMA8wSAOG5sFhxd4rMsmsfNdW35T3grd2MKi2syPxc9SUy7t2rdTnuqnEvhtMD8HZ+82h
oW4IzZstFRnYMBHxwI+UINHN4KzOfStQH4ZtklEs0jv8Slx7ssRdzFPujJlM2cXoIf9PhqhLiZ8b
dWdqHc1HoMlPRbpE6YTnuSuKoDY5/uNtg0GYMokMK+uumndA3OLcaMUMVzF0tLO1uZpWONAR9Iri
4RKzCrcdHv8/nf1zG+Cp6stlJ9IhIK91pPtoFshb1KYnxyn9djCM50b89HqPpS77BfllC/v5BhtF
A63HuGsQUokuw9yLs6UXvQ8fkZvH7dXQZgzjz29+L2ZPNNw5Ru1VxxTovTJfAjNefQhfPCRljH9l
XAueVOnzPmpakV29S0/GwpYjrXTwW8C8GH5Y2jA/Qs0+Hk2GJqhivcnmyRxYPQQJ9GpEEkig6EfR
AdQJh0b5SlAUaZYYOW05jeEjBvtPoI6a8ahTBux5DuTTtmQF9fChQIzl+n3gVvbgXUISz4S3BU+f
VR2XGXg1daZc0z3lS+hMoPx60B5E+6m0zpJeRQG91M7JiuwpmTw2aNwdKlS6IX80FlIqICZjJMv6
wjT49yqjS1IHaKGJ9avPnfdJNZ3EwaGQsRs0zScCaKmAAsmhJXY06fPuVk4iDaOHWhZqCC9FQY2v
Ws11VpDs5zjtfeMvukW08nQag6bL5aLU7cMTgzk8//tqvcbGySZdax0YK4kGjtCrj+JN2haTArZd
WmA9is+3zJyWwvW9F19/iloM+XA6c5erG3Ts0OMZJ/kJwGtSOyz/wuSh/9zxW6sXFInE8xzC3O39
n+USKHNVHKSCMg1BkpMhXvYY94X5pHR1jJ4/YqWrkLsNQPu2BvYJBvHW76XiUY1gYsUUViZ1mjCT
Sn09+voPu8sDBJRbzFS4G5eOMAph2EGeK81jBGg0yUIzyQrrhPCoEXmNRb0F+ZLrB0IduOVZ6cGF
1STVnAtSNpjqCy3+//GUCYzTXQ5LvDNhswT/4KHvheYF3CXk+KSRATbClF+UumbtLs6IYy4ZSIhW
jplG7Wm5ZMfs+GstQIdBOXQq3ADIlI4euI9S+6sLwTAx0LJTs2kHBWuNx+sET/jZcTHg1R8jDtTE
S9vfh2zT3P9/+aUY8N5xuGSBL/4ukGOBTZM9ggvG6Yi+eD0RJxfpefFNRKt7AR23RmjGtaSFgxvD
qxrWP7Rb2EcJzaQEbpGUDoDwUF/uftwtfA0JnnYr1fAn1Pajjzs3shw9d9dIfdkNL2gcLZzbYl6Z
GcSqpehKh/tUymQPzi9U3s+z/A3ZkAsXv1FJ8KL+firLN/vtYEM0/MxhUIaKsMnn7LdmNyCUPwlL
3nJmw8AHJXP8Jcjai+PveenblzL0hZf33aU9c7vBuJaq6Pk4PYqXFsvHU03wMJoS3QxUVVNyV0Nr
SkWXxMQGd8xszWhmvCnuB1qqGXDkWyuXbt8lJ/REpuX3CeXuQGGSjT/PQSrAHg4jsdZJCEo7xrif
tXP7nILULfg5AwjxdVSJBdSXwMyMCfMEMYtVbGISXycty07Y7TC0W2USgMxnRZdRuTovmoeWCh3u
18kH6YepjMjVLwCK87AWUn+qzVhhUKkfFwyK2TEoOKQOek3Hc+Ud+yhNXbtbJW2GaO2yTJQOLBBY
yu1q7nl4D0HYeMXnBcXzp543AyAGK6MybctAcqJoL5JDrlX9+b0xNdAIz885+VSYlM936pzBJrbB
4lwtzPS27hqdxZuiyoINC+M/b0ziSM9KIG14s6XYb1LkfVp1xodJaBHtUireOLxc5rAwfWd6fEd8
+ln8/xsEKTMchKCZ86a2kfQ8XDHcIpzQKfvUoBL2bcFlFtYTMMPMgaE07GUjxw1276eIpsjygmJx
FOBphMHqHuJh3oW9cOTK/DlSg3axuKRK6M6VTXPWoEHosIus14X78natqiC4aP7pNcaIuQbfHVsD
pMwWhBuorwm2B/oi9kNOHWilpR56a3udCO2mv2aUkP+K9sAVta09fAILKboEP+DI88SLNyBSrgUB
Z4xl4sL53KvdfHgOnjNsDgvZ45CEYi0VJ8JriW2rOKgvuOAi00o9Scj0GdMi35gmpiVcmwV0fDpG
NTXk8vifRwiHoX5WYqhF4helkPH/x06Ya9JrIbWYho1k2paTRGqbCDjSbb8rwYgy1xQCUHV39kia
pXL8iTIc1Zwam0AnE2wIrqhOz79ATTvoryA2QN+gE2pOEyu62DhIgV5n760+T0FfpfdQ72INI/hs
fUb26zeEGe8xuOmIhE7ICOyzEnmmXeXKp0EhmXK8kbutiYR0lk9e5iJypAkimg0LncNdkW6IOHld
yv2w++5WnCkN/wdiDWBaui0D+BrESZZWA8q4W8hcDEGKKLV5mQCpfQlc84HW0aXfUx02m5MzcBsI
oIPI7vPjwiKQFhIOCon5O+Q4fVTzgUs2SSo54OQN+6H6ac/HYdqvLFmBnTDiA2QtbEJIczAWDxP/
uuVRzUrB++65J/p0bj6fvNBlQ/uNYHKYQiV9/3Mc5AOUVdLVEKFHrzb0ToQKkfvc+KLTnvFFgdC+
JYDvNUBsucC9dlWlLwCfGinB/KUCz5B13Jn2xSwrkSmZu4kxCu34WNKVz6O3/NZ8mdfAXxSZvv4f
WKrOBoWCzUSRxQ47CZh7vj6qHjeNWiHJgiwAwzttYycu4LJKvqE7HvS31CteKqZhtkCjXQfNI/Ks
5wc7fIVWPhwfJ0miUx6X76Xy1Annc2mZlElgcwi0Vzmd8c69qEDls45xD1b/NIQU62Gzv1kKSd2K
b50SPKbceJZOWtnrtbRlLTtpdj/qMW0lEbsc5/Vkm0i6QhGH0Y4kye9Masl+d3bHyVL2K/eFo60g
Koksek4ck/wHPURp/iAwJ1F4IVg94Gm7Ha7/++uDiJmbGwvCMlfJcLIvzlOiUcMflpEkRfDMiZiT
7Jw4Erg+ziME4RPVB9KN8kWSskTSTxrdDC2y3udT5ojfnw3avKYpAoNJPPHTrG3brkrnaKAM67x/
jgMe2thRcN2k1TbCOICxPiPdEDXmsXxjhbNlDLpAvpGVl+LB3kXJpfewCCKVi2PfHQ1+87cyrHgY
xBo3MoLleiEjE0l7oqK+6HGC94Y9qnmt/sgSkvlpHYUhnH81Hf4eQAWPF5IMziMrkKO+MBeZLZEd
cp2tPkyPsx07zp4EYx/BbB/MsnvYobDFazj7gBNl2hdnVdhUQM+t7BtP5rJDEYzecXvFOAZxtGwA
gWge2TUTLKf+EjBmhiCyU1LCqa73rVCdjMqEwM0d6waWmiOkamXUXLYwlw6eWcK+nmaJtvvq9Rn7
4r0aGFDT8ePLJMQz69Mid5tZacgTwHms/Cqsh0V766JtyK5EWBJTHcpEZu/cZhlBL1OFmakYmYoe
67/JITeAMjN0DZ0cvtqkrkRnF0cWguaZt8DgOCaNzpA2QLvjXqqbkJxR0pQA21UlcP8a8zWUp6HX
CQBpBHzShs4EPyiEnBPcNXJ7ZY3AXDe9yBaor5ewyELudzNoj/PWgHcVTi9mBbo1+a2zY4vXMru+
Gw111GjDu/B9x9hZZsoPvRPWyDqX/Xvsr6PnR8eGinUI01bcAesGZIQTdQlMBwmmHLTHaT8AKq9A
cAr4iLeG8vjYhAYvcs9WrBYu6uGcOKMP35yELqt/gusWejc6pYPZBWrTu++KjhXGZParpMY1SfoL
4435r84aM5EAadiTWDQyqNuMabEAepACj0iFUjiegyHGU6MH8cbwrDlU3zASG3fkGDgWmZV4qPny
Nr/vZPe9x4d+n9H3Mbp56MHeAhHhv8UyrDU7aqvH3BlR70bGa4VtvdWdtYciKszvj0jAOtksQwvY
fnl7gMDMUsMnYJrEKWnRV8BeBskDzj9VMD4EfYWh2AXhK7C0wYEOBCdQifFGOq9qcuGKo+tDQcat
ax516d7U3Fi6bt5Qr/CoZyEzIJ4wcjSvq8HwngHY2ziYBNwbqJuGMDVa4YdduITfRmrSm3v+i1WM
rpNh05JrB7imwXxhnhrg1c+cMZIuVlPWyuNZNMz96vfU6irmc8If3YDTNF8NxyJaneRSquCLLYgG
BW9G3SYLXM/neWF3vp/mONXhLG1hxnqxKbNoT2jbibV1+773X/gVCyUfJRdavh39pVqfoR7CsFLn
LaZPTv1qC7FlN+PKfHcmde6OS2NNzpryovqLAXqMeSn9p9bBN3jej9Fy+rwo+qnYb5szwFaIwM5j
5RXGRw0lLSjZb4X1U7vFPkTH8zuOkVT6HBq4A3JQ1zVM4QWWftwQ+V5hp+zYl1FeXrE1JasLPvXn
LoYjdsOGmhgE+UYWWeOTz49JE4ZdhISi7TgYZOv6vjGeWRf52B9Uim67/MmuisusmW0u28pPQKtx
/udekNGXUywzDS0vGofpikXRU61p75GxIYMI73IlFErSnUrxnT8Cum9wadYfH67qCwJU0uTIDrwl
URnEkPF7KZAe4vVv2mlwIuVBVpqY0EmXYjj/3j8dJWEVPLoFsjBWQrk98iMQz5s+yT3uKn1eH9Dn
v1awWBMf2UYGbgTIHuggcYpXcUVnzvrzKgigJFiPKGiIJQYopuVKKocofuwZ2HC/vbmijJ674/de
6YOMq0pChCxWPxdthk17x+07BUa7sEWEyMo5gTszb8daR0v8SWK5EEsKOWmtasRatzhbHNO4feZg
VTpF90KNq0kKMmbhnW4+VzD3hJAjwVqIiVUWx0E6w9K5P+CBaEWp+Hwdy1gToWxFtcbCRYdyOFBu
QTZpn5rklUJTPEjGQpXvTEvOjSXIL0U+TW2XMshrrunqQFEDQ/01Pqy9h6dRwSXwRH/FXOvmBlRf
U8nHRyB514XZSOjoH30vmkmkv1fTAHyJMgFvYQVoOjnMBnAvKTdGf6F8YHrXOQWIj+ZkNDsD+ILs
DBzUyhbUCyuYLnICxjVYMdmy3xEW1zvcDx9NvP9VKYST491E9vErdzcWgOby2reImxEWUQH34eBZ
YL9qDXG2NMhiMXyEWzqhKbuuiVcEcNkQFTrPfIwVCAPyhL58ogELsCeXdWk3ZF1/BavoaZhLj0BZ
Ztxjx7LpKretEJocJttMax1+ZOW867GG1Af5IRvqicPsnqy7qUbBcTXgY6xiLm/oj/7Bf7AhtWMG
zMTIMJQ4kkLR6xEpU4VmWRGmURVhoYkHCG/as+ZOzhUfHROwaXgbm/7U4le2xpQDCIHOA8IqTe3W
kZ2HBOb3tilwC8/kEzKNbY+n6+j7n28XdDYf2m3H1J2f56F6Trws1kQwVBjFs30/XPiQpV7bveXI
4pS5j/tdOK4L7MkeqgogtPQ9Jp/iEKcvwZrHse2EoZG/hY7SSM47M8fjkIwRVfcVfkpMqGsJcYX1
5KebZorMv+gDEPk7TjHh0gyCB6jsfOi98n/j6TI939ceqt1tYROvseq0DhgZCsDgF/wULmvkcoCc
FGvUJL3Vt/UQxPBjZsB/0fM7TMpGro9x87jkFBJ+IhMKJfcHTnEJGiA5YaBplhk4/CipljG+viav
V6Ozq6QubKdtq1LVYbh2HH1qOQwIECHiifzIaIy0Tx5+QFYFa3gNWKMjgys34+in1vG8OLkRjzf4
IELCg1E20cm8WPSj1FXStTp1y8aOFQYFw4K8QZS/RPsp5qVCcYGmyQ7Xp9uDVYwKrE77z5klF6ed
VWNB3iZFuM2NBMyimC+ZAfY4QlPlizAcx/4WsDgksJZ45W14cYDT/D3dEiKTODZSpmOuRNLBRP98
Vq4rX9Wl/EOft25Fvbg77fhu/OlrxWVGvEMALun0g7tK4KFfh/vMdkgU2DrCC06QcKT9RowR1wA6
2XzIihbFttHSvz4UTaf+mAF/XJSvCKlQT++ENpnVMHVGIp6dbITwSkUMN9VcOZEkeXFIhnTbAnFf
Fx+3fbmn5XYOtEMec6zKp9dweOLDC0t1c29B4cQnNmKHJ5VPx757CIaC09mHQXroAtbYv/voEegk
F+gEP86EsjhXQ9o7VetTxqA0jeoX2VxigjoGlAS+bXSvFkn8ujC8D/vbBFegjI7C0EHIfhlpUtRH
fd78Ec5nOARg9hB58PV3O/d/Ft/WiHlure04oDRpbaisbCZBYUsoGjXf0YldtfE44DnHpV3ZIaCc
oj9iH6s6cSzMsOOeFl0UUcIxs0Jmm1e+7RYvpjPAojuMfTw6SlZovWKY2wobkKMFu0eGdv4J0f4Y
XsyR32Zdwea1eV/UBdwEyunEwoBit8VYNXJzCax6tuFginsOZRhZ78FcU/54hIzRimt7W0SHPvH1
8lV2uEw8OFHpY8NXRz0TCbfYhhN7YlKUG5SqQx+xTBkNCjW8pH9zIi0JP7fuAUqgu9SUScQHZFax
MdKp5WChKKY9957OKlIas+QLmLe3ajOrcV6lzO4M64G2XH68I6j6QlcEr855sP1TOTLMWgCxjIyS
JJ393n4fJuVyZz0N7gFl+umeOUML/yzmJPZ13Da+6xN67s0Srw1y6B5r0t/4vQ3DJc3FY1Gqc8wD
LCdI4bSAYc3rNUCJxHU03FKQm8ZXc9DgVLekDOI+fF4T53Kd0BBtIAiUwJEQEUP6A6XnzsOiwD+w
33tExRRCiFUiOXy+8A7ofij7kf2YynBaFFgyGERYDn7Iy1aii/LWn7bmj/TVDQyu3RXVvzAthALS
0vyF0gPeb56fvOLp1U3OmnVq6+MTO5FY5dFcQwWQFEBMtLB12HEh7FPD2ZQCpppAG1NMw0bv3aqs
Va6ZWjlNEKyut+cUQq/0O4h181kd/kBCdqG7r5oUWIoiJXRKxSdaWT34bK96ZjeCv5THcDYC1xM1
/pSAncylHtN5qmBratp+L6UrNV/PRYJ61L/vAMyZBCqbImsOaVZRyzjF/tWIVEf3U+F1mWWEyj66
eKtgBHq5DJPpHy2ln73JGDhCZsXrDoSvG/WaMc3k+bnLj0hJn/02bZ8G239Nm/UQQyLhQS5GhHJh
87sC/JIvxV7GwCiac1+h0lVh52dgfwM30hPwSzNtf9/etxLq55L/pHK8//BUh3xck4DkJu7pyugy
fjFc7XzsF0e7hpoiaEbARoxpxzLABiu4b0WLwnzQTxpV3P64FgSADs4IBwBZ0TcltaFqkURP59qj
F/bY7079+j/vTYJidmFl8eRiKxaDO1su5Ypky3ul3nKVHPnxPd0vD5wtvVh8RF9tQvR3aIGV6OPr
KNiVjpr+2h5Rc8kbpIGbxaolRwcGGccJLl0PX7UlVuG+731zeZdi6u22shWjXFxNzL9l4p/eL2te
6QEWYmTcadHaUphW/iI4Z9aPXlvBC8VNsFK7A05ZgGs9iVunM90+BDzMNrYrPo8nuIiZFz3KiDOE
oA6LmAvNGHQWMVvPUp6c+51LslbcCbN5wheUQq37CSdSVYrXOfIXsvgyVY0RWKT80Lx9lvjLSFyf
gbQPyT0KD2IaU/WDFMtWWKGywiudKwFGcV5wKHR3HumaEmZmd6g5EDs37PS6cM1iBPzDZDWGQ3aU
/yjJZ5mXPUv3xpnTz4CpNLUBprleAxrCoBh1fkDdbhT4LClsSi7y1jsmeWpw/c+PoflyRdDGqAqO
+g2Wy1Qay6GOrWa7v9VlXcB6As1g0zYExbwcD3BBYDRPoRTA8q5unMMvDW4o33QPynXjNHKcUUU1
XoivAIu/MT7fJdhC8mHu2KWUZdlwy67DpvqQOZ/60G3RMs9GzHsAFRukhnkGkMdG1Nhjozxsahcl
vQLCJWEy5xl9v7kqYJw1f9LtnqPJA2x2xkv2ze7eUdlQtqQJ2WSNV+slpR+w9Y/P8No4CppgZ6at
7HOiSlLcyucyhYAOPfThxoJyw4+530V+KxlW99y6AMoVcpAu7reqxcK/xkliYUCCrS+gp7Z3bIYU
5QfJSrJCcGYaM1hhH2f0ZS8UH4T2GRPLIda4EH0Y+eKaMd7NUI9UKjS7aab7UIdlf5OiF21U3nKC
poT5PK+HGITe9w4623KGumfhsJsuJv958er47Y+L2L7d+orfEZQxRdYOLeXtJUIB1bPWzGF9oPu5
7ZKEPK/+9DqiJXWvhJOgW4N+dZJESmpoxBfkHtsah4VOmySksSX9Do3rcqOf5c5rZEaHf8Da+dow
mE3V+/MokJ40UgMJHs3oEXEcFv/r8PSuu/Wg+2ABL4AvpxcZN7ZM9yzbGyFrGm6j44PFlwCyFbkA
YU7RDYDNW8d577BjvOZR+OpnHv8zJbJbP1D9r27uNqg6keFIGtDusjhApZa8I7v3zDPSBwNwq/40
BCg14IWH5zSJ+kRsW2OpagkjXRvXHBcw2FATC1s1Z6vJQSVEl0rw3S0+XO8LdpynBDK8z4tpClEg
c4sqe0amUnsqA1yDh8aRcn4e0UXnUIGiClObJX8sXrcirJfxQhXRKskU+E/ORRQCevAvsMTpFTP/
WCAVd9hVNVncesjZihL49ltwh6rpxHqrVI11IdiBX3Tt3XCEiGXxI0m3qBMGb6jtWSp+E8HBhpWp
bJLc0mmgeS4QV3+m18EgvYRv8AmZixGdNaUnc2zTizEiPCkQmIj3oc5rEJ2Nh881JZttJgyMKV4t
QOi/PUVBLre2YOCRloIIRWIlHWqvj/zpc/cp3egWqnIY5vImQuHPT3EfH1/VsBgRGiOQD1hL31Sr
t+8kA+3sOSvHu3bcJcTC4wT+z+q1CZE/E46Nt4XyBgMEJ1DN+4462DjbigG+XuOymYAQ9QP5R1mc
ZcE4hBJagNek1lMnpIgFJwfkZ/Nyoqg0r1JIC8GF0CimSIoPrRL5098s54Ur0E/vu27p8ktmm02r
YCxYH8FEKWEcou+AGCwe1HBfZjSJ/5s8lx3lCtLCMczNVuhHxBG/vkjz8UKKyLP4iSbqbDrDGsXF
idI13NobTcqWOdIdJvj776NdjPrYip9p+7haJPWxhziaYGaE3JgELxfdIF1QhdRn/4nfq+Ob6kbH
ikxkGnW+/n6BCRQqfaIq1IRfiUr0fYuY9iPzeygemhTh+8lM0HK6yuOD2stuyeSOvMVvhnSsGTGc
+r932ZgCX1A765arbEf5KXsFt+0cO3XgyrG/yvHNCDpU0L9FlYx3KasdWkLDcwLWImdegRJaceZp
YdR73t/CZNTZwH4bP88emphpHhOM0bIULZOCyy+7sM43snQOGokYpazR789vM9V0wN4oAQYeNzkH
CpHSoLEJWBzGTO2Cyq8g8AjvbLvcYdlXwaGucH8mzFgEwYrWm1sJRAtqSSW1tkF/wMiSft+sVZbc
1lVQYHCz7AXJobuNcKqbvea0Uq7cX07rcn+8NXrtuQr4jW7dev4NKd8+EYlT2ND+24IXhtPG+QFZ
Qx79WX/xX/pUverYtAtKvY3nnsBwAVig9Nf9VdgOsydhgCgln4jMUrPITfwE3YCtv3sb4p3BO3Oj
C1PxOIVIeWehUrUhANQAKeV7owqX+IrTMDs1AJvViUXK+iaMnGCRlJGnzjJbhV+2zawil8rk3CwS
otHbKivLWdi6WcJipe+SX9Jo5fS9rfIteoPygYlDq3x5LNGRhw3ww/MedorkWbQ5F7DpxJlEAlf0
m8VzIfKGQrD5pjwu0K9x9Mb32JllcNYqz0b9un7bYpXdTTvsnCvH8bYBMMC6QvDJwEKrsJOXIFRN
ubuJd3utS8f8YrXQezckc38bnowfqZcUJ1Iek2c3hOIzZKQSB+1lV3GCrWo1HP4hqMfdzRvkFl2E
4O3BcUl6WrXF5i9tFOFKaqSoLFaNmeV/fPTdXxl5L9a4iW1ytKBhQ+YFokVP7R+KrPoDqZveNYxk
gMB8axPtvCMOaoskWzrCN8IO+qs4LSZiIQkBEdgHiJF/J+Ycl5VVXrfGO/1tOFzjfLAgNhoLhHmy
Fx4mD8QmMj1yQdK75IPOtzT2ND1156gl/2ChnSKqrwxn7ZmSxUU17mgxufdP4rO2xH1SGicKchXr
doE3LzK75u89AKRY9m3vnQEuT2B6ulUYyRXQKHw+42rGWKZ6Itix4MBMX7QfMfGETit+8/nxsV8z
cBfKGwrcoIfMNiXAw+M4sXE3uRfAmKgzO/lj5nHY5/sBOifJB6jP46SiqJ0bHA/66RWOZXnZfzq4
Yv8xCEbY7JWSIYWDthEY8K8J+ksiiKmUzrQa6cWmcEhia1N+tRoseYBaihDgKQ+yZDmIexzxzEig
KMJlgiTnEfYzYziMqVeYqrLjg4ZpPgHBqVlmtZpWDZbl4a5DxTMlc0sVRbqruaXsrN02IkjxSgvY
cbE2czBPJbmYN1EzZDpaeSoL7Hlqi3Sey0kCHOwyiFf0nh2bU327E6Nd81EHN+4c+30CsN/OvoQk
yaiYylmrR1EWCo+zVOAZE1teLsWpGZJC+2Z2CwpsDXIykcA3ETd53wT9kyZ3CwsxmL/bJEZrQVUx
U+zrWm5wLUwlw9nGF5LPqODl86yEtRSKXgkfRFIfRjsEPqnWFQkIDmFWeb6EY6dX7ydKbQbVUYh5
BDEvpMExe8PiVa6Z3WhK5yIT0ehTwtfAkuwPQ6aWUqyiBdhmT5mXhpuP+x62Qaqs2se83OUncksH
BcHKIy2Fz6sGw3PhRFb1zLvF98YNyAGMDKWhmCA2PgdGwllhn2DivGC9eDXBrk8pEnSRCXVgYBRh
HWpJS7XJ84cT2dbZ102g2Zd0hcYrNoa6Qm2q+sIEd38vns3zAilc0SZ1LVTxg5Agl//+1BxM7cpB
PlFPbertmXcakeKAW5boHUOQfIwtnOvGxIbcEGPuLoXBUqeRsGSK3JYYWUZ5SczP1gx9bUJvpqW6
sN+9GdpNvSguepkYtdbEkcUWkhtBYabqm5xATQKNPOV3nCHGtTE9l2q1vvQVfBVa1SHSQPmX3d0M
C24kMNMaaD8LzEgJh4eiMGffcCVjFQ8n4arzq/u+Uc3MlJ8vy+dxUNbN1xbLIju2Mkt+bvhRhtHe
yX2x8OaEOTjxgKun2vlNzsX/X5bScqxwe2xHSyE2vJVmUiA7LrsD6s5yaKl5fW1lk8nsKIxNn6Pz
lWKyaRsw5zt+TikGHFycil0VAkUfqJZtytsoda09tGPY4efKcF/XBmlrUYivUU/Wm1tYUwfkkIia
uMI3xePttnGst9+e/g4PlkArYGNEjp+oJdABS58GGRXmDDIxSswOwQbcVMh4cg24fxHos4KN8U7C
Xf2r4E2F3G6JkzkW8UvUsE0JR27c/0Cu4OSeQ1PEZbe4OeVhkF08bidPn9DM1U4mtADXhIXOKjBM
2KLevhiBG3z1XgjvRcNaMTs8U4jWtgvSTbUoj2zhbwbJcsfJpjZKWmHUZy8IKnu31iqj7CR/IvDy
wrr/1KRFghSKZvKl/o7+ok2vRX/t5T4NacZMsJsF2RTYlf+rQKBDJ07mEJa+gYTo5GBgRSnS4rCj
cYRUevQusfxrkRzQsjOt/xSfn3qdPtnV+BVKtFkDcymtlkww0Xyz4eqdZBDlW/XkKS0qJyPWnoPy
VUvNcSFE1CAz32JZBoUG6NSLbOQqdc44m5wECaAGPbdkAIoSd3Ie+ynIRmpBdPPFhVVtyLd+g/gM
bQyjkpuZxNfK2UWlOp75DRjhMQEW8vLbyXxUHV2pCjkFc7JjqV0LvKnoxa3uFCPYo/oaJ4ZTgOIS
6DNsG83CDJ6OYru5AW3EuH4chaZKLIm0QvcvxjWosJqPTFksOFR42Tx+rk4oOn05ibxDvu1RVHwX
LEJiz/3D+9MG7Bl7NcXgX9MBNf5KK53h2SijBUo92p9g5TG1n2Ln3eT0areCXaUH0/jUugPe+Gb+
goKNR2r9my4rTBUPSfgny/kQZMiVfHWRbFyLXRP8k1aJgD7Kbv2qw/1fmIEE49LGqQZP3EIHkuyg
iA+B/NE6d1BdDCD2otYpzQhX9FAsIALJTogz1usp3E4kTQNaYeplOrkZLPyKMjsQcHBaQxo9auU9
yuhVD5LJnJXGTy6UrX0hWB55fg8fppRo+5ztgpFg2q0U77VMN7SoktHBkCPl3IoUpTb/fawNuGmp
TTt5i5yveTP/LthlycGB1rU/0ipBXU5gtwJz4IlUJL1S1S7ohNgvG+hQgPnIbuYbiGHauMY1eYxq
rAjL7UTozDQF3jNQV3mdlZUzONNuXLyTTxmGMxQ6SpoodBhnj+fXqBfS9v+z32zYjJn7VwQ6dHGS
84LvgSdYi7LyOjNNCitd+S1PHhCXbeWjTzCljG9zCMCSC4Bw5vpgFO4/JVce8jY3+OMsmZoSj/EQ
FFlG4Kmqkz0J9vpe66nr9QjLjgdzou5vqPnM3HadGe81NuZ/5AsuyF5qISRXzJMpAy+t4SR2FtaU
j6RIy/N2MjH6IJlM0gfNZg4GgkOPAbZWb9GDoUionGRYntyQvV4RL6NlcHqRZPloqdXTG/icV2vU
lCjPABiRvlOZc0a8z/IsIkMNJCNUcif/OaVaJK2QsoFNpjHZSaW2sPRZWbz9Nv86jyT5I3O2LH1j
WuI92ouFbLS4JPBQx2n+3SEV7GXuySrGQgSkyzn+szJE0mqg3EfBZvcjTMdTY2I2GzITbcScQvc/
Te/pcfh/F+b4ukArhYX7IBiqm7iW/nJCJDJThDjGTsxzvmDl7woNobaMmF4C3SrGHmf60mf96e+F
76Gk4zk+dKRiZSjp2+IL2IPFa+2hlhiqqkS51oCQE0FPg5yNMpmM0z2Xfgr+XSqpb2RBTyrawO+M
EAE+h1rCa+HGaXXsckPnKfwGUqQQZhP+kqBWdZFmxjjHh93W84+f7bDHZi5v8zeqHBL6wFP51i4o
zOIBhaMASj3pq4eSvDEnagTOIS/YE3FNoUVYs1/mFWRJsGG1pK0VSrrZPAQxSFNUXI+FJORfoQJV
KmQ8BA/5oZXgqLXVLhd5EykGGGngZ7bLFudAN8Sd9HO4puYH/knjUjRUdZDfnPh+aeq44WGjVDFI
cDYgUz9dZBQ/dcwKYWbbdM1MqnNsYwlzyyrQrxK0irn6bGlNNpGIIEythYhsUpDQMS+JpXTZ1Eoi
5kxnLifHOEtSVct0i+nNYQH7anZ93Y+0Awzm1sxX9jqbdgRSfvO5jHRQDvmAUxtj2Ex2HFlGrtdo
Ty8zGodByICvpLxjk8LtZPXzn0/pxguHd741im5R5/f7RwTjQlgq8Gb2vgaKn9OPf8fR2vU63TXZ
quuWIDhunIrqBsg2lv/4rqmTLePbvUKGDPVd2VQamrECmOydSTBShCgiJklOFGMOaGhisdIMtoOG
XxlptumqiJt6eLeBhTqKsZtatdgp+xhy5pRMlJThIlitiPIs4R3IsjtPpnovuyhTKiDmKR8Mw+/L
s29St3RcxTnGEkM3zgK9YEvPwYHYevsKh6v1ArKLMoqdkTlZujkS9ywT3nlNAY5d3HBu6uHuj828
MQpDw9fnUNVUQUiCs9/N8Q56jmzKA+A3/fzaxe8axDcl2ZvnlEvY1jgKzzGjdn8BX2hfl+x+8ZOy
wesfdqcwiYCH2SFj91h902bcxHxxf3f7g21+NBZtPnen+pzym0aUHMXDvcRVwHTCvtUFlNWHwyS1
hZf2KBLG0MKVPYYpTCj+j2b78lFNTceBLH8Px+8l5/qxQzFvfRJZtq6Cb8OeDm8G4KqiEapUIiRG
rNIKhYaLf89DATyWKkKSk6s6gyU33yi7zuIB7s+gHKn9LYPkfq7TExvyzj1+ikcpq6E+aZ0QRl5S
b/YGDeDGmEwoC7tU3z3qZqhDBWg59o0oWENFqzbmik7qA+FFaDxQCBC53BV38SU+AwioCPazBljG
26FUG7+rtvmDlwSrl77i2A1MyGZwb/Iop061Ywg3/1bUVhsJ/GGtXA/mAcEk5aN0gglziVfsFhen
5JAUFbYofRMahVURM1eSWCX36Ghs5V/f1qGy2Mzd0vPfjdkcb6iKA47YBHOxo/BGooUn0bBiAACZ
7nLWK6zlw8/ZQe/SLD4jtH6NmBktIHyiEStO5ejriTQlvDWtBbIZ08ueeHc47Gn720XfnOadovw8
XWe2JqAZUMIAsTeDwCiuWv7SpCUtix+CS1x16ieTUlXdcXTlLyKvThyGsJSwqXJWiAmw2OCekhcc
NXugTQoc7ZOxgMQ453Z6gVAZ8I8YPPYkdP6TiAQdj26IzSdWp2HsFp+eAM6vfYgK0Gp5ZD9Yh1eh
pZla3oHwqLykKCDUT38ntyXx+kEGliGvz0IMi/8QRmYItRxTD9DspyzEoig0OOUrz4cg0aqw1KXI
kAUgxwedx8K9iTXHDOWbcMKbihpG/W6dpN0y0B05ECVEeUXwj+ByFj+7npUUaUr1vj5CeijU5ook
B9F+a5BDFjaurMfb4oc9BP1LKw+nVyCyfLLPb8HAPhWv3Y6bOfYqTz3llK0E3hRoJVkBmbPPrj0L
jjfigPLafCCX7oQeqj10jjHuNZ6BztZxy6erQtuiyx8aHxG7weDk6csY18aZaOpN1YlZRRj/SyVV
P0nv8sEEpjHpRc5hKUuDfxdbkikYqmtXubnW+IWz+DBpy3/2hPauF72q6zQBT66rztzLeQaab+zc
vhlVN4rpnnjHa/QMqiBLzSC2DnPq0oEvhayOldHYCWTMaXhTWqapYy5angNs0577e6wLKkw9n9TB
4LD4Yt6pZaBIBaVQDB1bfJ4PtTewe/aFX6wXP0F/hgHyugnlHQrq8gfzGDZ/k/iPvE5VaP5Q+DPL
NKBaJc9/12/wi0fohMpJKVv/SO+WweQqbwC5L5JiUZdoN/wJeQ/wr+trbqGlXNdNnJG/xn2si8jq
vqGsgX5buX8utrO9ADi2MdIqYbs/y+f4Ftwx4gFweYw0G06QCN0Zf0WFvXJVpm58LyvzAO0QphHm
QWUmZHsn5OVZZYpzoS6mGW+lc/dqdmQaoMyW44HNwqz0rKkYB5nBOlTroTU85cowK19tSB7FY2Uh
W+XxI7MeUM4bELcZPaCwaqToxqm47xg7jWBm5vTIA2bq/ot3nfWPcpRQlyDZt/CO9hjfIKVk3ndH
c97zQdlRSocH50FclogF0iVhIDE3Q1sMcvjsI38SUhkLfhVyDd9fdensigUGRjdPYOIW/EYuTBo5
vpdaofRkeNE9AnoP7S8MUu0Xmoj3TdGVH4vuaWZmKz/w8MTCRgKi/9BYmBOFenwD5b55336WJzZM
J6weW9iIdwf8nfDuCedEQ8wjvlTYqMSS7HveoB22bzKVo9x5BPpUqUPSANWMHI9AHM8DYLoRlDpq
DvYFex07sS6eAdcN7/jInRzgQhJdNL7cDxKmoSA1dMEGTBI0c9O486K1I6tvaKs/xVJhzLjWf620
FRriSyXKFzGqQnpd3JS6Hktz1sfGYseivEKdHeHys7xq69U2JimVBIZ4JHlna8ieczveYykPQPl7
XWEIiWbLKFlWVEHsCiDZAQpuYIEO+JsFfZb4meG4aEiC6HA2Foijo3DKigTpgCtZPXvpg/hqTZk1
hL0ggUA3srEwm5I2ML6Cas6pAPVhNp/Rgmb6pxf5St5OuvfZzMnqcrJpm1UNqsg5TKv4rVvJqSd7
+aLrLs8eio4jm/CBZg5eM6oInCdGJByR3fdt6AYnnwZqn4bQtrUrvuRD7MbBjMROZ2pSfunvLqxa
Mvj3kRoAYyC/488agay1W6upudkWcj19aXelG3HkJBczda/zN0wjueQ7mavWntl+uB1t7Yb3KoCC
l7UQeQjIcAIFAh9XfFUvnKzEHLbMCm70aN4uSrLGpJRJeM+WJXO8wUWq1M7jCc0p/GqZsD1O3gG6
j3SFLp32FZr5rhBEcnI8Ft5WCPDMbqlHdKXAazJ+3TBrAqRdO8lq8BkMgtjPYMlU4RVXjmQpU3RQ
Pna3gbpuHkwmBltEgef0JJ4wx0K+cIbudCSfRoDMrQXj9yIUR/7VG50594dWdKp25GD33F0ZLjip
NhjqifzGtnWodL7IVfsyKI126PNvF91fnY/CAxb6C3dlU5pA8bbuiNdpj/JYGbHOT8uoHqglE8d1
PLRgFMIPg08nxNv97WuJk2OcG7Wo95nW8FEXG+XtEqjcOtXyD/73JF31h3mNBMeXkVSdZ2rXUVnp
UmuJJ2zq/YyGS4fp1iIf8e5xa05xdM8ePJff4IIiqx9QRRa3sQObzO+pV1WBQiua+UK7XqyQS3Ie
ALoBwMdV4GDK5VDEzGdAAF+rjYe99xEkVKoS7S6NSzb85uQAOqBjxn4y84p1D6Nga0OTrLCojCIT
gG6cDSFWHQ8nvYthizmNfg2+9+mTAGOiTFgRkrj87EOr5bUb8dKmp9lhpdZ7/70kzHORYWrjGcCu
BjG/JxkNjadgmFMDXAMiX/eqvra2J/jw6/52bqgJD15ShdBy/E+eF1W1kdr7ZFi8sgjdVUU3FZFn
8iu/SQXz1Ef6iJnHPd52DRqymdunF+m5f4N9yhnwyNR5YxDcD7GhpxmIdOKEI12UanyCRgfaIdQX
fH+V5Bt9Xn+Pk+/s7GcK3nGQjXP2to8siuFIyz2ReMowCXcBulwiNOb32a8zWt2LOMN/VPkBckmL
Yjf8XCNlGk6ZZMoZOV+7Vi6rZnNjpLA/yegSZqFR9/xvB+O0RVOkrCn4aaC9H0sWrKQ5BmKT2AI2
03Z8RJynqVBTFuQgfQDUFoYSHIg4+/Ky1XqLzIlO6olpNIFB5YFC1T67zyRXDrdAlxAhBIl7hrxn
LxDeit15otDKivHYZZHuqwgaBtjVsMekc89QteS9QMdfLaTnlVCZdU167FsN3xP9zCymTf6lviGm
/y/4MrDaKQvhC4NFl5F8HAmFraa5TkkCm7vmoAzt+BCu1qfKTAvyq095PYZHB/oTx65BP6Qc7Asr
PEVVWj7QzeqyPFiRZFJ8M2uf0Iyggy5ruFyfZOxzDTN7GlqalThg9TmvUamppsZVtqSjcQp/48py
4Sw17Bz6SuLQmPN9hZ9oGHX6o37jO2kuoBFFdfpiCHc73NGs8LUxkk7V88JcYS5nzvtFbbqavZOu
SUyzENv3bRLfuMb91gFSy/l2Xq6/KA7m+AO6JEvQfN0mBUmVY1BeITTPTjJayruj6Mshi86mzmwQ
wRnVCNOy+M2zEeiRtg6Lh3HLC4rDTbJOzoyAJRDf0isdwBBttMNzM/BHNRWzotcmfsI6R7BBhxsH
6L/GXXjkUF2crl4vSnN3FOjA18vZlSA9HFWgX+WAh1MPDNpwbwtMvegUGDo8baxWJb4vKHcrL2wx
i7bmVaoHC8+WVPx5mgUUusf8tLr9Co9k5HI77DjgbVhgmmWaT8QkBSRePfyb8iD9zLdmh/3Bp6IO
rSFwh5YYZbaTptG+93Iy/Twy98CR3oDmpnkIIt3O9yqjMcrVOcGtI5y0A4pYqv1XbjUAaW0pbxco
y87uFb4k+g2zWZ/ObG64oSWgBBYBdxPCzsWbLxnoQQ62sgqUOf1X4d7GsxwcoDKZNENiItTPv8k7
WicIsMV2re/xrPO9yQD++l4anWC0TsYkYkrpaDpI2FcJSz+ytdFiWRCMmHoBQPeYPZY9WtaUXa5O
3oVVssNxT6EcCk5X3UvsQsqQOcpP006K0YHixdPtnzpypo1Xz+orY+VPW8z/bQdMi1fySOWIl4sY
oJPoKrPKgQicc2oclLeJGet/gNDZjODAbkVjvElacMGqStVQjHCEOACf/xiQJepjpVvj+HjKw6vP
85FXVBzIR/rGZxY/R39iTWBVXqc5HZmY9gwf+ALDhCTSkSPaAWchR1ebc2rZ0ISzU2/PVyx/emFm
6HeIQ25S1w0kLVjpwKtG2HVwPdljlvmpYmqE+tDthoQ8SQ3+9YWNhN/E1YKjc5P727Mphjxk4kAO
Ig4DK0Yk5UfRGctkHaBVIr1PwWFBtg2d7ir7XOCbvm6uzSGVrygV1yJRIUtZz12to6upuKRtH2vz
kPkZxlt1D97ckXWUDp1YnNCoq5eFXLgkzoQzJxlFF2iJc3qZODczWjzJpb0I1/v8s4n2vQO6B/bK
aSIdxzFEHiDAlTzExxpj8M0rRZAu0xhMr4i1uzEZFtXMEBFFT4fnoAcMuBcVhk1AV+5s3ISbCdnp
AxJTainl4LZEbsKsF7CIg5zRNzhhIvIWLsiDNYcCrlpAScgJkp61hCqCWnblDYnNF9tTOxr1YgNL
786YpDFSYhZ2I16qGvbRGOk/zcPZCouiFOzqKvCN2nuAJZF0TzONlPQ4UzviqRpX/6y2NiQuzSxP
wl8sdHbpxUPsifw/Y6DWQPpK0WmucwJQLI0sAMlGRbqhdjOU/biDQfgI5xmMGenmuzLkpltksMsC
6dkVIDDu9XHKTBnbJXW1xK9Zl1uyg2l9MViWe4/SMCyPUIpRjx/f33z7kzgDRJX544V6bOl3a/e5
FZUwqrwkChsLp4Y2OfT8EOCR0RSsZRQEoaA0LL1ST2iPtIvyH/GP/ua447qV15OOIeznfZIu2t/k
KAFSBGNF7Tu3mLzDBZtN/nZdEmvd1+661afX6LRh3lkjpWxXpbuzUD//ndj36tI7PwDK7IaB67rO
XNvPnazDe+2u0YizUQJx8WIHbCEtYqD5xwSqPNeES5BRLDp28sHUiBta7GDWxf2uhahurYxSS23P
a/2E67QUyvZ9D+IiwyPzZBOiWN/mSI6IJgyFZ4iR8IAbIcKuc9AKZVj4/pvDUErOYjLZECQ4T/0Q
ZgDFLWjqT2A3tCFJSmDN8YE6k99yXly5xfmR8TRUescCFFF8R1LyuKA+OEBBr3sRbHmGvPu+HxIx
868XbGUHfDUML/eTWBlnLHYcFyfjkfElgjIzi1dqrMNme3pdoR6B+ABEC/r/q7kG985FomrB740F
M+Xn7UglhuWBn01NCh9xodqXcDMluQKGW/kRSSqO+YlvohZ7fjRrBbYlOR1kIlmQPksTc6tg4vjy
0+4k6yEbASgSi0JPxizkrfGSdly+z4L4QJ+CTBJ5tbyVj3e55rIcwvVFGl6mJchv4S84NthJyUyI
IH0QE0kDoYzQiwUZ0tMngnPmqv4ZosdxpD8YEsfh3CqaMv+PI5QDSdpJYRDLrbVLgxHEWzPZR5ni
xBasW+b3e+hsl67E1faLYgspKQ0DAzsqzP0bNC1iY3pg4e4F23KYVjUdcRTJQHCNHpHEIoX04/0B
Dg3ah8FUxYvWOV3RrsHnKnxaBuCSx+xgWZHaoWMII4fpl7MCiiHquJ6zpc9tHcbBlPUoSAsUXGme
WhCcGt+efbY6s6SznUgaVjL3wce5p0JQb0dw5JdqSG2RIEkpHutcQ5GAE4wPSeUeHfWFIclHLFaE
l3xC7oFDX7Hx6vQsOProgg7t6oLkdqZaH8daiaR1tKm8MwXRFS4u41rLz883YB5WAKJLLMOLz0Ra
E1KW6x5zojy5vU5qNM0OzIYaOSGGsieaf0dzZ4TjhG0CTjZuXUgztFtxS4QWUOUDgM/D6Sql5agm
7JmamN1B2rd9hEks+C24rnRiUOhuDZmOcbKyzcqhoyU1+64pHKyJkM1819yyS3CJ95kcOfIYwDoR
9+2YnFBwRDEvBFJ82a2LoosWeZVhZQkQb10egHf4/SeB8ifwjb14YnzFv0aKA1IGhAl5spglwD0X
3NP68YvlJnegaPYB9IIToTuQXTpa/R+xMvfZXaGHo6AQv+2qAYutfHmd7HRuJ8WnSAKPuiXCUDqX
yhYROyJAny0un1qu8vEFFRnXcuXUtdNrPOOyl9sb543Y7jH/ND50aSFTXIGaiyq8OCaiwYDDA0Lw
Lnw+BKSywlQkK+AXtBrwT2/rhx8dDvD5u4EUO6p5JhlM7AaXC8G94SYX/1E3tUZR/6Q5zCGWxSp0
qC5TQNVF3FURR1vb3kXx16Ci4T40JzzOXHGvyb7k7X4NSrQt8f2IOs8tjLKWXrFHYkVpL/ZwaXKE
ttTv94f2qb5RBGyPLtlcqwLfekwbppoZbgUEuYcUpSgK1ox7/UH8UnmQKN8Bj9OSv9+VD71YVU9s
EG6gHYyVTXWC/3YcobQxcIyaiRsq3C2hV7AGtc5u2jxY63ig7c+xCXdLWybPQwXHktp46DHrV3wE
54bskU+4ATFzwADEIUa5g5O/SLzCimiqB5VBmkpVbN7M4v0cMzXIcwmiOI179J7Z8540G94cOnE1
6oi3Y9ktV+X+gg8+of1CTQ1/a8D2QLx65YPTozB02cGEpyH8sSlD1d+FM4O9tplNagQwfy9O6WN4
H8YtHYg/XmDTohEVRArDaeeorJ4Q4Nfuq+r9bjtC5tn9DjNjwSfFMgQzCOH41v+FvrIuvLZPvIm5
RHXrOgy5sn7nxBZf4wBn5hpnZa3AkeE0cu0plW7ZXUA4IJGVOlImnaqfjkqr6NwuGSoTXyTRX4XU
zsEZ0cEJ9XIulL0Njh3pUmdtYX15YjhxgwYoDCF5ED+jyY7QoLz/qCh7Z8ZzgfDcHaRK7BwLqgg7
NBoPZBoGcY0QFs2fYXgMXbuwn0hfFzQCyzPU8f/IAMteZ59F7uS8F8Vbc+QLX3iw5RKg1p5p8lA5
CQGWkvjiq4uMrO9sWX5qRMKD7vc7gpQ4Zj5/UJDlG1QL93coxghpUwUgWU36zT+Yo8mcnFWbhHil
r2R1gj+D/KV2ZfyXLqSTKiWSXwj6qTVgC/ivQkPaP+bzIqldDBdT9Ys8dqVLNBeNxLCNtHR8Krb3
5nVHbakMDSRBpmNJ9tqiQip5pvH1EhqkbGSnaxzzw48pwHo5BVmUV3Puz3+Jw25vpodbgwMzrrH/
zjWrL1+beJxdy7ty6Sj9AOJ299EQMkLy6WR2+DUIqnjEHNO8iDK26W45FavLScxM+DEBuheIoJKC
0U7hirTDNVenENunodbaCdbteT0PZMoy+RWA3FAPFS0LpO5ROxJHsxMj4GuphP4mDqvbiA2UWvEf
vkQjzzM+9JxcSBbDikIFiADwi9EdDSM/kSmZlSE3NmTiY8gioZ7C3WcEwwrjpCkzGe29g8amQnyi
GwG8bPTkx23gofbziOWe3cOdAAlf+hA0KBgLHfdBsk4wnJKbUlQ5hkYZ9mgRqdv6d8WCXJlobg8t
i0CdPGuraz7lfH1dLT+5sGhoplrchxW3+s0m1ce0WZa1QgQSXDc6NFVJXiifWk1K9txjcy+KAtBp
XmSyaKpLtPpCa0zpmv++mAbAHpFxLG8M7LDBfIaK0RkVoGLkfnEKhHyi8e2AY+K+p3dB3U4DKFLV
6JGa9fUeSoCi/j1T6Paz+b3yLYkP4t7CbKGrHmuEwcP5ABz6FtuX6RH3kZyWPGbFYFaVW5TOQbfX
fQuuDjsBoAsA9RyqkX9Bn8NEzMYvPXrLXs4zz/t0qDCoujDYyc5NfRhz9J/TG55jNvt2ZnkbJSup
NwZPhxmzz68d9Kl2D+fctR1UkJdTP1rkMJpzn4dGE/mSF2H50JY9nAg9HqyI0mWcQUopT8O46okA
knUQPzsCHzB+vwgtex9QYj/ZT18cWBjlLHbdjv4fcTIB77nb8sqk1jrmzD5c4ML+SidLKot2Eb2w
nWf1FhyvDlqgcMpxLjTWJGmie+h4PmNnni+xApyULere0uPMJtxmZYM8IIYeu3QulRMIl+xFBN5k
zYhFGSNgRFTncYL6osS3N2dRv1WqpfFZNDUZpG0DEYoMx01WsvDsTTN7+Xwpa8/E+487gEOzCiWz
uzjiYVit/VIf+FooyKAn2P0/FRKmQPrJyGUuuHwWTRQW4PtA2JoeqZAR+iGcRw8LGvUkkR+7WutC
CR12gVP4HwiqPS8+8CRdgjljSE0DLmZ9z3Ghn9EQU7riQfy0VZIamQqFEnKAUIvnvg4tTb7lSdS4
tRIAZUJ/xZpEfajU3E+FS1oY87a4u17ZtVtIqt01Z6iHeeKP7tx2+FjA7BlEQpVrQMccF+C5O8np
HFx0+JAc2OVEcLjw/fH6OQXs39xNdRHfwoF+zmRFQymbiqi9DcE0uMosHkmxqMnuxc/j2S73iEWE
7Mj5+MVqae6btgrKUQAJuz9+WkgT9Z4dtn1XQi6Hy3gyiNNvHaTGFZAcLpSmpA38zYHr+UhUUVWd
Z+leTJg/DXQM3+P0WRTFLniFHvL2S9CDSBDeOJZmX5mVWxLB8x/6gm02E6mFkXlCUONOLO1F6sf5
GbRHaO3rfGqthNaIdF1bJv0TUkT5RG/wVDdidB7+7ubrKyp3zTY097EAi08YFvoCyEr/h+mtB4e7
/bqYC7bsMeDz5r2zpZd9fd5D8LAz8casr9E16P8/GF6Hq4/VNufVqEINX/WeSNbINsuKSjpL55iF
1fMqrylPj/cLMrEJnt/K+Gobjs6MKED5P5Ri8g0vegfhOKEtvgkt+inzhG35PssFM+rMy/H/UN7f
Di1No0aeS6LNkedyrN/iAxB4DmfKVZHDp0yvz+MTZIUkqkm7okSThkbLsIYvKHVsiP/O9vOR6ZID
6Y5pAYA3NqhFkEEBs73A00IiTK3fsIeir+U+B8hqgjOIfH/VhmbhuvN8tglmriWwCRdsUtDuxYmj
pqDwmYzkt4tx3oL4RFYxjZ3qzTFkCoRI+95KdbBsP/3zsQfoI3MQD1ROeS7rG31yX6T0FClLSPge
PWACcuwRalkEXgkqC1nRoEMw9YrksuoXIqm4hNG49l33stv85op1WJHac4zGyzFzUI/As0m6lqM/
xBIAwzZ/tDwOXYIY/mkyooNH2tcdLtVW+8K7aOiDyMUrWRDp77LLklw7ZFss00XPhUWY3/uv/vqV
tpRpGc+fCcALOcp/D/id6R9bXOC3HttsHO2XQaNYjIo7C1eHcqwXoNq641hQ8AHaWUUPO+ZUwwk4
ygDGRPta8XN4eEwf3WTf9tnwh1rFHYasb7E8WUWbj6PELzycNNPm96+f6xTjLtz03JpLagcQwHlM
pYcS5IICJR1ro0sbKv/LkZKySHUjF8FxaI3jTkVPqqpcxt/4LQ0XgOvQgEh5UkZpT9H9/3WOargk
LuPyom+eWM/fOOuEY+qU3wZOOduaNPWJBPMgcsgo+pMLO29nDst/Tlh1R4vtGb27XU/kNfhNylUx
BjPg3hAh3Pxk9LNPrmQf9qslW17+bidENOEAr2myHFdTX1Alu9dHpL3oxsMx7FhsFdCjSHKipwGH
QH440kYVy/k0qr7HshEu3w0Qq6Vxov0Xk7yYmkEtYpeoqUwR+8Lu7NMOrKN9OehQkMNy1G1/ZrIF
lVzeUA6wZfEszUMnXbDA45S1SYnf5Ic2/57HzktSHdLfmyP0Q0VSrnzFQOv7fMLJe7zz1MXIB+Lu
C+CRFtd/2GpteqgfG1eKg6UgxLV24DUB3xQWsalnI9frW7cUqAizlTMrKoZy+pMjalhzu3J33I74
oyG9uyd8pttB1Q4lXEG12JP2P4ADhWcwgEb2E1iLo9TRPgdbn7NnRSYGzdKgg1jmFdfuMuU52uig
NpH2AMqzPp6HP183IR/4o8/kVc/yP13k0EriKXx2b5Wa78B1OlY3x5lHPs5QyL59azGEs+LiiFHW
V4ETKvvLp02gAyddbJKYamw3fic7CJ5bXhzexOwceCIR2HWT4QMCzgSCQqRgsTbbe/BZ+IOiB1Om
3SzyrvaiCUTM69Tyjld6HSEvaOqvDWHM3pVJX2JzW/tI27lvewKehyjRTq8h6qYDSAbUQHxkuCkk
gIM0r9rZQqlrmW/THrNldNquZh8NToHrSC6kNQ21/2w57SJwljGjghstvwCRBw9Uysl+8QkvUAzv
/LbBMFmxzNNHwApCaVIs7bK9q2f+BiH7Ztcrs1f0pEUODLM7mo5o/zyQosnpIm8cl4l8ysLohr2c
DeoQZS5hU43cVugHEC2LmuGIE2OFA5ean6Wq5LdLpJZ5Vttxiiwndm3vqvsHcjwgahtJmpQkE11R
uESELIueda8y/swtgTjXW5W4k783Ji8ZV2qnO2jLWRYuYsajlhpaQ81U23kXyib+dhwDjvqQvIFe
FLhD8KTqdYq+qZ+ooC2gY4OXf/WGWjn9xJ7uH0JYJxOVgisvfb9Tu5dxNMX0jVw5q1koj5i0tXs+
72FZShCC2mIqdojqJISNz45ucGEkPjlTBuB7RJWhe1mVzG4j22kQKf34x5jiMgCeBGYs53YddAfk
bBnAMg9dRXuKUAx1otjXwboeLtL4nd0Bhp6ZlfR57sdyQKe/liqKMaKqQhWZ6BzC+mKFQfMbf5tA
lZ6/H4ZSHdh1GFOBdm+vrX8GxP+X1uvBYB5ffxveTcdc/KzRZi28PpRJi/L6Q1vLSglXjt50/xVY
mwL5w3xDjDEl0cEGzbL5Fink55EJpo2d829gAAGXiMHKVvat3Dy2QSo7/McFRwI3qhH1+lnen354
GemqRtkEK44JFvBTBI5C2NvfhevhJD/ZCI/UT1Y8Syc3Nbzm5u+S2KYn6PsuXItu857Q6jFP4A0A
VorsMvwJ6RPs5efhgS/8UH/RAl8/EgwPeYHffrU7m1NlSPDTS8iTDGAL479Ux7RRBn18EYabZz+N
x426DUq8F+ozCBSLw9FIFcqR8Hkiwdsw7TzAG72johW0NU0gw1zxM9EU9XAntiSPkjDwReKF0CxP
lhJak0lyNfZyEa29m0LY9+xS4K1xvoW0/4xnsixehypi8SeJHGYlQFmErbUS8M9IdOOB7S1kXF2u
kPN6atrSY8iR8sCHWhx4s+Wr/YRzp0/YJY7DnaEZ9qaThQEa56R+2jASh0Tt9mwB2wyZ5WPpJhgC
f0nVc92ulfHmDCFeIh70GuvP/0on5kyysrMjH0g6bQPlUQOSW8NDdrs7/m447ZthT2bR9L9Vm7WO
3E4U1XA2oLoQyhvh9fURhiWfYue+aBHebOmLqDqeD94tN9HKhuJ+xfHnz7J14hlVSHoNAw1Lduxc
6CLnPV/XgLk/qoSZzyPW/nmfGDtlvPqgyP0jW0Zkel1N4h8P66zdjHFCotH/A6K1zcUvgEhGeE19
4klTlGGvkg2jTJXl4NX+cl2v7NIUcCQhRwFk2OnejCweLoo2X2hhbR19FpSK5e7YpCPP1IuFclaq
XvK6orqcsCwuv9U8VsYhdOc699R0cQGHdCVMLOm4DkNM77YMtFJdOGF6uCM3bXlqR22yyAW1kPyp
KzxTd2IQ1l+GVft5s8W7L6BMHO54TtCFLgMOa2XtHwOaIfR30nGRXJhGbmSbjljQmmU4ltLPzWee
S5EeXR7K8LowRspUrSQchOgn86DHGoCDouMYzeXwo5SytcWxgvYSCCHHW0RYd/ls3kop94PEzwIv
V2h2i+F/c+TmjWuqQWU6G/mvU3CIWTw5wXlgD3ZOdoBzXXBXO/rJEw4gzYWnju8JGsQIfdUVBMwm
NlMQk2f0N6wNPFq1jlbbPcTzkHu5zGWbQpwHzHfGvBOuIuwqOdo1HWnijGk4ZawWcXXbpv0rJR5H
DkmZnfBWXXxrPkR0dDMoCLqQhIoNGnoflnH58oL7VXOXThXUQTyqZ/G7XOeXlHzfj3vv2T0EZKim
KXE2f6WdlqswJWT0tFN/OrMruBkGGIzzhSVxIVvnmWXCdkuGVc1c/sLD8M5D3P4JXTOW25u6gdCu
txL2mpqwAmfVUaLnJcxnpNPRDkclIUIOgeAxgXHFlgJCTONR6rdL0JfhMjz5fEdPCX+VTvv3cJt3
BxRlOK80tjMgtaMAtsdEVncXZzZ3+IbOrRu1mS3Ibv11vUuxI3sbNEjP0UjsYIIBHwz6Nk0u+vlr
9RGMex+fQlRusGlwPf+EA5gL+i7tIwtcelLqlqufkPCHSRYFyywHmGg11Ek1/Iq/7mVGCpWJtGXt
BahFOWLB8w5kxIMzArUJajkM50aKGvvikjUOPEbvPXtlUoASMpBDBs9vMxP24mkUqUoDSso0oj/M
+5GV2z6Nd6tUoCcf1cpD165dh2A16UbF5jJmIwEVwQWajNJpsiiEEeOK8i47FmdgK++5gI69LaSu
oLJMFtVPI73mN0LkuB7Pj+P4TSZjzJPuf3Y5+JVV9WW9d3Golvg4oDrm2TudSELrV7fjRi5lFbFE
ajc8OMKPflJADQQahFcFfGxKC5qJ71+ovKVz2CIyGy3G/LRO+fQWzXE7eu+DjGEhXC72PntYu5Xh
JFcSy3fsh9W9sZ4OvO9T86D9SvuhOMvqGsODFR9UdFLUfOdbleLfLg2GVWQbxXNavwhz2g3JICPB
nqrV6XisQx6EMqJ4vN7ZU/eWzFXk2HuuW7YE+T7/3r7GpyOcR68qVX9jjdxbnPGp9aFgzdBCRsRy
+yw0iypggd4oKcFcOfKBWwL38fhj7Cy6yhNsBvMX2mHbJRGE8JTsAgfWr2OoFEYt+3oHM/+baEvt
Fu4I7Z4L6DPXufKJxqr2p3nHJ5ff4VeVO27ahcoslO++kyCdl++73SSPmOMMm24fxgj+6cjfPcCr
3FqV6yNmhl5Jvtx3jOPAi9TheFxPL3k8dHjqjZmQT/P6r+wgFz5EJdRa1fcv5aIitOSwxLFCbROx
3qTViD4JlH2BtZwFnQxDJBlLaS58CiW5+EbfdemUFIAScY7EYdcUxzz2p3GLiyugAryBdJODZ55d
4HJP3vf2tKqUiP49EsrxT/oN4LwtdScucOGpAdPlt0LH0g+sOXHdxk+OenmYNE7/mUUzmRfMiNn/
ChO03zsg3oEftQ4r5mLnjadC/TDDCv7dyUGB/NGVRRYcxPu8VakbBC+jGwqyV2SdkLRcVPrKKXJf
XIJczN2PvSMgmF6aP/DRLr+Xd4sSmw5FMSVZnpAyx5mxAcqUK0CFq6XAwiYYCzanvh3lseu1gxjc
VroPfPi76inj6oUdP3QAhoyh8OHTFay6olwavIDRKLehgNzWiUA9PWA8hitKgAYZbZsi9G9se9HU
pP+2MdMbjy+wezhbgPlDVhvcPT9VSnZwEQlgm0SSRvG0pE/A7CpegnWcCgrxyxj0rkcHWF3NUme6
83T88xi9DhKh3Rf++YcglrAFX31+L3J+nIDBZIGorKygGso+ygCZZ2IdPp4enY26g3QSyeD9O03Z
lO7DzhHwnilCU51WfgLbke/W60FyDmUuya6hkP901q9DxRkWX97ovRFbsRlEOMFYUBc2VVi/y3ye
79X1rqwCBdW0DKukoLbQ4wmbavAva66QBfEbChbg/fGgHGy59TdRum9B7oJIPUSlOcOSSzIJVZ1F
8zprqS4FRapfL+Qx32i7ZvMmA5L9dljkdRV+83zNdaLfDVjyIgunizN2Y08IdtugVeIZPWjnU+s5
M3Sr9o1SdW+XNUhTWwnH8qxi9MqwaeIL3kGP5twJMd8HTNPEc0LXEze00wy0JYAkfOJhSDPssGVh
1r2VLr6ttuhW7rj0T6gPp1WzcSQcvsiRApxnE+aaI1zjPWOHkpu3R11M3U03tHuuK09Xrzy2NJWV
H19rKgKf+6tcRgAQ1+geda9pZ4aeKM4q0R/cyRhlxRt/6fZqizDgJG1ufWjhT2rMhyByvYKxUDJo
MoH1xIieIM6fdAqBM07I4rInQYekmGv9sO3UnUyAW+Ih927I20Nrq510fu1rGJz+natcPmObZyDY
Sd2KESsr7vzTGv7QcQWv79xwSsOEfb2mB/J+E6torXsqANdVdvPqBXj/XR+kJp0hBXFdHyu28F5N
CCisI+4mmxkwXqyhlnjnCVOfHKbBsXwp9HI9pN1TGuNakkECa+A4Ii+/ixGI3P3QexGvtNsIm1u7
cPnTQ0vJV2mYc2+M3oKDro/LYILViRTXG6f82v9RC8jciZ6PPD69kh5rz/fHIFiuv4rDPeqkbdUq
GPBeVulbe750NBQfTEGD4Khg4zOmDJfiH9tQvN6OXSK3SHnDjmQK2MAMid2gsx1Kdzb0blqWLWuM
rng5Dbs7WsumCCB981svZLLaJkvHWDfTLlOnrYEXiH/UOhUAqO+QiSX49qd9Hpkp7R79CMVnROVm
bIzwGBeb3Xt9DIAZDt8pi9m5bNyjxiDb68Um2xengmfMFvgFW/X/g18aBMn1HLH7cKdrGjaVq1gK
iyKl6D5+6+L3LTHqXwQfQrK1GMgMdsDhY0VnIJFDWsfS8ns6iqhfgjmPbGgIPTcnK5lvQexsYmyW
GaOCvc+8BUMW3dOcqElljCFlgRvUNIhi+yMPIMimTZn7S8GxEP+PzUuwi8p/x+zv0V4cMoQYTtmJ
SnqJG5Z9NuQrNsYktUm72eObrKY29P+E+4ROQuVSsU/6r6DyTxH0et5ujXFXiFVRsFgjS5HieUS8
V3UpYH9zFwOTmXysd/HvG9Umc2VLcTybZCNSZGYlhVr9OwlfvwqzpjUJx3PF8ExoAzM7J6hcDGCu
n6HqvTfSCBXi+kilLQ6VrCEme4PVzr0xBrQnIESg2f25rFgCKpJoU1i6bfLeBupZI5/EBAlh4IX3
hPEjixNQxstjPd8/R89iINgKcqwFVvXxRbzdQ2cM5ByHz+OpFlUeqEWp1ncOFhyQLydNyDRTGtnk
ywmARfjUB0Ii9LdFPgCIo4btM1v3fvuwFR84PPHtvOOXpHHxNIixpDG5b4o/Kv33DF+AZEvEIHZe
w3bCKVIGNNaa9weaK27KgnoiSwrToo4VeFzPfopZOg9FRf/A6IhiyxD3NRt06WDqPU3/62KWh6YV
Ye8sJyxXLzk6CKK7ihCRDwndTBy84pFIWi5ZacoBp6MVKrtFIkvb0AOUARqAgA/O+7UAfzK/jtiu
f0Q43HXU16geRql/yf2TOBCr9h5tdU7OzoFm/zMh4l1EXO2XJ650zanPwWjluzIuySOqXm4Ipphc
n+/wYWhR5gjGfIbUAZ+xybcSGQaYjzndwR1Xlf1BGlRbDgDbZ1DL1UAxaiAt9X3+66+WFh66OHm6
ZAC2QlGHdIJPrWZLoTJAaAGL73Imx17pqchAYEgBaIuThZfSiBFQepJdaTKmIfBa+AtP9rgqNS2C
ERsarEKgj2FgdFwd6gCSK8NYPGh8bIfWeHmK2nFR9ZRpHygm1qFPPrFiT3QNVUCWaPeeywIIU4EO
oFtOhgay27Tf3jhJawd/SYleBDD+Fd5pQ00KwCj8xe6kzLCYDFyRFYr5fZrTPo+35WiztWa37uy/
tyWsk7qOZEHXBX8awOKSZdh+crw2mTaDbNmp9zpFm94aYMNsbfB3b4ZX6XKBvLknJhsRWFl5uQk4
1pqU/lTkp8N525usoCaXoNaEVMJFzUPyStQU787xlzW6fdZu6qMO1qd9TV0MoJRHDkURQabWZvtS
DV+WaMbrCQa/O6vd9ARWrmL09+xZcsk4Iva6diauayuWswc8TsMgUlBRFjfWZwp+FNgfC4R5MgHG
pAW9075Rv9Vap9coIzXXdywoOIy8THFOy/f99YgtWR0/3dUrmHIoFFLRd5JK75d+1cMTkTA3Ryle
IfK/Pfw0lNOSjN7LJ1mpqkocePAe+smtUAk+ZW7SWLe7hGIcaYPK3GGJARRVOFaWZcIfwXAhCgIj
YIdRwFQjXDoLkyDIIbWB4XdVUV6SfRhCRJ0CIJMA3AmtQIctypNKYpOIVDeJEGqd0lbG6I713Un+
qrOSb0GN1qfhH4B185zMalJ19ELCOf4bG2SEgpW/i8DebHpRJzQfGqHZOKydPkOkOI2GT4ywup7W
2NyASGeKX6TdPf39TMRpvPEiF8FRZePcbQCmfP0Hp5i8pFQs1BKM7PKjRksMHRycfKLFDPg9qoiu
lZuOJtqRk0vdeVLoeeHh5ZxL9gID69KXZmeew73ghrMztHdiVSuOCzw429fLtVj4S9HuWmMb+75v
Hu2eEQ6w98bKrvy5bB0cDNFEm+CttdLDqnm7K3XAREpWqhWzrEhwI6UJ4QZ4DRuIBaBLeYraGRO0
g2E+6o/rlhf3LpEELXgTyDm/5e7Za+W7o+B/u9s54ALo++GDyvt53JPrrV17L/szcLynZmw/VZSl
QUnbjqvlzEZKwxwPYaEKmExVSVAZ86AZIoQRumC6fCEWOfgGSrW8I7+F/rAnbBJ5Y15ZXrMBTu05
xuaiDDAwBMYMcJad/cliyfMXWI+5mV+9wwD0mywBfmR1NmmgWAV6KBQLK9n/WAxKKoKFClY1ykMG
uF8nbvJVYKJIjn/geqoDq+IFNP5jXDcDzNYVIbnEAXKq0s9ZKy8dWf0Bp7BhIPoasRn50eBLIxll
pphsiGgy/IlxVJrQgVCD7dSCX5MP2uX70PygJ1EOw0exyparMhuUbIRH/XH/4MN6j8+aaShdmrnh
sgeCjN6UL9vekIQMuaGJxnLcSpzVRRpZ3Qu2VVP1qmQob4noCWVdjDrfrJRaeIyyZKbAn5h6IQBn
OCZNB7lxttkJWeUU9Y7P63lumTdLyFYZMM9gHHEpv/TfCgxU0T4ogtinFm4P2t4bsDafohj8EclZ
Z/i+qTW0pM19bVL7+RqnBeTmoJGIrSEjWx0fB5WyGQ+63iLzWk/0KxugVBxXGx/UztTXhZxAe1oZ
2lFOycdoQq317ks1RX+J00HHAmpYA2e1NHwE2/+3d8HrkipJtNOiMjGCugwLAOS79ykwid+u2Zuk
CtFVIDSG0jZpzyFumqMxZM3EM5YJ7WGd1uKYLgDgI3KnS9b6HKlikEk/jaWeBNuWKm02MkI2odKq
t1KbXPaC81TxFLAZdkE6gVUykLQylJP7fgZ7s0qliTLhpH2sB9rEIeaNwiqGfm0CJSobwxRksbzd
RK9DpYK3JRNvGbHxkYlnI0q5vK3TuKxV0qyqR16qB7ch/b2fgznich16dQyQ+5JZ2mWi8P58TEPJ
yUxPAgyu1ah0JwWzHWQFtDgDReKSRrqVuMzpRshuYfUo9Dvtyra6pfyJPYKGavBdbimuSxmFRO04
nzjJpvrl5IUeHo3kjbi5Gy5BCqbPxdcCNOHx4+ah1ja6ga9np4UnNMRj/G2yyrgXLW475Dpo3Pw7
9/j132oFEGgNe2WzzdZEHz359xdowJ2VH16dHEyhBCwkMFcrN4yPAtJ+v/Rgx6GXMaWSZy28VGBF
L72OY4GQ2eUY6H8QUU+7zNs1YS29hfX1uIaOAbYZTTZ7DHqnFXKdqxZWWn7gQKWo7Fxhbcpzg/2s
NsgZq9e57llpg/80T/LF9z0p5101k6phAb66JWx/v2MsubV2mSwtGBMQ5NxEkIJP76r5D76bmbWd
x2sGYzU/W3Is4tKZPUUGn2jgZcaSEFsxqEixMGYvxBgc45r2OR7X2GmGbSwSTE72pyAojnL2ZUTm
Rxgz1o08ky0B+rOZJukdbY5sO0PSWqdhoVdb5zrBPg0bwHrlZep+AlC269sur+RytZlBEMevz9en
74XFqNyZXAw1Rsr5yPLSFC4qObaPkPQlb+EtGWPwrOvanRdxTVIC1scq5r5cWkn5axKTg3+iS3gz
OLkGDP3LydfxcVito0f317FHlBrskWTde10OHaXFEclqTfXysWQnvyg2g20gjXNKlnu++0mWpCTJ
yQ47I6DZaD+wr6cVV4goA5O08HaOWWSQQjY/XCj/FP1F7cuqqUwinOXL3/C/CRAeHdt8vuq6PRMK
woyX9/wt+yJ7obtcUzxfeg9JjU52SoZkQL7b/2UWauSaa1x8AlLSVikRvqWoP4lDb9GH+BCFylye
sh7k6zv/TVBkMYmMOO6aBEzcK5NcxHk9yZGH2JNZKOWRRZxtnYohjvwf6noWhuskQ/QcZDMxQ+ne
eqwHxaIQR8pc+deuZutqmU2Y7LmF33WzVg61XekNMc79zR6BtCoCAtH8k5ng47No2F91qxM2hOa0
kqpBh9Ubj1QzGsygwYMtUWMgLsDswcNtC9QH6UdiTScnjR240M4JCCYn3ESzwMxFCCgv4zAcCxzH
8vW8Qf2HR7NsVOZYzF3FsZQhDtrj3U554t6j9tEMOSQwZt8N7nBtEEsI8X3mDQqhhYKfGQH/EED1
fAKartbY6rkxz8v8kX/sMlVGXxIiwG9MN1f4vNudUeTEwcebmBUa+DYFOiGNPSjfZOBn1k0iTEoc
AquqWQsOKkhLtaa80jJkX5ST6e29x1b8L0BqK8T7g6NntBOL0IXst+1/qFPcUwq5UqryM8ITnd6s
Ycb3EtzjusIAH60ZASTGchdiabt+ocTZI3fN68gFvbwu/Ep27E1XS3wpz9aeZ2vwkROHjoREL1Rk
i0kXMqHFwWPrsgzY7q9TYOheEt+QTwQmcQHZIq5vxbiDpjZPQwKMqExlWAvaJrxwmwcGpnSK1tBu
jF/R2DRpExFepKAFKkDBCpC9AtKxJwMbY+TT52VzNsYKQcFp0q5h4m9RfrAtRkl3gOe7NjG/VboA
Ka7vhuFzwXiBC4A4H+WB98ctyGcXRlB8eC2W8lTijx8Ka8pj4ihSR3fNxrRy/ubfVSMDoPUyD+BQ
rqggXUWmgTBF0UHLzsyqfUm+BLBI4KQrWPXMF+O4QckP41Lkal9sit9NqJz5jx9BaR4UKK1UAewc
Q3lWKnm7Rt5zSLA4Po9+6p1VVNbtunbKbxyFaj2S78/slX5xp7JbwsFatoIdhkr88QWu+DjEWPiP
l1CY092X5iirrritsGnGUk5ynbDxllN0pn/L4TCXYwMwApf02dL6MgAIUfo2p798va7mQyRXGPeO
fS7vo8HcFsDwT/wgRcklOGsSMUuVsNv12e2eoRJZUekoXKO72fhib1YAvktxaa4EbZP0wwudEJ2g
qGpAfb4O0g3NiXox9kRHJCWf07iHSDw+WelVCwaXcRuAwFvDSxBzBo8HJV+SlfH7dAXnxlCPcN8W
sqzWA+lPXQK/H4OVfKxwYmkT6reSF79lNB94CqTd/0ZorkfcM1gcr/hgIhS4FwHgo1u1snUIHU86
EKisNJE5rrYUeFUkLAeRjt2HBhCCvQ4+bA2/hlI9/dddKuNQ5Xx6TeA2SuMu+cLqq16pATa4Vmz/
iwPw4vVf1lk6bKSOKXxUd6GSfT3+lFsKokXlEsX+nPQml9Ote7SC8rMki41xGf/RnuubAVhvrnHt
gJg0fp8CuIOo4bKTHgzSHwMzQ7yognlJu/++LKonBZ2JBBdmMu8L3fkLOPplARl+kiRZmsr/LOSs
IrnbwageLqwN/b+T5x1/zS/bi0y4ad2LjWwdZkexvOBYd/P8ipwNl2Ho+CCyGVLggzEQe6kr+Mvw
U/UTGXJG6Uas4odAhgV4sl//9ZwC+x+c54ccP5+JJEzGIOjS7wiOW5J/HrIjbArFBHftssxBApg1
pgKtv2gHNJqxIUFsBav90vEvbvQY2IPfAS1AQ596YyB1Mp+DWfHp3lDQ6zCPy71VC/HPl9ObR/UL
hnqNNpDVIXu2GxKvYJq0XW89UixFtNDVpkbFn+kPm5FgGrBKOO1cbtJjkrkJ8r28isd4CdCWzZfl
hT0WE6rlMSNKvuOtXj86v9XKR7rO0/7laDoHRmNZ4xcCeUbzD1+DRzFZqIvh3kxzb8xOwfczcvKT
88+9moeXhp33mMmc1nD7C3MTPDt21/vfMKgEWKw5BCm6ug2lxZ8HKc93/g3NzYwg0uhmQkaM+QpS
sOV/a/shHcLVdf6i4cGKjyyUzKVSELrHJLe12CXBbvbwdwx++VjRwUbZKQxBSvuLvu0Y2s3M3xZC
jm0B1AycrcjB5VqVCCjuAcOfsZC1eEfUhlCdlEAEiGEcAcXL1/OtR6irjxP3eJpaHF3rp+oA1izp
5sKomwZnBcXzIgdaxrHRlJ6XQahjHmbFw6YuHG3LKtxYdJuhkLqqmSc+vnh2mKiFKlrHbRnV+WaO
w55AdHCJHqRRbBaPqlCmc9+9b0BP/g6l3niXdWLXI734q6rilAvLr/Jqpmto0o59OIEYIJblb/2h
Q4sBdKeKy+CyiGYeDZI79tzCagFBbY2R3bHoREjD8qqNx1HRQnT8tJESBts57SBctXIJUFoN96Z5
F07hhQhAuyRFQofONYPIWy/uAGkFoOYnH9nOK1v2hMe5x/o6U+dxg8CC4uwUDQDccoYnv0EDXpIZ
fXROnfqRGmOXjGOi6L1DZv7vZAzAI9wzitWb1qwEVLeLGbkxz4xYFACHx/uhDGeDyXvrc5kdNq+M
JlRlbMJk6NNp3IWzBU1fHxaNuQR24bgQGT8cOBt1XDSN0SYhAqAF/qW7CB88yc9NJyUZiss7g8bi
h8PsWIXZh1emLuFysOy4F9wbwhF3eLCVUJTlM2hYg7qmYmDj8UxoMZ7t+Gt1y+vzIAEgGN4+dgKl
EJEQ6ZrO+ldNKFX8NF3fEvamV7jWUAAfXRIvfdOjQec0kV6l/ieD9bDHpqYJ+DuG9ztGujgTj5WA
Glp+AlNsvtkvkdyJwXKS1kWQSlKeYrhi77DMNFCNmAlB6+meHIm97vvrkzr3v/jiBuVwittvvj8r
wcLWRmviaPDtkY88Go4Gn+EmN7GCPb0vzYib1NAQJTcX0MMvWUrC9ofTtDDIwolZ2W3xjEqm4NFG
lcG35LYWHF/br2CF57B6hfD0599hT2o3XcSdXGsZkkaY3aXeknyNbPYFcUaPw5nKG8CTXDf/jdr/
KyYix9brkkD6S4Nz/Iz9DUwLEOTXcV9NgTFQZ/AejlVc5iMo2R5APeZJnTTECbj+3shVUQpxIRzk
ANOMuu9p+Xr/QvLGrZW4D46dzKWT8Gt1aTvvkqZ/nNxsGSmjfmY6resUWGyus8Akc+N3QdfmF2T6
hnMK3qwGhMK1fYIV7J3QYxbM1A7diZlfbk4awlIjUijHap7PJ++Is/uahPyvEQdSEaY9T/u8nBhn
NNwKX+e5tJV//hIChXw6kUEuMDzW7ruLyRLU8PHMfZM1STjEINg6HzNMmJY5b/UgE/UhSt936NPQ
iUTHqVwLSYrxd3woUV0LsgqOVCwk0G9aVsnAX1vyBCfvY3e7DYlKpHSh1Q4nSIg4bP9YveMrbafc
3iKTbjuV0ufHNTx63Zr2j/tszFe+xy5r1TdRwv0u/Qi/z+bUbRRVO7gVqRHWQ/S96eYOW5DeAddy
7zSRSyglqIWmghaqzu9eVZjQGfvQrU6B0jzDI+BvszZYYfmcdWU4gWdgfhuh5//r+mskQJE2hn6U
+4UyHiQnSllV3hf6RteAO1Vaiq/Mg/AS1cfRytGTxfA3Pew5xa9yvdMCmR5j1HRyhv+17ztEzVgC
oJWvq9y2TihtfF+nF1M+2y9nMwGSReFfNt0jfqa8fIGG9zXpmxZGBdSqMBAhxza7HG21u3ZkOKfS
zbCIZLIad+it+4GXIMEigyb5A3v3v/ftTKS1gIbCi/PGP6ivUdzV7fQXP4GVIyTYtYHsvKX6pLSZ
QFlBCtJf+uBACMdMGEE7IZGBGKSSRwrlegSp1/+mIeFt20I5UY9PHageEL861URin368PbTmg9dM
1ayXzOJbZjxWgammKFYFfPFWWMOza9lJKCHzVmtgY5fu/+GfDP9Yl8R0mVtQ6wUJXYAVVpIne+eT
bXIm1t4ajfVKk5gVQqpEa5BhRtRxgzcFFH0lfLPWainOcSHekGyOrWyy2w8lEyTqhpKXVIieCeAz
27PPA7R6jHC28XXg7v6odY7PL+mI1v3OnJOLmCoIrpe7g1p3iIflcpFxJ0ovOPr7QVKuYv4gzldP
Wu52UhdIhTQnhb3fHoeupbnV8RQYGYjy/FQYLQVe/NQ8PL6mkOJszFKrLi84e2J/W00NomjkDbhg
lEVHchClO5I0kY9SykQgph2te5y8raUUJ+uRZ9nUYJkcY6GusboDjPsW/BVyT5riaBW0NqpBZKNs
14+rNiGo+OE2yYY/WFFpEE5ybaISQzTexuwvO/IMe6CsBzWYkUAhuusYN5Zot1igpYVs/ti1ZkEg
ayy2N9Q0X/MASxjsCyhyJa7qIHRRTBTnjtZPQVgadpMzmXIuvmAfSaUmRoaa/+zLBn3k6cNQ5dxM
0pnI097cekFuDSyYeNgwaBWzz1yV9vW6aSquL/dG405pp18bGBoj+XW9FBcY/TSyUVdOvWEMB6JN
6zZjxYhzb6yoqp0Kn8qFK4EkHuiFs6B5swurie3iPwhHPj9Jh3wpv6fWj27fmUbEL8MqzW4CchT7
bUgnatqCGdh97Fji/oHEAuK4ZcjDcSTYHi33U/leCopDg23c2EV67usU1tl7bNqzJvBBPMEx05py
YgURnMXrxU3gaEdXVIuUjjQuRlHFT6B3S6p/nQDtmomnJQQhejmvMWEZ7HibqiQOEASxol+9vj61
glsSdwg33pAKx0NLbPRGCCPI7TICI2hpuCbLMRf++VIxKdn50p/+3TJSp/RbSZEuCxQFaSgmJ8cl
dp1x1Jd9Qespm6RvzgzU035vafwgQsxgl2G+WfdKvRc3LZ3X3DYPYQCuvloulNFUMRyBD6eMAGUd
WJ/gyK0+odUQYVjgR/H4/XfFTjIRt0XWnQqCrTrBBT08CmBSe/Ld0g8+BKFKit+d/+7zLIioLhJa
ZYfJqgurNoadfrhha0J6qfepBnyB6334tYEcq3NQCglxVe7AEQxg4gMhFNudsWDRXwU9bQG63E2W
ZwfqT9q8ZcA4LMEguorzDe+wYLmTwAEdyhiBpbAmFJleJs3JCsCqkvdXRUnLVJVxiP67cj+DmQHb
eukssBqP0B9lgK+Fln/1/otKgPfWYV+nfU2tGhSesgEBj3FS8cNMge+A/mglwy7BIq/A/7qOtgNM
cb++psqzJyqQ2iyJvVJLovstzNBwQM/ox9QHnVr7exKjaNPQbtq1Yj7CJ/dFiI01RC22NjumdXZn
UBq8vtqkLLZ8zWUa0zF+2vFifAw1bqAIYiLX6289fBxTeWNK4zSfNJ9xrEVic8tZ3cDpwhwhHJeP
Sww3Ga73vRA5MvsdjZRNI+fjXhm/3E6dI8c/RQPK6FJ/UKArd2Kld9LaGzZwD3pN0xJFaEi/CtfE
ebhtUZ4QregiLt5oC++t4ZkKDne5qavm8NlcO/EvriLosOCgIXxbhfHbPuVJyJgvyLKDAW28h9JC
HgmXwrNVuZf5P6VlSl6gbHNY2J8uGsELvHrWh4Xa/EH03B/sBGvkuWX4VPyVQphxkHPHsGbP9iE9
ezh3ME3J6rttW2xqi3G1TdpT+Nwf5f7vrpFYya7WTFxR+PcjpseenXWUj/Vx8jDX6CkaQtxo9fOW
2SmtoU+Z0W5aKsNldgmCREoruN6vC+zwqAJbc1/878svvMGmshi7oAV3ljzP0v+Niok14CGxKyvs
7on06+UHKU0TBdpXAMWUn9dzohK+hSVEwwQYZLrZs8h7bs0IIkhnnmmDyjJzDyt5sdCwwgsGnWvM
zzWGcjaY/Uj/ZV2dJdi9vFB3eqcnG4ualEw7N4qtHjwEDXFUZnfHLmsm6VuqDgW0/YjJ4PWlPkMl
kb2y9tWa0xx/JQ+uZ0u/kXc9tHzarhJxO5Qwf/jOtnldJZMBJUlTHLoo8HXh0E1D6UkO0D5K4ab6
EFAUDNcLtJVgFRX7yJeTLLWe6pip/90lUvK2jR2xkDQYakCUBmTJDbEolWyhscDOoAgqFPUcxyNg
hGVjODMQ2dILTl1/5PChSrVSAlFupxHKPHYKSRAE1BATPeYK3P2N1jXToddipR7/UDvW7NYBLm5l
DtLcboiGjnl/g7hUgaqJ6pO4jTuj7JTrTsMFK2BgEm6KyOhiuFc7dPfbGl323g/aChk8acGbBjt5
5RuziujFvzTDdH0qnrXyVFh8DSNO2ohBhtLo5fhNoa5RtIvORfR3koiFkI2OiRHzbq11r47gVcXD
mEdsNa/ApQX5DPNhwv2c3VkiKzNUmmayUGw4yufl54pE9AU+xBaFijKqigcDMwVlP6WrVSg/Z5gH
Bqd73IxQTT2anG5Vv0xdbcfMB4f+cnV8zF7h7OzEVr+gxIvdTE9EitWUoq0oyfOTyk4B53qNBeG4
jPTUKy4RxyZIOBXQ2cYn0+GkQCCBdDLqCYkQMeQWoG37enqf80yBW8kF18TtwIRLF59GRY1JyX+8
Z0PWVa+bHVk8wyxmJ0buE3F8eCeJ0mlWmbij7eYOcBRZwNCL0hSE/6T51WtGGzXs4bqqIV41p7+q
AM8N8bQPJ+cv5zqk9CBx/+7khTAV1Rxd7rRj0ZucSwlHYy2fTQk7bQeb1bhFYClGB+STxlSCyoTY
/AcXEFyvwceQDU0eu67uRP0SBwb3/IrySTF2mZD134j60AX0C+mVd2OZmCk1Hd8kQqXgbh9pHFEz
tT0wIi4CvFIibW7B1GNUycpvqI98OMDKOWdgqArzA/omR6axb1jMM9jye4TBKGK38RHakPflOF8r
gmy8vcUM0dHuCZ1T5MTm64M50YmtxiVVxtqRxDE1T28kIba6thRXS/rGNEaCZTfqOiG4LyU3O3zp
lvQd81YDoi+nzy92QXIkWg6A/zBrhtyPde6bSWy7NOYlDuMV+Odn5ooB/Pg0kvZXO1lH7zznJd7X
Ii1n+78DSuTTcsVL/Xsp1YAWgyFk6WGcGZERN4g8wqH/Grp0pmL6UV41PBQHRXcPeSLBFUgyJUmf
R3gbbSUVRGju+TPjRTuYO1LsaYlaT7Z8q7d1Wv6HPHSJFrWwKV9g+AH5HxvDsngZiUNtkYMoaRSf
YV7CuBmDa6q9Yab50oRJULFv19A150O12PchB4Cd3XhbgJI5HQSMJjvphHmMLriFAWweYiju6xEE
b8j2fE/0eBfFHSLFQsp6rc3Tc8iIrp9f6Ga6+IR14Ixm9LLgRSU8xq03F8IWlh0PaQRTlOJsZrru
/PKQqKF1Y/zl2YommHJ3JGNlpSiQOxRsLFzMiljBSHSa1t9TP1nel0dV0LfPwiuzAx55WLMzfhtv
EscxjQj/CA0diXsVH1oo2c9ox2aA4GcgC54Zck/+RS/rzdUl9+f75xUX4Jnzh330uBdoE79W0WMo
+e/x3yWcSKf7+oGb6/yXz1cRT7qrZ5pxVsBLrHVQuOuo3OOk/BvWHAP4pCFA1D6+57gh428y5XUd
Ogk+t+YnNMVH7Ad9qCpZRxXrYwo0Q1pV31BCoSm+yCAkwiPJ88Koi5cNp/kdRHSdEck2Wubg828M
pCvOXCz1LDDTl42iIkeNvjOkJsQtxxgipVHvtrvX9tAC0368N3r/mV0cz2tsGL/S5vehjz4NWB6S
bYSYzNMt3VdpTUQlNPkLVSlPd1TBwNkifPKPObNse2txwIDAX8CWeOOmrw3ZTThSX5bXVsbA/dml
gV3betnFeZ7wQAb+E6VQeR4tMx+4WeutZbyo8J7y0Pr/3q3teArd0Mk/INXZZaDKhrEJq4syMxXf
5J8/6g7bHIT2PjszxKJgqpUmRkK4zeYgyx1vY6g5mVxpmhbY/EOoILQaZE9yXk9+2cP/2seEJSn6
u1FR48upS6EzpQ5HUgOXxgVFlvuUGy+sKRm3mTHsmEmvm/UfVYRpdMvM8w4slqXuJsjlgsshs+Jc
A765IEOaK1vv4rFYHOK5zGC3+/RYDW3Wm8q4VFGV4qUUh8G09oPiY8cj6iECASWFx1dIWYNnadXz
azFkzyu7Eekz1HaVG5T4EfvskGNHxy6orqSUktY9gDs9CR21YZfpqUU7AulW3L6PHk0JD58ZoAWL
Npju2+FAuzEAkqkWGFL/JWkekFTkMGIcZ26+Xr7eU7n8kGkXwW94aN8V9CWYWCRMYNM96QbW/BBu
k4MA35Q0yi+DPdtMzJa7V2Yud3/VO06iuLzDSR88oVeI+dUFc8PhYKFKnu050hKXYgjdZJHAfzIv
oPh1VOFBuA+AAbFG7q35VmEsyOUIg94SxNHDxUeaf1J4ac4C0sZ8e+LkCUYgUp8J4EsO8TMr9cbL
ZjJJNQYpBroNSwmJc1yZO5hjKOhxcN6z7WvkFALhYOj3Ydtsp4wectklYunpW7CsjMsVBtyITZSe
UQ2iWqJ85GIVdkABRInyGkptRiltQHEaYDMdhiuk+d/4VNBp4X00+gLAC+q4hjKmHslwmzNeguWQ
fWBfGlifLywhc1ETbveO7DTcK+28CobPDWsIG8/JWx+PLSLB6VMzEo+zYIZ9DvGzhHCsj6cRTExz
Wipa9AiFF0ziuppmYY5BIeYn8xBYni//8jgBvotoErbzGZ7wc5PwmVQsPRRQ/0eCLY2Fl1Po3fCI
UlibEaexvUVTXTx2AdCXbRhSkbx3A3B88h2f2c/GKs6r4YOSNx3tiKWCZS6qGp6i8MPIcXx9C9s6
iKnm2vdyKsBZZsHpMeZzuizMX3cThrWaYxlEELHFr9UhtwgwbmW/8/t4tl/bZ8r4rFFA8p25Uuma
Grtfo0uiKmw0siETudW8priySJQ27RG1cVZnmJCV96pHoxmqpJ4vSbXF2V+CkpUDdjAowoMu2BJs
PMQ0FLjMbhIHKgFPfBGdDr1Wx5DxbQ4c70FTtnS6GsYbm+yGSNE2nZlWdTtFz8k3Hl8sTrH7sw55
2tQBeqlchiANAPmeCX1PPxj8E9vpfBFq8EmDBI9iAzIImHjfS/8Hw3xdPgVLItagGIU7qy7Ij1Va
O5IY/vWXAvbClfrRK71O8VkogDfRG7q0cBT4PRCm2Tk+anZ3epKrGgvuI2VUbYmjZXCWkSoHa2Nr
mcmidLil+aqAtGNlmltx52JjyoHkULSHkhZJ9FmdBpRBDvwjX2n/S2o25m2GaZ3ouuTWtgWCaMEy
TB0Ug50eMoEF3/0jbYjcUFzPdo+xkAjqtQYl1Si8BAa9wArXypxi+MXas5zq8P3b5SUz3sk54hGP
3uNwhuS8MzKuFzENsA68IYvRYgcJPFmpvx4Wjn0NWxKqXGE3ObYPTKNJ44GxvuNeEHul9j1jDo13
w8ZpBTb5fNO0ryRFB46Y/7pwnglQoMMpmptHqUQTz26RI55QU1HWvqouaYDIGe6BX5hpKUXfaehn
Ky+Y2abIaca4gCqOlzfGS28/83pFZKyCtnyfq120A0WensPzBCYPnWHNEtQiIT6xe8bTUttaUn6G
ruPxKjZzj+Zfar+SqysqA/aaF+znTLfM2bSxfGAnag0MT9HjE34oAELqLzJthoqwuzZ+ujt6h+IY
kYSsCtLcRKMagAX82pgJLYOfSIEanjmBTLeMxHj/1eoATcjXzojBBozX6SZrCWU5ktf1WeSMyDCy
rVhHYbHwYgTp4+TU/upHtfnHkcaa7iQQHyGg5bKYID2fYJShpiDTO2gdg3LARGT5LsH+cmJuOa7K
mWZ7p8rW7s288tMjOSGcKjnTEeS0NpgUt8jPnqURFqhbeN5+zQFHh7mFq24us8px08euHD0BL8+P
+VEXJ6OumnUukv0s2/afwOlvBBCpcosWn5Tl2avpnlrSeDM53uc03fo6O0U/qiBhN/mbVB2gr+/V
TRQoyNRA6NDUZDpwNuWlyRbCgfxIlW59/jWgq4ayaKhYUc7IMy7GrhJhFhGPm7RyL1hyp17Uh6jC
Qnf/g6fTS1aqtun9C7le3PeYCPpqWirzZOF19VTz6Ph0Apm16MVsitOE+fXyfw0pTVwKltPnjpec
46JnaXv9LRwVRp9nLRtad5G9rHdRLwLaESxgAxz/aOIVkr9pCTwNGF6my5cfYRu0q7sv1YvR84Zn
4Dmx3DeLQ93yVvDzGoucQITV8CGwbae+4uV8Plfl+UhkNsmU4E95R6nJB+HY1iuyrAYr70Vr0YTc
LnDUt9HbFSu17ZD8UkpyV/xusVRNXoIqvaJ6L7Y0+fU8kDMKAOj6wD1K3OQOkCQpIvC7AvFUNExu
w85GyDnhezRqqrzBtJgUQMfTOmgHUpLfLXvZ0dH+uEJTKZP/sKjOxuh5d57okWsPd+sDSHqdm8Ox
H3un1EXWr8w+j0KqbFBDsJlS0lzLB7mfTThzQ/+Uqdv0k62X2QAeLKgv2/6rKneoZqPqv+KJc/6d
dwDcN4MGDhWjKVsTgHSTJQWG0N2ymAvl3rlvbIRIcraDfUyZSvPSA13TUE56CkjMhhg9zY1WzPeM
k2c7mGjQ114IbXh/sBtxDlylb7x07V7xghNrTSmx8SyfHygQy6nHmkH0EksiU9aHYR+SPKfZeB9W
fnTMFmmBcqTdrHZWRA8h2/RGANfXquioe3x5b8zHwEY0W19ISbxlAOlzUBAqwEqRiqutprYLy6Xp
OhhJt/pGh4TSJiEMC9meyT7/ahWszBsGDNezzHJvqJGPscTancQlcywsPTdlKTInKHEZXoY5+deM
sF49dZ/XkzafHxRbYa/eCz4Lr0uqO2JFn126XDFXMBpc+yKBr1w6bzfZ4x5TjE+JAN0Vs3Ltnr0d
zDqBXJpCXzykUbKRKjN8zGpBG6G2Qw7cjgcA+BpT6MN2i0NIv0CXl/x0BdUvH8dIFPuLiGLbUC86
plTCgmqS3ER0bePBszjgVgocu5M8/Tb3SUohtp5bfmiGWBmp10BUSd1gARUgIJ36AQJV0QRPdbbe
0s3ROmangxJeZGYjAWVusuNBA7PnV8PwCkUuGDlaU2vWM7cKCSMGOvgZKa18UpCPNhXchRKOuYW/
kMSFqs8FqhXifXryPvdaDOxzsmPHokhWSpYCp0RPPNh0V3NoyOqsFIkcow8Bz+4k6oOUAXDODmpo
DPY3Cg9qbhFufga5lhzb4VhD1zko6M3Lmp+rehpRm1TbRLRklHp4HS2zG3v1Y/FqvPCN/yzzWoNP
UzATtL5ItxaE//6X7Q4oq/0EiTxVLeLXW7iJujpL8Z6VXcLTO8qymsC6HHAltnTfATjbp8BQ13+s
lP2wCaEtL5Aa2MDxqLFRwzpki7a0BcmcPe5O+zL9/AZO6eWl17ErJ5N4lJlGIIJbMa/FvjcIL6b1
zU8ukVtSWwQO6carTu3uAMhNr2X/vUfi8iexQbTFJpZ1vmyK/vWfLrWBoRbsixiJ0/IW7JQVIGH4
opAtQJi3NbLiKjvAPBmJv5zxRhmeEUHTRwUeIuSFqEOfOSlTaPocUB81CHriLFw3cbo6lyfNxklD
Lfnb3xl3elaVrHfgtT6ai55buDbyplgo6v8oo89ptQLfX/riWHG8maRdqltKrIUc2yTzT5rUq0Rh
u9jUvy4aJrr/HvZ+SLCmXTpuhf+0Gd+iiI2szuOnjCi8zWIsvB388ILpw3LO03FpJbNNsZ4rQa6j
Xxf+HriI10TiKZ6UaT9HZ3l3cI/qrdr7hSN+6yHYiftUb1C34Z51mR71fDvOVrgVv8B46PX4pDjx
GT2nUFuWgYwpAH9yE+FBx3umhB6DsX827GiDt8IXTtjeVgSSGFoJITW+zKqjQJbrXM1lhnQJZs3k
3YUHk4plcY++ZkBKLgJZ9s0E0YA4bHnAmsueeQ83FS7a61ASn78mI6Q5eIpc9Rwtp61wexwVK749
kawEbOiFIGVZsZS+PYibxp8Q/CABnFkv1vkb2BbbzilooWZJdxUiBRBkXDvVZnA/CfzLaV70GLLM
rnX3kFPVXp7ZIqzFGHE0fhsA1FsTj4bZuiHY4MqpDkujrEOFwjgMpa2l7/UrDK4tbGjttymCbBcP
fyBKkFjNMf7kTWk5l5R+5eNl7vY41gtB5LLwE//69SVbb90MIRa7KKGFtV8/Gig4GDez/J8kr3sC
qB1ao31Ne2mthbkmPBUPnXp0/oVC6vYmHzl+Kxssg2pRD3NzmqNVcuFerElU54otWrS+zDz+2boe
dkSMNlLxsbnIlOTCaaN0x054bqUWkCBIzho2BdxGy+QOf6NQSIvaCLdWE+w3MnKKfyTp4RaTdzUa
bWhd8i2EqmaVGIR1vNNPuu7tHdr08S41nnnI08iJkUBSlBG3QN6aqBbpUO0J2uUhlwh4UFdEBnjx
y7x2R/VWMGGDx72rwKN8ukjrqIeuG4fLs8AdZ6wiOUiKRnJUmvyMHebbE9yqApwf/v2pJQIux/Cs
ApNMKg3vx4UZNV5FtyjPSibDvpeeJD1I3l7x7PA5rZLusKr2we21Yduh9U0lbMXX1KupQO1dcR5C
L+ksiupf21hBGIdat97B+hMMW6xX7E1UHocPzKVteYo6Bm+KN+l3qjWyB4wt+M6Wnwo3CB+pzo4O
MTOiWFuB9QQyZjAN+5kt2SNVYIqJhxbWuRR2oC3YmuR1kheJX6qjXBwK8/sozeYQqxNukKFfFxU2
iFhu80fBk/XORNHx4w7zBxLaptEohbrt3qL8fUkCQ4KH4PzOtr1SNph7QQHYkSD/baDrTewY/Wag
crxFSaQFLJf9pbVjRH3YAVBYG9HMYAiXnVILw86hSVnNOJILtxALr43E04XU+shJ8RAmgaKHv12t
6mdCe+G9CkN31uOBYij14TxRM/3GK6elNzr7+saao915ZOCuc3pmtEHM6uQY927zhxdnGHeMh/Wu
k5foes39g3JUGdYsRltj/L+FIBWJKPVB9PRou3Tw9iy3SQn9/wA+GbB187SGeDO4nbzTB60L1edZ
Q5AGMy8rT6Ad0gf045mGTGdOcRwyy4Qq717uLPVwBCSYOWARzt9k7BF8UggDLlcdyOEejs0mTxCt
CYCQZdPQ8wHqYi3m4Nn3zFKVWaHqWCLFyiz53zDHWvcF5J3Ma5Xw263aXvMrsf3Rco/vcT43WIGA
ufVLHMILhmKEJY7mpABlnOq9AAqvmprXB3tJsumqVG1MojRjglX9XfWsWEnFnf0nCqWF0NHe2it7
uE+h+LsALoJYSbDkHW2IEBCnRJhecpd/ZPE3inI7MDwLJ/2HSJYZb7uD1260QBwCYdegMIJohgzP
V+LPUVdO7Mc0h+BnHiuGRqdqkihLjG4APavYQfoiEbYkBxDoBBPzmdx7KWzQCakRjDm85PtHbnEi
NwBbx5+wEdzArNoubMTw1Ev0Y6OKQqMY9tITgwk+zleJ5pGR6dEAnc9+F0SslKBYpJ/URYaUN7+k
LOPVvzPo1wVnwBdy70FuOUSEB00IEHn577v/JMhGX/scNtGstrox+FHIWyHOXrrjRPbnBnYVUEWs
/W0sg8rFUs71zdx7uXHYCvQBuefCWZsItFMd9Cc3kiNNDksZL1gkSgfRsKkMkg2+dCv3lNESQZ07
nZ2unY44ZSdH6bJWhP5FjPuCmHQCgJDUV/Jqt/udRxpxyGywlv3aq11RPte7BJt6kZ5ATktTjpxt
74/ksUbwH8O/+gVgcSlWB1sb57QYRYJS5VgYVr5Ls4PUnZn+emOhlje66oqq/ob0xIVsi4fsag0L
w89SXkhGSYpg3QjiWJ+lkhzkJYYok/ORBkNvQ8DMYUaUSLVcuD5Uu9xBYcDyKH6OLEwpzLMkCaO7
DcSx8j9RnvOvPJcvFHTsR9g5LpbqrxKZKYBXb1+RSFfd9+obARe4AONlIT7onrIHVzWXig9Kg1n8
23wveqJYIYtQtOmoZFkYNmxn8KogTEyexGmrZkqs/r507o6vKR+K9FNB6qqfdZMWbjUsKAmQtHeJ
UhCyMqFhrOAmrcMVxibMvVP7JZRdsYqB0GlAX/E0nSTEebuAUXeQFUU0SAlUDO4kmJSxrDhKIp/+
XPgHbm4kpuDKD4tmjZznWMZndCkhIn7IVl9FT96ArQlMyVAwaKtVeJ5mqRLlwLt5IWlnuFBJ7A4r
0U1X7UfEDfZVfXzRHbUshZUCEJF8bG7YOnsGHgWwyiDQ7ATdpXrl34N2PJXCB902uRolQ/eGzSc4
ZirOM95UEISP1fUXRaTn3FdOdc7zbDq3h4+WCfyz8kxPPPLZZehJa4blsLJmiEiVvHoCsMQZntAq
V0Q4eTNTGWcnGqfhAhLGnyppYyiiCTWRsQgyv/FoyWug5U7y9CnNw9JgvB2RhWuLHobSGVJhGQA8
OV8vrXXaZGB9pf9RsN0utjS0CRvtor2hYQtxqIXF0jbChv1RiFSxFdcdeZnT0qZNjX5HufR/1jtb
w5pS6lWbinmH9ANe7JZmwLXeHQL9DMG+HVuROmE2g9TEpQRMIt7fapqjwyW8kPUHvLcA26bzA/Xe
FCVOUvV0I/aQSbNclIM+Ldliugv3YePqreqgQ9J5u2izX5GlDAUOJvRvj/3ZmMR7UfNjs4bSKAe1
A+4XfUDggWBrGPO3mKd92BU81NaO1JqPUzNXp0J0X3NSdrAS8SJEDkImcg12dRVB+YGnNJVN6N9I
z5v9Pd/1XCacQRroW4394qZ1kARi6Dl2TN+yuVP0tHhCeMLwPUsfUZ5oEz6MmEqWNX/yUdt3kOCi
5Xiagy3WYfkLQ+ZOqaAdKFllrkmiHimOzO24aUegSV9/fYS/9ssfhmmgg/T4BAkJhr3Hzb86JTn7
Vyx0UOWZ50pB4hBzBeIXOOyqiQhPQhYkWDhfcjgClWXl/ZcqiH6D6GSuRj7GAQBDlQN+yK8zvEJ1
FLJX/NLTvBSqd7Xp9hMAzNnX7+FEZK32FJhpQC2ZCWhcxUKsbA+kWoU6wjslFLtj3NIEzpeAb4yX
DxcUrSJIQnMXFyiurKELNQxjAsXnnQ56X0jpE9d/1oOzok535DnGB5qvTN69O4J8PZub9wS0GPsZ
haRdqZN1scbK5R4xbfwOZ/5z+HMqAxknyx2C4gmKACNKjv4qHDJ+tx65v5Ogb0GWSPPaqYz2Lv+p
POyaURsUlk9Z0jl6+GT1cGc/+tJ11AqDM3uTBTf8gvCtFNpiZAgXT8+z5MsoEGN70OGnZUYD9nlR
nG0gtYcLGYsWk2klg845TQQDKpPL1RCjHriMp6gY4IpW64S7SBd8Q/0F6YePFh1Yh0+bpydkEVuH
Zt6Epc+wWhFbzTHlvJ0OEk7uvPAG2cjdl7dRogjfNwEb5l7yLc9A67m72WdXW/rJGTCOv9ZbFjQB
yWCR29BNBhFagJVZDaEsei7IpOhvDcB8aJeLZm4F17qnWLPddP9i18m6NGHxoa4eNb+5JYsBZDIW
8o7yxb4fpbsfECbB1poyOH/4H7UyGz7dJig8UDqF2A+3YMbguhYR/tBxfEfzI9T3hRIzJ2E+Qweu
bXMskV5BmfI8xT4pzEIO3fCaxoqkemo1frEh3BbB+bCIM8dKLzv8ZBbA7sHWfwYQMPhDBLksijQV
zWoD0CvS4kpZPz1/A6aZpjO80f3bdgCwa/zgCJvgg0NCBGzM51yPqNZsdRsoi19LQXV58mrunshN
Uwm5ppXGG9ZkdZWxSnyEbIKHoskQAOzCRfARqF/6BLruqPCOk0GzcViRgah2sAy3idIWa/xxS+TR
f7zQLi/9fhMwIJvebLkV1yF+gCDCUvr6tqp1Ml7Sso2bgOR6VWvn0ArZuy+S3qoFj0BXbRxEcbnd
87sIfDhbNozyI5oQrBIuJJi0v26jmh/guB1VigKuASZfp1AnzuL7gZwn0Fyflpq56XB5uQtrbHcE
it/IXnepT7g9AdtT81Zu2gij+9+lHfq+iJXxy07rdgQBhicZG09o5059nL7KErvmGvwbXHn8lwQW
RZljLPkB3/hc952l9bLWDyD6eCp7ArmBZApS5molTnuLzM/yBuLGMaVQNaju1594NLTsx5gASlDk
eSS2KVtn/WtpLX/+PRdRv/UdFDW/ltLCW+vm09/bCwVlEIJAi/YzTFuKPKPCD+yr1KDY40SanXNR
yIfLOzkieeTkt02V1fn76yMiSPryHgIvNlzqhnTBbLroZYrXF+GpVLFaNXKVmWcrWcKTyGZz3RuA
5k0VtdS+BgjackQ9fthyAZA0nzqWsUHa+l7/aPUBYsVYcOInHCKHAoETDMYLGk5bbc0JTOJrZCFG
5T3Dbc9w76qTZDJDtbiEWNFMw2RQ68NggvoTG0qRbB3+mfTeLyV7PtTClu0z68CQjyylyJmH5BFw
Vd2IU29CW/XHcLovPj8aqefxNft2jIAVOyMQiZTCKoX9cvaMqpwiKickpQJDdvDAEOjP6fUsBh5U
SkrDqP38cyQx9uVBzK0ziackqvOWdbKRTZtcI/um83NUhGfvzDrUDmGyuc0Hd0pZuCQIPf6Y2u3U
18PfQqkVLCZ2ddmg8kXSdWJSfQNPc+vo5kI7NptfNRlxZslIW8o5paJL76s87Jv8RtFFcNj4y1QV
aGimxhJY5YVFLgagIQxXW1ivxqMTJHomQAEnOidJcq2PaLRx8DJcCsMjM7OlkSfLLFQW02eNxwsF
JLbot3EYCbdsQ8Xa7JMSPUS4KRcMqtpoKfq+BarEX5jvWxiFOL2Rna+VnFu/3mHJnK97rtDR+2mU
lHtlJOktFj1rR9/pdWzBxxuGQ18r0OPIP4pV+ivleGxsyDuaviZAb4qdo6q5HCuTAj+i/oSLZLJZ
mNf+3RYtZ1ZKK2/vvaimvWJoh6RmZLmxaI8+EsaYUxbBVwvw+nRfjWPXBjmy/wwjjWJWDuEzfsD4
eackkffIgsiLnTUVdejFTFSvAwVazhtwQ0/hM3OvouJQidVBDy0njj3mdG8z8tryH3lEb4tJ9+KH
ieicJeL+K+0jbZcj4RfCDKfJyJoVn1ySmGqVJspajgNBCqWUIljwf1Qq9MZVyVL3quJmmXAWuOiP
aSk/q8C7GaLS4Qh8jn8Y1800h3QwuXoqdASJubMPrzgEyF1MBNuDQJBqbQyv8nmpYMalj6nE0C6v
2T9ewBXRHZiy1AoBlcvQEyumcloZ1kzYpPkwk6frJhHZyZdlqJKXc2d6mbWHhfamVwzxERYqVY2S
oSJsxg3zpIY1uwitpXPwTpKYtPKeUKgf1xfVPlww1sPtZiwT13mUuePD3wVXTulueWuS75inNApM
fUiIOd4gvLw0Ro+94IoN+4qIUmrI5LsPhdmlSd5KaPm7NroaQfGc7On/i/YzfLRcBCc2jbPafA3Q
SghcBU5RBH9jgaxMtRUe5kbjP6npcX/SIJYbrfjiQFtwrqcl377VGpSh8cPY0OxxPlPhrlilZqrf
6XaVvgwqc0PqkfBi8jMigohnCMFLdymz3ngMx9BLQeota+SjfN8TETqHanslSHLoBONaT0S4l8DT
ovyjqV8sZW2ltQyaYU7rQsGRbMxxTzi2xktgPdmeOPvuP9j04QgImWDpGgJMvCE5cbtCRc/UvUx6
54iG9S5+d3CtL/MnQ7vVxLm2uiKh1qsthv70OHqmKmrFOEruS5QoaTDXRaC8uVWXo8t60bOHoQrX
3jJr3eeOlLGVjNcmOCkn4LZk/NzkCXWCYWY8/G+I4iv7MDsdZbHitmhHMeLQI+zjcbE4f0Fa146K
OSu9C5gUUewtBMyiiEhrMm44x14detkvUc9FHnN2K6DfDmTYtntmeLbBJyolGcD8ol6lY5Yrn6ow
ocCKuTTSMB33gNGfxSJKUnkk6uVuSsm/8QY2DitNKWEEZmk4RjCYookvFIgwV2V7nkjjxHiK2Rik
CxnXhs+5GJmOdIksq/g2Ym4/fH27BEMlgiyyEqCfu/FVpp/+D6StI1S0nSdBH84bQlHJMePE7wMJ
LN5Lf0jus2j1zVAM6CCbCvqagEa4EuyHV+qjdLqkHmU8ktihBErxEfUFurWE6sJSA3tIqtUXKszW
CyDZ6sygXMzBGOQuMF3ou1VxtEmewGGrCkn9Y56d7qTGvEBjJkmkUzI+UdCSAanzbDV9RStl+17E
90+AjUyyhCCvb6ES3bO+cmIJiLBPkZQqVYTB82iwEOx+ItmQ428mUKhPbX3f2hycvqfPC5ZQ1gGZ
He9o/aBk5Xt76jwYUJ3nkZegHwWsCx7ic1vMLtGI6dUcDX4zwqZCioRf7Ha9EX5+6zabqITEDvuO
yBkvZibz6N9rCuOIByS4xYqVkpcHeVdAxevclVdnC0pv86I0KxuIjUtOXCmHY/jFilPwnhdlU7HI
6TQK6LybAW42oUGcSsoOpdBiEPKIpDzkx7N6jj1PnvL/PE5SlreveNm+HoYrHQdfs6NYzenSF0aj
ph5CxQfi/zRfBImbU5pwesGmgS5By09ilzM5DYM3FM61LYh8lXQJLRtEbk/Zm9Dw5rH6Xr1hT5r8
q8/1P/PN+U/zVD2kLLrWCdestUEUBeTWWoSBRIQs2jwS43UnB3OdwoFQ7j8l+FEupMCdV08mDWuA
LY2FtGi/IRCxWJVpPRlUpw2pWSSV6nV/iw28zwxxvw0+SThd+hWYl1ZwxvXT1DioOTlqAoq87AuR
pAcyEOxgqGngAQTCbtQNjL9hUsPST6fDhIb8/kQp5qXUxw3KHQ9xeHnUnF4odEv9i4G3a+g8Bgoo
ql9FOYSwJVWkWYtbmf7Y7N0tckM6pA2lazLlybj4CBdABcZ4gptOEWbNpRxWKUudD8eNbmZfD/lj
9/H8Y2RN/Zf0XjxHKpIxmR9j3LXhYBJMhYVP80KSAG8CujYJZ8qyZXe4mUrHzRRQwMK2wsJ4sWL9
MK7azyOuDqPe4O66HkPxoFCRVcRHOMmjer/MSFoeH78vS75DKqi0sDR4+F7+E1+2xo1R2dmMfhcA
T0nKv7RcgHXv36Qf0gI0zaBQLJFrin7N5izBh0niquH4DmTFl++8aYeGQRYSI4jwWaCpgGWN54ff
Cp0LaHOIfJUwlNxsBHWg88c3Z75hwbdtQDT3dWPbgBM305E1ooQnkOE3mQZJz2e4X1ux38w5At3g
AXzCrHA52QE73cQiyHiBVZZcxRi3MMsnIwbh4AQGBPGmf1dYBpjgmaynKGdpyQU3o1MCue0KYQQs
V1u4g2i+Dp0KsdlV6x5XAx+Snzn/awIbRjLl4sDb10qfzYZwklaDzF1vtG2OnMRZL+uCAX9cW2Zs
MUlNsEC9z9lTf9KdTip+FQUoMi5T235/klh9DbQHDkUibRoccvrOad0mweY/Jpf1eEhshXBLi6ya
OoUE1dc9KLdviGMrVrmPb3CaNuZGTuKGVJWGA6P1mU5vt5wwwpSphfY+EC1mg+iMW4R1fB2Irwvf
c7QGselcPPDBcqz425snsHdP1JdtVJSO99jaTYM0yBAFIr4YnaDeqxjVxMln4gclpjVoITA+QiJ/
4+fMyDa+ntrKR+j3RSaAWowjog33ExNR3Cy2fAJU90DjMicmBKI3adFlutuw6EZO3XwfhbI76Ek5
03ABkBjD/4KNEJAxHNeJqAXunsQNp7R3Xpi5ptMDe19lvMVJvWVXZTyi9oHU4fqd6sizeh59vqJ8
BmBuueVNBcPn1YBF5uHcbHqJcLwvwTZgVKYqW+6d1P9DqYav79gYp96Ua/WgEM+Fx/XlM50HGZYJ
SkR2aXorWjJ1j9P+g5rjTkwcTRzC/dhpnBXznNMxq2HrTX1b36VwtekbQGEPhEjIYsJmL/nR79dL
3WhTe/o7j/5QoH937ZBc1nTzgCFVCBl+xSebYPGAyFLglL2laEv3YS74ZIglPcrnF0oTR+iDPtbT
s32eTm/iOWjzxiTbCUso2CVuYwNkLHoi6Z26J4vnR4Vj5jfFCgw9u0kj1sXXfXwZNucY3g932b+q
8+x93+rlkz+F0rFXQwuZ1jPtiFCt8M3O2YaBTNYV2UyazN1UCooN2akofk0hPihrnKZrJaPrwDSq
W7TrwhoiIH13mRFj/YlFl+THn1sM9vNVbDvO+xfkZWJlh6rhMAyTTb4205HlnQ+HL7DF+fmwiXpf
M1pZtlClTeyUj3yDleo2GBxt9TMIluAKQU/ISIjV3RgyAiN4KUXWz8LcVt7B6iQfFzrgkJCq0nr2
2H1eUYnDXgOAiRrclvgo9k5nHyeGOGwceQgMjUCLt5/F1k/pN2g7v925k/05zlhXkkOwYEnGp/Fs
8gRg3u2w3u2pARcOjhOnbGRMIOoLX65ntDQv81yDkU85veRHAo6qOa5W6sVWNmGx9KCM6AtDCgGJ
rnmjeQaD83tRzgsumj6MfvvUbBUQlZOF1r6zT7gAMEDZeETVdhH3GFUw99o6VM0rv1vr2Lg6cC9M
6IBx57LMsbaVjkxQXRUh697vIHy47dxA/FhXT8K7EBdFReaAgYxVx1B/HzDKcQmlgkBefsbeIjE+
ry0rnHUt+NZ97cChJ/XWj5MXyG1NTJEO46AATaT/r/RiSEvPUbyIZdy+7YGYiC4C/Bgy0Mq8olC5
1GQzQMOZw2i2WxOJFaXmQjUhARUIVfSCKV5aSHYJzDTebk40GUfsIw5KLcPGPvWg9sc4bEvI4Nww
ikRZnWA8/ap2C/AK0Qwn3cEKPzIBP9KLoKikfr4YfGrSziD5TNBlFMYs0JUI7+QToQjwLjamzgQO
3i4fLGI0+r0h/cAp97q7AYORq5siGi+w4n1aI4R+1oxvZgtaGmNfh7ntzAtvQdZaspCwlDKgKgjp
ZVWYa/aka3n++Jn+Xj0P6yP+ZGBcHrANmX7DZ5DDqFJ9WRPVQWisgtYA87YzJVJufzUuxaW+7dQN
Pb4NLxIWVMRXMZjEvRYO9uQZOgOmuOiYwRywRZN6/Q0bCTOEB5llvS/LuweFMRZjhdp+bRe1Z3NO
Ti6/BWUWTeZlepAYEw0cSFPOJVMfe5hg4tBvqaFPPgbXUMERPpOfIgtLVd4Xr8hiU/Qay9ps15t3
NREFwF9K7o/U/pQ3w985NkxPlh/wa1oKzOamCLE2+4/eFs+TwweA8a6MauKroQ3eHvCmZBwcRDaW
nfaIBXu/fIicqFkz8xZrnstNV0AN6ssES6HjI2d0Ww+ONUihCHO/S+JL3AWSOtF1QU/qdFEaQ2zr
cMVth3/vk42nHHAfHz18XHOCqxPXsi1t1DfypKTjkNy92NSxgTbBQILSEjgBXX2SuwypDBiLAaZ3
k+2UGtZx9JCfY1Opw/jpvkUGm/7n+flAlycvim0rCpxgEp0F+OF6HWxY5JM2QPjrXfrXAc8k7M+D
I8cTGGDECRFo6jCHiSSVCVAgOwneT6PuLP29hx7dVLcNRXAXBm5XTM/yAlwxboHlYSZ+FcY22bQw
tXhRiLKtX9g0zAXb/ePuOIbjSFyUkukwYMl7JUZ+nDuM+dTogBmlhMgJZZmfwWWhxl5M1huSNRTc
YsrpMdSTJfZ/Y6VsPsrHJ70h6SkohS20oUfVZFegEazMH/lG7SG0pN1ZaEk8tMdkJHMSiHWup9nW
NMDQfSd6KakUM9+va5fCB8KMYbclM4+USFhNxBmu1pQb4ecGE06O2La3FeTkqEp+EUrdVth7h0D1
QvXERCmaEdG0lPemccxZAbekusT3w3xycMJ4KER4+m1+ZMzNItQPvQXh6nQD0VIkIgS+9qgW1a6g
znTiWSNhlS1AYjSW2hymilvA++Pct3sEr7pPggCz/FQ5ddSxHVQVnHLx/IvJ4IZXSQTezmj3l6ue
7Z3zSZKkdLAjnXlFFiWxsFvo4Js6acKwva3MsDPei298BRhrniBs+T7LNMq2wWjJPcaPPFlHlXv2
hEw3mmeq3k7QfPds6ESJkt6wWmVeCIlreEpHWPZycGll6qvgHwZD1+QTrE4ZwoMc1P+Hd1DSi10I
otb+KttnGWAsF9q7qyBFZw0HM5jhHdBawKjcc1bj+h0LkuUph4DHE9IYogEvZtX8u9ljU566pV5K
WOY0jTE1zwz3hWnORJIs0Df20T6RLiuDu5wE6ODoxRM6TOLwros0OEMcGMYsO3PkR5c+y5UnGCeP
I/bIH1UqX1rDSobCqVrQqoewgvKTc53UHbS5IrgS98RJpxCD7dOyiKkO32zMWv0OLfzQMFJwJHBr
jGh6FN17ZzXbbWZ1csmrnmtmB8BAulA7ZkOGb1jCLHC2hL0tvxGmyGP7/LmWK3MySsiY6DFjSw2S
J7JvDTIMJa3QMxStSKa1eprbo2z0riTChFaAeDG/LtsSzP8DtBlREw186VCD2Ue7jQb0/B538UeR
8I7yaEyuEUfmQW03L52Xcyvh8ValwW4qwE00F1GMaH993gZDnxj9Xqded85ATRJBmbUaTo1+mnCm
X7AzZWflkueh7DqYnlGRNp+MAwTGhqPiet/XTJX9b/lgNvQSZKCV7g6hGHKmZW97ssiskVTgixWH
r+RLPhv0GVv5MGjgksJNTcfHjNcob9ZpWJcbjI7LTfrLG4Fbidz9ulnYIgiREf4SBomSMjJpDPjn
6/gKELK4p9Ml4kfkAhGiPJXRll283wfxtEfK23lHqqNXrsu6bF4IXcILCpjL3Np5Rs5M67b7L11c
JI8aABL97dJR4YRao/cLMn1XbVONvy3AnrTXHRx+Z6QyWISbEHxcec7tL2V12hC8tG6prj6SYsNt
3cyZRPh9sHAbAF8UbEaYwrXw4syyIEzgiAiJkkr/XaMDCV7deBBLodE359fdGWu8lOLr1/jqyQIl
Bgeidl6fGyAGAujdeaukWWWxm+83YXz4yZIkERjR8sHjCBLHq2zcvotJEcd/+CMlm18z8pU6oKy0
tW/pzgU2K1W49oP4saQyxVwa7EE8hB1POmUKoigjTXlErF5VowYZYyLCcSozBlaaFwpWqtN82iRh
Wnj43JEx/DwpJpJlWp/37cirm7kiJW8Hzb1DrIf6ELkYyIBHXacvo+ilAuASTb/EWu9fB+6buS2l
Y2Bl7uD5IiOkB8FbIwXS5+9pdJjfTAAuq6bdaqy7cJ7RosPiqIMxHe68WlUmo9esFg/FsDealq7q
Bra5B1GhoHHhXJyjiExjI0lyu7Rq8dedVcolAkT76vVX6wdRh+GO5AZVIgMwADPlkJq0nBOaMaIN
L0kSjTfZGO3v47fdNzke4WNbLEdWLVR9m1XisJD/5IFKgzTlCTLASHdv248Xo8/vVvtB4/YxTD7W
zmnerHUpgs65/CocvGl03RbaUUhmXuoKAezwk/v6nXQanOQ8kLsN8HoEAW/QR927M7iyHaKCEsZE
QLdx/HMfYlgrHvU1lvl7Xe6Q3+21OhbAcAzxUjIyXqLsHD2UduAslqMI0m6TJe61AFYax/vzh301
1Pqzr9/bzU+z4vP5B4V8zAjNRRCvH7qlGEifpLDrwRsL4WuHyeRQ4+1CrUhjYrQyfKu5D3uoD7eI
gWW/zh2kUd1ulqjp3JzZemI1oZwEB9ObL6fti7JrGTytcNrWtCpGcODJ+lU/B4vua4aDpXAznNM4
yOFfKQGBTiiYpUTKKvEkdERxDoH9kLMjf131IuxeUR9qJZqMIL483SdlLhody/lezfPHlkhtFgyq
o7ZZ2S4YKINH15uHP6Y8fugUlpf0t4WGc+VUrm9MTQa/rM8aQv/re5K6Bj36vBfaYQBbFjSXATFb
VMmwoY+L+hW3nUZ+nVSyqxJZVCQeGwjwALKaZIaSd2RVvHcGcGo4I/zQEaeLFrK37ngKvN2RtF7/
FmDtt9/+UywvcKae+CtTqQbSgEAqbGy7A1CPOV3yezh2aaBLeskqRSoMWfU8mMqwHIiLEOHc/5+I
+vtBfCCpLe6TR6y9DJ45CnYjVTi6L18lB9PY1gyubxxi318kkyP0oMVk6eWTPVaLwdhChGJV0Kt6
haMpEFIpuVH9ty/0C3IgOW6qQNNy+hVU1ynnBuyR4Y+fMiq3pRXipDNkGYLZk5Ph/iBVAJD8WPg0
px/5ongBJ7/P0DHuNoLBD5tzLDpKgxXmWjPprUz25uKnKJUNOqJgzVv6C8Ki1DpYi2oHZsQqIbml
75lvMdyvQ050yGuHG5eCJv+h1XcSZY4jDPEZlyJxL7XqMI+IlJ2fhDPa7Gr8aTjwb6VgSRMsuFoj
QCfiQtTIws19124gAVhQKalOu7VDF0pG5w3J+EuyOFyZ7abUy8m8t4DDZu4x5WdwMFr33sMGWpTQ
6bnHlTdh4UOHb+drS27PnE+vi3NGa97v7OCRcQJ1UQInkdiZxHBmkTM6rKbNLUNKaTd9yArXxLBK
qetO2XXqTocJJXTTQPUZzAiy0j+gSY96ZABvws9IqwGZTwpbc0JpbR5IO/WydtUanKEg4+bi1NHr
LSgThiqN7mLQF8g1V+VP8mAirhacVruJ0iCAeGEMln3bA7k12+6k1Cz7YNgR5oTunNAG0khfyLcv
l7MpDYCCSCCvlOzWGb6ZB0Mlg/XL+tOwvqVHVcsnLqfszQduMx9VLZe0EVt5MAb/VOE+XAeXzFx6
3DZtmA7fTmTfoVAquMd75NyLJogFpgB8W7g9DaEsXBDTsJ1q+rgdPHOSOfkPUTS1GomGrLPQ8ZvL
JV1v1deOsHG3KRKqWBZNvmNC1bjzVRiQozMdQIoKwL9LsKjKcyT7XFu8LGsHUhZm4j0fLJ/lNmYH
/AM3VM/g65FIK8GzmY4XgeTo1b7JyLQvucfOXm5VlNKMB/ffUGVUdjFnSAxzzpTWIfmf8vyd3Hbk
DA+GyR7grptpowZX9VfC5XwCKjn/PIMijkpyxk6NBM4OHaIXQdOKw9rdVgF5HkfHCtdrLGkWmjaw
roXQ21IgY29tDjQyRKlyzuj7AUcBbwvq3ZA4stzi/BB1+Paen4hbna+c+f+OxvK1dxnVnZALasQY
ea96wi32kHcq4YAqxEPxdpNClENcJrlgn34S3kiSBYlNKUu+3iy1CheujdLAd+gZ1N1kanGDARWa
y31o5F5jhKhYKMn/V+a+flG4eAka1YSDRgdZpUXsxrOv3cYTjcSh1KXXyv17ypC9VJZYgLLlXM3V
b5fUfLAMKcZ6vOMnebfNsTQDRQegB3sbbEM4FMxH7aA+ng+s1QUDLx1fL+TH8eAAhw1UTui/KMCe
3hfkN9mWnGEnECIWekZk3Ssv9JjRGCpJOQ6Pjbfr0g1fb7ge33DP7N6LyBqX+2UEGAfkNkRnV5U8
2dFio83lkOQto/gdVHtotYd05bAswR2KjFAbA5c9HjfOlxmcNe2v3l6seTAuba0MEv74N4oMDx+f
mGu+b8YcJ50ln4TS3K6nlG+b4Xw27jKtQnUrcjAkpfg3LGyeK4QQZq0FzPBMZj4x/Af30d73AkaX
pC4ArV3G/LUsS6Hh9kWQlzy1IbK06WNMnK6CoLsj8SHKGBn24nhTK+vren0Xqv3ipsHo44AMvqZ8
uRBW3K9lio1LmrG0AKgl8bA/0VpPxU31mBnGYE2Z9EsN7DSg0iB8J/meFt+GsyUdwgQbAu5Y5BGT
Lpc8b4RQB0/Ncy6kqRT00gzahCA9Sc2p1ELq0mnoXori6rKLvX3a1KQBU6GHw8cJKNU/KL7GfdEO
AGysEFPJyuABbtBAzmMQ5uBCjDubrMrrHxoiyzBsmbVQLAe7zfL56n2xzybmL8fy57k3M7IGQP63
RpF6ZxPyMKh/v95UiwpX6p1IhKeuXm4CguFVg08z317nBHGq2fcUC7SfTL81cwU6QL/9GDERzIx0
WIL+xLP1Ht5M/ksMB7ZASTAqQp3bEormwzChLY3JYByzNd3ozBqnUhkhys17au1GG1Q6gvM7Kcc0
EyF0iW5NNh/OVPKcguhNsoIWgJjFUHU4/y1W1P7zuV4DkBGWofnqOdpKHipWWrVXnZF61VF/HEBs
UfHjP+UDRj2Lbun3QbVkXeMCJI1dEiggXo09wndL/aGOjJEZ1dc+ouCACYghqYoJ199C8/SbOT6z
k2856gnY7JyqoS/AKrrdmlJLEa4Y+If7cpU95Pu2K/VTBr35ejKsG8H+HKIk73mTqNfg6/tLvsgX
OWnDfLUkQfnvVHJI9/rmnh6CQdVgBelWgFg4W3SIJNnkpmR0dz45qvHQxSmBzoZiOQGZvYZ+daxy
xkjHpN61GesT3gxzF4MyKLR9Wiy9xIVdEQLZDgd97c8ZWgVub8ijLunHqX3Yx9RQmIUYD8qIDSAG
D7sbcLLAxeIR/KCCH4+RPsCL5HJfco53fCNMs4l7W8iHSAZyZO/SP3PlkZV7bhJznUyGjwUZP8qB
/pg7mnd/addFIGr8TV3ROPqfRLNCxGXWcGvXheNn2Q8d4R+ImZPrL7n9gv8rzHW1WzN3jLfB1QlI
mh5Ox3OrytYTOWmdO5KCZfKpCuGI+kGLYcDMQQAwOH2dgmafbUq+OWDnnbRLEbimGSp/cIPzqbzM
abp7WfZzIe85MAEXd48rulShLk6SX5VRiqGH85squpPmwzIJWVDhVHlB0mOaH9elpyGgYPndtmmZ
9oIYSB5OvflfV5FHlSbBZ1LG0vyw6uy3V8HrqqZAjYDBmKnBlmeKnB34eg/8maNq6hPElsFlPZ8C
WzZKFdTnNWvcoYzg5/IsuUITgnfIKybbLcG3K/4jMBwrvvUhkcYFYTh2Nox6e4LMFvXlMu8sns1d
YwBN2/4t3As80TEpSvuKeAJWxlvguYL4i+4gRWXeA/v5mDqck9IbWLvlcQIpkE5WhV8QGWeiUUN2
+FZn55JZJLUoy/0DvW36Mt0JIkSwQLWiTqxcQ+FQXNIeIP1uYxCmUSJe766w9UkrQIbbyAXtXCaq
PAv45TvDrkY/6+8U1H12Cr9BKrxAM+bayTKbBWo0lEwCFZFllnF2YkHz8wzFVSLMZJdQ0a1Nrdrl
gzCVyr3asi76/IaYZs/YS53W6QeYhWIppa1/LeQyzHCGYrJkLVbZtbQ561sdOgzQoinlypQ/Mca0
H5TtaQU5J95BcLKQQarMe1l7t2hLkEoqmmdHL/z2Q8m5MXmDRqHTZySJY+/+sUivHJ/wjTLSZTnT
anPifl4o/hp/pZZR/KvzzMIrUHUcfNYWqthwu1bQdvSDgcSyJIZnNrrWRC0ozgNsg8RjjHTjDw1e
F43wsK6xSUV+0RoCgECjp2c5E9ae/q/OeIEtHNVW3RLTZhqtbuNxPC39xn5Y1J0d7WNB46yVRX6R
tFXwCWSmSo6pzmZICcW2WQHH2094PjRokqzNtozpEJVFHRxWksGilTTm3L/HbEkdAlNnvTD+96zN
SHjH5M0VKPUgshpKGoKzv4WfGL+GvReuvk0dN8g5vkqQ1PH/D7emnlqkcBF2lYmRmbehqgcyHRYA
4O+7HxDZwTebiDIy+whr5zhWoHZu9c89sY/qxK/Pghhzp45AOisjxSG6sjsbgjxK/krAfIujucev
fBmcSvRR1JKTuMF0jmnhirv9M1mcpc4kAHNSi/GeLhepTE2uZElaWg9B8lxlIH+ifYCer4bGasfD
h6/Iy/o1NJfBmZoqxpMAGlESVd0eq3yicvvIq9HvVJqayGVDBb+StM+ZkRu42gSxN8kJBWB+NZG4
zV2mtmZ18OXxZjOzfjlqIBdB83Abj29jkgzmtbK9cuZB7o9Yhl0huAgczW8CZyEn33GDQ8kjd+XL
YwDcd8BV4mdFROEMODA/a4HB38nUJzujHn1u0llgCCTC9SUnjkISj/CTg7MqDISlUeGMTGmunPZq
dFc5QGIihl15QnLlzI+dn3AwPAnyKCLIirO2xnJa5HcicCNz6LsRWgazUwMLhjGvH65qhAdsBF0v
EaX5GZQkxMLNDMDx1U1n8cAlfWKT3/bhRECK02WeB0cZ3pREpDnTdtTHucq3oRkrzsRb8WiD1XVa
KFg7KhH05S5mF6GPlLR251O/JJ2bkQlhC8B90O+Fk8YrljQDzekjpZMcP5xZ2ruV07Di4SVi6+H0
Bn7LODshpXojczE9l8IeduO8mnrYnrxEvE85dn7lOqCSWforuGcoBSF8C3Qu+BdejaJoF0PzlJGb
ZxahXgHQzycugG6kMaGhGnt8WbtqWI5iPOYouxA8ZbAJ5D3njvovLSLF3wRNw/5AZVYoFIDv+OpC
IJDRNDzDUxOHieR/5DwJ1QqropTv/dB4Gz3BSFgqlOubszwjxTadML/iKB/k5Nkji/vHRm5CB6NU
DPVO9mMyy42s8KsI/jtxrNXLtgictFxAxIE17hdE8wU54YFcnz3wjhNIPic3BnmjFlOw/pmJgboH
BXF0UP9vR+iteyHA4uIJqOwnntZeKzYUjFRurvypGKFzTGIvY0MpJQXy1BTl2NJWWGt+NI9bP99v
enFZlE1FZsKmlBGw0Ak6RY6XZ6CZ25zcQjrrk57sRa11dVXVpOuKJ90ZL7vmsqoqWsT9VUlCupbg
9lVE4Lq619l6OIjq0F5uiUNkigZNn0CswQAOXgCPj4NIxK1sFGya1BoEkV8S/gmGggvQ3Lmu0TYz
V4B+axaZHjgL+yvRkQpv1/x6DpJiwoIuXjnD012uA/nhi6OFezk0EyzpfuAtfJPfAya/t8eGlqy2
Nn6Vq4YXX2Ey3Y1dm6IrWwBdbhhXHrbEIztoaoZUjHpUJud3S9+i7CAuy3HxCsIaR1jL1OsjnrXb
qB3BmJRT6x00DWVakJIxRjHLoavsnxaNz7uYJGmljbMVi4Kgr5xNi5fnJI6dNPiBX2l99h2Ws+Wo
geS04XCTwwtqoHYEWACHE7uMRVlWKdvi4D/yZnFdvdUEwZqrwQB+i4kWBiZDK0yc6HlIl0q3xaWc
oQ0yJPJzsfejzXwxR230F9bG5cCriAVl3YV7e6wqn1iKvlTojGlLJwf4gHb619Y1D+wuqfmM/lv2
LsvrNozBDe/R0nYIMw52av9nmUu8pNTehzk+2HuKrKO4cqtuUBS7idtkyGMdorKvOnFIrb7gsCuM
ZyMenlUdbEFMCncWBFvsowgEZpRVVE6oSme1Y8vn7MX44v9pGxCEMznewvCXe/OaxqU9+N1hwmm0
lolC3UTnzHm/2cXYciQ9IgJYbMgiywJ0wkVw+uq7Sm8JwTDMBlQTz3IfGodUoN1XiwiAx1Efdn3J
fZfBdrdJWGGOCVvtoZzFjZ6JwJm1ghiCn947AxaYjRV0p1ejhGqCdh9S307N9OjEu8x+qPHbD1bY
cFXRhN+bf3U+Se6K7xJvnqrLGZ4n6Lq4M9HMfnX3f8kXXMb6Zd8QXv8iyUfhY9QupCLbFi6wgLsY
08YAuXtdabQdRKY9+kALnGnGQ36Po6OlEhFhQM3OpmRN7MvaKYjEQCNCf+1tEgS0QBQWk1J/f1pV
ygunrTfMtImyRfukopKjQXgY1LMJxmDaoJa7HWYd6NGAplqFaAV2MT06tc9lId39bpQnD5IY3AqI
mrCM6f8Yg/XkRUdg/tqF8R0bPmYrSfP2hXD4Y6ohGx+bW6e216FCHOHlh9CYK56VziwcTWN9ly0D
almAP33FMvUVGON5J9JW3OVSKE8/R95COtFENX23X5DnH7ue9YsCdtFLNi/7xwMgq7uSahay3d2/
pNjOE8oZ2mykiVW4lU+VEMZZpQH3cjF/IZGHek4YNn3aXBnyK7g1w/96NnBaaFAu/ALWFzSyq+k9
Hm+JBFTaUETrOnFwjw2DmPy2eDEkYYsJ9/5K/aiVTQm3J2xBZnveTiH791MFmrB/dXO1cUPWnr5S
UMvJ8lApjSBcvHBE32VWGkH1Kfp0Hzy3VgDFQ6Jpuvf+Fnd1nLNgMwiIE5fJq1p4jDJMul1orjLY
cPqTeJbWGgL97wB6TACgo1Eqek4Odljn45jKNcQUpjwLsKvvtkUAaOYTZyz+bRcdAjbbO17XJxLX
/1BKLoedOB4DLiXaQIircOzIecNhGNx/XwQq1+MZ+VL6Ze5+8fIDkaLUhNR0MVZ6jfHZ2OK36HYs
2OrI187+4vFiAAtZ9ZDh1mIebaLOtVawV9yAT1Qt5vJ2I7hQUGz6zpvOMI/V81zeu9pjkjnd5wwh
EQGL9bL8pyAh93+nCLa0IU+N78q+i97rtpMm0j/iR19nsMKvwGTWKJYDUE29WI8/1PSgLj6oI6Fv
Y1X/VnJAt5J0Eufjw6S8Fnqz5W6qkOz0atsRNkITq4dTdL9aC7XxmU3uDdkaciBA2aTCn7/thtNr
phmKApfM/OiRdv9/OlZucpv4s2DU0/HEGJQVdDkCZvH7QlKMTBbFWJh3jsSXsMZgZUezJTQuujBD
51ecJqsj1QBaQUwT0RDqcWcQNAO8LDmeoIUKr4blCstz96sNO8RRlIjPyN7ZTtIsdxYBQCdS6x1C
qt6bHUTOEcdrTuF2mSS7rRYYJKOvr1hqHKEsnGg9MSVfNH9THXu445ndGU2T3ADaITRAywf/g/i6
hvuxCqaMuhEgSXkg8iQ933odxFjTHuLW0BG4UE0YMOKyci3XxNx6v0JisH+qKuYx8CMF+/hzLUeB
cjCGlrNQKhcRMk6EFo/I8/M0ECt+98kJJH4zIfAMg9bXPmY9gya5lUixnfsvx70runXg0Pj0v4/a
0hFl/0/mbcPLJB0mzwVSpH0m3BhAe8v+lN3d7AJxM8vA6bjU0m6iBEhcU1hFokqTXrsdNXWNeDr8
p92BuULIfcPygiqtsvTouzM82nEgFZmK0v3vCBVG1ee8q9eXLl+GeaYvfQyaOTV90xSt2tPxDxT0
dy/jvI1lWeXprf19g0lvvADjHtJPfarTvkHbZ/H4nKCERDdlCO9QOIAtLuaTZ8AVWFyY1rLIwn0A
DX/swY9oa3M2DiVbvJLwkYvQPA5I5FuEyDW7s1893HMY9ZnH7X/LIqgHgyJ1mSP/fuskXTTfHdhV
Xp62DfrN5jC88jcY3n/M72WnulcJCZdKyYBGFreK+kPN1rI3URXnRAfmmg5rityMp1WYPEWniOJE
sgP9J8fnOS3C+DqEoXPZhpqBBLUJRemxj6je7nEUGVPEnjZigfdtKMfgABkYY7tQ58yhxqq625rP
bY2dXYAexs/v1BJ4Z3sRm55P+HK5B/vfCSXU89rcikAF32uA/bFue5imhUEI06o4WojV3GaS9K6m
W/SeJ+lk/fbfsI4CVDwARZBWfxhv/JGD9cJHtXmZ0qsUnGfsKsL/zOXi5qYsZIJoM7bHPtPjrU9s
NletCcE5mdn3TVme9oDsGXG0atRGVDo6ziyyfv23g6e2coxkL18a96y9v5gusulyjBc0dRcaH7BB
ZvaPSPvaonL9h9Nty96e+fYuR3YXs6pH2nkbb3HglL8eNRt7+4MHtPwd/Tet2aZw83YTf44f84Xs
3O0WT0nCrC7pDqLBJAwqcP7JPkPgze8tWF3pRmqcGJwfRVQWA97zHW0Y0+59Tw3J2VwL35ls8uKE
YtBpphTKWS+h5j4kltpMfh3EQpsqnxL+Bd/5oVAQHrUYBKgIOxsL3NcuaJBGF9Lk2bL2cAjXsQit
+V2BQYJDsHKggHRcjtG/YaankKfNQ3GoWmC7eRr9TXqZtlqDBREurtZPMtPkeBt9S8eDPpb1mPcn
jpTNVNL416BwXAGyfLb14NkgyPuJutTYRVm0+p1CDf0bUJ0hsuBGlj4zPIAp+ro5nWrLPZ3zhp7k
0NEZki9M+/eFLZaWLcAgtk7EOvcyDgADkc9QFukrot3JQQWJu/lG3dwYHzF3ZiBN6VA4hTwKwxJJ
uw5xFxkswmKboJRiQLQ0uNnsPDbo4VH7Nttkihkmi8bRyy+VeI7mTKuoKAXdj51aK6EEyOMIna3U
ZRE8KTdHVVQ6l1/X7udNeQZkJcgwl2lHdfdoTPKL87bROH3/yDtxi82UtYHDsP5AHLg+wByw0m0c
P4NT1fy5f30J72u8g4l7EVKvcU8kVcNRIY84hMD8KhGA5lRx9NV8G1bwR0Fa/2mbQYZ6fRJaqFuQ
wAewey8wpjIumE9EVpqjtiy5sFbbLgHPlJdoyqzj+1fg2cOQ2k8zoAi1EfMvtz/kT3L7nK/RxcQu
NFAEaTcfBLy9F+ndjm6FVQy7fMOvYjigCZnq+2Co1uvZ2atplcj1K8P75LWctOTax8nFrXcRrTDG
llxrahuVjCWTwcaBz1tlpstYu2aEjCBwZcaoP5wHVBdYTynEkuNUk5JWuvjpMw/hCR7zUyQDmg2G
QJj+7tb+LIlsU/Jv8wolxshdRlnC42wvG5BZsge9iqEkEWs4uiq2j1ywM8C5SEY+aSRbEJFolVi7
VaG3mDlGPu2GU0KMHxY3eQADOVxFkF6o00cPNoWSC60NjCHDL0mQqsMp95CfBtIx37ACmi5n9Ty8
dg5PTVEbuwc2Lugxoq85qQah+y8bxqN6DGhMZRxVlAEUzJjozVHjvtjG7QWH+zPlmKd8rgI7hoqq
a+N6S14VTBXrtcKtrUC7bCAdkkMaloWEXKfFSci4ZJUuMzFxSpa0ia+2d8qad8Yn7QnSKfOSHATL
TEYvZmD0OZGzMmVOb8uVTKguGrTxNXyH67i1PpPsGMMxTX25MmjTbBah6AVnUrDEA8dkTl6BqycD
H3D5xLIce/lcRsBidS1bf7E1kZSLh9pQ9Q9WJxd4pL20YitKlktLGhvAjtQE58pny5RCYReJlgLj
rwl7ffnwph3Q8YaWcrpJUbj0fxtHS6LiMIuxCii4uHWHpj+0fZx0/7NTNKxmdSyhC6txfpm1EkAN
qjO89H8g+vqpJuYwRjNf7lVU6RzzlvE6XPaUcrq8DCGV6vJ8+AyKZZqkCkavhntgHA4z5L8YoO3e
ZK5BEXuEAE/O0i4ENRwfz7IMSXWvFp1M69wJ2kWGZ3ZJae5IZg7000wzZrZ8yB+3f4XtTRuEAxlW
ibiqxTD+hidAPwJ3g/HEqyLMOg3HPouxUhSdqie+bIZGDd+UrpOQK1jQpQucppBYqvwROVRdfiMI
8ff6KENUG05rlwXDAe8s5WnsYB8pXJwqFrJ/57YUYyYeQpsaCUuIfBNObfAapK0jV0WnYj7UviWe
3G2J5xNorTozQHR4eyIgEG0jHyaaY59bq4zB9TzYBksfVbyKPhoa0NPsMSfKg0gpm18bRI9oSk//
k520aUhAsKxQ5gaMgIS3cD9Ulwl37THS6DjhBrg/Lr60MBRmqop689UwCuz84IM1D8OaukqrHj1Y
/xWstzed9qQ1DLtRR8+txU/Q4liY9c+Oh/+0sjM53kxTMX1H9fkwStlzkkpc9jFLi6v0Us2rqvwn
5uZJbzBR3l3V15F5YhyMg2vUmSxLh1ZhD0lSeC0/cWy+W6zxQHrGsLEut8tFpKgH3hGRQzDklrHk
wHKNlUDKSEjHHLjXZY2zw0cnpopXvw/sGSzc61APOSeEEfOFKdkOrdto3ix1PwJyOeTrqRidfyTF
Px4H5+MG9MbowWRZ9s57i40Nx3kAwjwxPD0rkgUTNU0UiHM0R0GhuKNGmCm86cFeIeuC6AgFg09Z
8zT73lt1oO9iLbyrMTXL2Vgbc2QJXbC3W4BUAD/g8odLgyP14VUyCZuUp8tbOw0MJF9wm95nOJpw
3Qqu1Y1nUj3vuJmG6nxIbXAQ7/fwJD8i2NAOYT3rwJBy+uyNpSxAxgLZICUqpm1zQ7VsPW1luIzZ
vrJQLdf9ehRXO47kzMQxYILEfLP6aHE/ZEff4xSKCYCxaQ0OXFyneo4Oq0Li18HAZgOoOLpXTWMw
RN0rzsHsRMZcVGz1kkg3YdVxLuJIb6oFcw1p6GEymDQaZ/nzMDOso6KdD0VxsAkNxgPMOgQ9/sSe
gz1z84oeEapXp1XLLbNxSE9ye6vUyaBqNIfUYbab1VxU8N1DJPTdPs+jvX8fefumC+mU1H5AMlir
2ipVnxWjnmVE4HqUFqaeiBVadPl5VcVrDwLyH9HqbQVE1sYqaZ1TAV8DRaNwlSisLh+olbJjkayO
hbnAPVrLJ/DO8bn4Yr24tVX27OHD7vmNALR0zmrmDyfrt6g3NX7LOQb5+//tAc2ham0F2CABfFMK
0aXz5zCup+5fDUT+n634Qtg0mp69wmipo37i1LZshPwWDvuRBKZGw9N/IWKUuyXPz3MNG6+X7PGJ
gUoZIUJxkYL92sL6OyKNjoWDwtx3DIS87jF+Y6FYrLy3WgiIVh+SEtNItP5W/DjgPQRf6E4wI+iz
gj57vm/edyWafL7JDuFfLZqcq7abx0BUk7TMnN4UdpRFhpw7N/ZhWBqyvTnnPOvMZncSpfBPu1hB
5V173qf7Yfe+zwh1x12S3W61qA4OZXfativBHKLjmGyOUoEyUHFFVVReiJYhup6Bkp8hwlh/zAbC
aWvzyuY1f6K4K7b+QDqRNeDXSVipCXaIplIUMnBrsGzl0njQmMi4DFTV1txi70+wTPxNnsULCi7h
8jeBl5E/8+z6OiqS2X0fZ4I6GPcXPHDVl/U4McImJ1kynmi06YuMhf6b3LshYxvuUh3L/0yF0ll7
v+/ABWkFhjkw76C6w2KKw6/rvPli32gTriE1js9W/0ZNN7kDntvUGHqttKettJpNiCfoAkt9SXwS
w0mT90m3H5YwWXYTWkqSKk5JLjNjZCJSLxhlmSpDyRv+NEZJLW7G3y1zK3166avB/8AyAV0MmOTl
9mU1+yPu6AzYy2zbWRQNF+GWgeBz0zzSB57QQwr75oJ4nICyUaUO0SA+Y2m+k/+4+CCYeA1NUfhO
/pYszSimZXA6Bqg/xVK8tKwcvTdyfexjS2N6jVgrWFtXmTh2cMzxIvGr8M8I/IOpW8BmoutGxiCS
OvJrQQTVfGwRJ77uhEwiAOnVZ3JwinGI0S/HGQk1/jakmPWp+QlSTFrchg/IxuXGx1PGTG21OcrF
/3aZgT58/n9vb1FSgNOnz3nKuI9MSitID0sq5sKOKXnsqRB9ige64nPZo7s264godYipl6edmDGh
Bw5oY+6jxyIb340GGsDDVDY9LRQ6hc7k8wFJgEJXhB7fV0yNbSqw5vgBpRWUKoaQ7RUQLQUUlsp0
/nFJXsbNeF3S57bYz3MX3oYD6B4SIV2/Jk2b2HmQSpk9t+pnF8iKCsHUyjaSUwbsi/FUIDih5Plb
B3gBKmQh5cTAt3dAlNCp19r4sno7F/qUlGEMze5h2UjS08vZE5dThGWvdKWi16B7a6XPHW0JqA9U
Cq3SSixszd7nnjmJokYjbq1zI+GcYgmb8EKQtisaM+kksv9Gp5SI5til3ByMpsL49oNgrf8zFX5F
/8gzMbPhfHbOeihj67Q4cv39BExshAs0gNoUEb2y5kpjaYviVFyh5WmE/LpCrjrFcme+9Gfv9bBx
L8GGPE+l5xZycYYo3FN9wDXRiZiaY6OLlr8ijsTD17ijrNrPwewL+clUFKO0i9rWJ/6q+11VbtAC
mi6dUkgtPGTWRcnoW6DfqhzIag+l+aq+2xPmR3F4whLW2q82S/BDqNApDwbmR8ctlXXGJSmNAx6r
uHvvuZA3LTs3nbwvQo5JqknkGZj+ghZQIHAaYzbxTD5BEb5wQUOfinPLksh/BL3sXxoy4SqInF0E
5L8+D9nT9rhatZp8YHKXAmC8+Oi9zTdx8WDDqfCtmyHdaLxe5Rh0WezM9y/rf24Q2UToebATd1WH
yXFLag2uAXD3sdEOlSz+49xXgShI0IuWB+ixPlmG2JdVrywl1Rmsy+xF+bgLWnIwatrFuYEu1Vmw
iaLgoAhEReeATOHTwJT9y9aiDSviDtaEUa4mTGyRMAMRdAjYeqeEEZhouYQ6wW6/L4439Pabhmov
AzH1+Bp5SMSB4I+5XOnP/56p8ta00lzSCidsJKJ7gfMyjwX1jxey8OH6utkpAlFPjPsjroHO0muo
JNvkV0q5veD8MPMR/9leoH/nlieC0VnA/wC0CEBOglHoN04kk61C3PVpGhcLHRnrZruYRWxEVYRB
SwkHM5DFwG8NzHHI2hEE6S4HIFhQha509QtpMLB6Z7uG8PRSwUtTQmx9Rqd36iNNgrYZF+jAg+uO
7sBfbqnmkJmyxrZwaeqI2mMC9FdNpDrX/NxdwsDC4nEHycsjy12IpbD2dzuhrVtNwAXrD3I1HJdV
wgYCsbkro+KXB0yYLAiHaXO3wqEXr2bwFkZb/q2ph0ahLcNFcABQe+rYzznuD7SsMlGrc793UVB2
lTvfen8DiUxpLXRgYIKtolSKJSSOTVGKW8MlOJ1GfHcOOAdv3BJSh3CWubZWMhgs9AfL369nXcJN
otPvNzmzMmwX0GWy0kTuUmL7eao0dFIqZa463GX885BSjYyRkd5xK9CrDGgZewTyqFUD241VVTWm
+ZvN09nUt2B+TNy7eeO60NhIYGjJ4yrQtl239XJauLzrpB8UhGbxqHTbTKH1Ql3bPf3I3MN3vJZW
9HVCTIfH60LVf5fzAFVQhCSL2j2B9r4EChOTtaW9hXJTCJbKP/uiZzlcPcn+nFE87OCeQzrj+RNQ
+pAb6ERfqdg981lZbofXULUE/A1L4uxjrEMzDwXO5EsK2UsyWmY5I10LwpmapAkkdJQLhKOKU+nw
nf6gAOY506Ni2Jc9jxCToYKFAG3yqfquLJV7zIB9vHi8Vr0sHhQ0J31gZFnjTioEpXYbWcRG5Q4C
6fcmpt7fnL9vs/t9QNpnLa6ClyBoYIBBtWkAF+NHxbztFUnhiJJISsCm8x9DUUa3AY9YUXRUXI6c
E80x3NIdSXF6vWam8+W6rl1unq/9PPtuek+9SsB+l7WPEngzSm6F6Ch/YdIvTX1zrnDXtZ1obJJY
C7nzUlHmnwYJcln+C6Q5cWcFpTIIpRXh9qUhhr+feZPiO8QZ2rDJjcOW481riKFcw6o1d9hcgaIQ
Xvhb999S8Hrefsvo2LXru5vgTGrDHIMdXjToMpt7zsDnhUNx+w1pWvRlpkS8DnmxthnVOFUmV14K
Mj5HG2YVKtgojfLC/CveJaKEF7Ew+dwS4rNZ59bwlLr8r6MGpTYDLz64yMTjXQhGfuchiK/4/InD
RmuuchXX1az5eDGQxqlKTkrhujfdFkAsPLhUhxJwR9LVr09VWu70bA5bOlLE6rGP5hB9v5PFPD/Z
J3k4yh1qn7iHh8T+x5lzink4/9YaDA8r5HNn4vT973X8xDQlD3q19FtFuLrg6svGuFbV8vWRC+/o
YmnEpmDkSyJTpigaE0Nu6HIy7Jii/RkXJOI+fJswJS7Hj2VU/ddhC5tcbshnQoNkmbUYMxjKV2+v
bn2StQLxJsIrfGosuGbsgCj6NgM9Nf7zXOMdKdF0NO8+MWrzMh16hB92QW1fQKW/DTOCOIBQAdTi
2sk6FKXfE85jpToZWLoJ7vf7Qe0AddtO9Hmwiz/PB7MI/KQOBXRNVz+9dm468r4gPZ2EWpDV9OFI
0s3V269yhMPcp3wWqnij/T2GbDbcqFm0PEfKJuya6S0oCmv4QQKtKgAOfNWGL0o8k+lElR5xGxqY
oMevLDBNNgy9y2upMxpbF2YS9tBryArUvNLZUPkgwrStlGHkTNWhqvBl9Ra/K8N6jbWZO+UGlBMG
WHQXXfUTZ1apa9GcptQHerEjXDElXrCbLI3B+ClYIiGC1cPYgRxbjP3dmcaR254IqFdlBOHJxOF6
1J8vSLaZ3kqR6W/8cL2JWBxdLezBzxASNin+QJXXaeSfUEPXuQ8SeeRGu7vJ5OV5vPrVPUw1Jt9O
sajVu2qkMoDxpcGZZgzUc4oXhJ37f4vsY+yu7OI5RguiEc4Bo+HqHvCKx8amh3cKtxK2CUboRYxm
oCvkoRkQYo0NzetNbWHBnKYqHJ2L3mbvRNmLzXBCVSQdsGyp+CoNbTQ8DStYUYLVNYhZsoFYXAUn
fuRfQquVwfiZo5F/QrOhqrWasnM8aD251+cywhmLCss/gdeKhqP4GIHALHMDQWDdvarJl3zKVE2k
8oxwJujAAW+DoeHsIEYR5j8d5ws7UQMLh/rzg1kRsEGFmE2PBpA4VMzezXXLDSN+kUKBDNYE15+Y
wC3kK3u6sfQRqVnEPU7IE9Y2kuAPhihcJR1lJFqBdQUt1YZQt8DaXBCfo/n7H11S49MjBJp/2QWN
p6Lew7j6S7QdFmDnMswHeEywwZbxbn47WiU9126mFYLtMA6ZCd86R4Zek9xkNGX6Ba+OV64Bofmt
S9JcQ/rJlqTzRw6lGaIBpR8lBQBEQdHr5ad7pmdPb/xX+NpmTI6QKESQgo9vNuSurYczj8oY/zyk
g3j5CrjwlCzkCojXNL7j/ZJ/3han6+Mb/JVLpzdOdx3LrQPZEfggAiIluSQc3QTQmHfuYXXtaOQH
MKMHqYJ7EQGGwNlepz4rcmASelqb7Q5+LsYWoUoNuSs2m5Z/3MEMMhL+MwUtiaa8Mq+q9/ka3Vd5
CWEFQA/vxe6I71vaJcC8e/UEDA96GBiBkdAFgz7uWXL16eaMfRcpPMkP+2ubA0bos1PSk4vaGC4f
nNR+QUmBAJ2ukIc44EQ9AhPahgR0wHtIGa4y5uBki5HhOUWXswpoZPpJJOS8xUg/JQDKPRu/BY4w
kNbRh8tE5ZdupBTHh0GRI7K5dBLxhTWCJxVLeeY68Y0osErh2aGEJ89o4DbvSw0pS8s+oesehkYA
QGJdy8TU6bH7214DkKRFM3c7yn84pkXn/M35SiHw1nlAi/giJSQq1hNfEOapl4+0Fqf9n/InqM4E
sy/cvHp9hkTYibH+FSgg7i1HyShY0vyydjri6nC5RNSgPV+kjIrj9NNd5mlFNH0icW6alxKm1oLc
60LfRU8854SzE8UP37hmmY8zX3o+PnOLvaiDN3weZeakuC2Ni2JRC4Uuplbr0jl6uUT0jotiTn/3
VaffNWaR+S/Wc62Mokav8LUL4RQey26/xNvuYOnH4ivO8vnKW45xmVQEE3LigxOf8LnomycdfSEb
WvXgvLAnWyZq1+H/axRJXnfW6aYLZP1nCRjVQnNHEcEk+GdM0NcfFy+VQ6xYXtu1Rb4dwHvGNNHO
eSZPpmGr234knUONaTneJXxCGHdzxU7zeoIMBtx6ImB+kfm55p4P7mMh9B74al39vJPzu8M/sJJu
Pvz81kBox/tJpWkw7bBL4gExjuuzyTzgwR9MMueA6rD+rJpN6b1cKnIVHY7FjPouDmx1kmwjtTF+
akdiYBvcyJ8jkzF2T6/CAq07Dq/ZPuJiFGncvRp+9Hfxre+TnUUwXqfyiEd2VjlsE3GxCfszVvYb
jkwgNomCYYgi/lRahRg8HJc1kJ1BPXAAP9JlVN7v82eJAs7mnBoYl5edtPpVg0k7p17nqFqikT4I
MOvZ3PJ6vEDv0wfhlG49+dtLMnWBegB28e8aV2ro44IFgacFTiEgv2OIbZDfCfyb3o/7/yZcCXRp
ZcuvYL7VxaSJtBEI/hf7O7tLnxGp+UQV1IQCwTR++HFsaaT64Kr3CMrNEWNaUTVFBW0XCmsI1Jfj
ayzUvSH5jyR3F3aSLDxg/rEqHxtjNYpyMa7K6favjkLCYDkdv6939Ciu+wCga0z+qajZKOV2k79N
MsAPx3fSiFPZkguBk/wOoDUg1IcJoOJTRNRjk114RFEe7UF3R6+9jTP624sJBzNaxsSg72gPWryO
6FAbOpXD3tlymz8x+i8sprCrZsxbRnQUiFGA2aLL5s+ymFKKh7NWv17t5r+RcfzjzJhCTXJXv195
CV8dkofjB3MaioKGcTxnoE2FbnJWs6+3dtLMo15bRV+i7yJT/q9MHLpMNDUCuod9RhK27meofSzd
khN1dUMcprtw54CinU/5JPCTSMiVyq0dLJNR1+V9tViBep04zWZqaB+IcXXJd+VQCrNPD4k5Q9zJ
Uf2bYGN17xxGR37EAfDCb770VdDo7M3pvEVHbHPf2m8O2ZYiYwQQFV0Txk1VvQvY+ugCTkfuvda/
iX6J89ZYeNtWA5wpaCkpmVgiwyfVsaj66OafNBE7rbGZ6pW2wbwxQnBmpIFwba6ciQaOI4WX0ARM
9lPMZRimHXw2e4pBbP49ScWgGhz/EwBZFIsESSF9DmenLSnLPh2QxhpUiiiTXpvUAACHS/z7FWUT
Qge8xDvKj8QgHCm8+PYS/bZgL+olArq+F6Syq+10spct3/QYwJk9XFHKVtlW1cVapmC4IsCv20dz
ihAlvG/SLGUxIFLQf9l8lOsKYKZUA2KkM150fDYEezC5gwtaZHjju1A4Mw/hJ2YKdtSybrVUIILe
D9IwPqpd7I/WYgKliyE1aBdlvqmabn/RTfYCNw+7YNzeTAfmCbDZxmKAPdzIYjMI6RvcP+WbeSYc
61nBfGAgOKgz3ucmXPILvnb5NXzHsifktdDob8WV+hvjTj6RX0HQKLrBygk7h4Io1MqqlLJEB0G1
3zwcwhTfTvkQSJWq8LQLolGtfdzO58OM+G89tLjFkcolv4l2FVsROl6eKR39PXe6Yb0ddgl0Y7nG
3AFK9l+csIr5UP/o3xu4m5l2N1tUZKo/Tr11NeVSnxjwjGkzHc2yZwbz5yBL1uDOBw10VP2Y4XxS
dbX6P4NMAj0xEM1i+EzE3iw+OH8CbDezttMUr4AxYJRH0O+B9wtuoERNDEbJnfnenWQOMaV7Ukwg
4pZpvl9PHv0ZilaUS83VCgPViOk8qgCZQxBJDiEnf4t1JGg+1T0ayX9TJCTfg9w2nwa7LjTHDBCg
KHrVJa0rD5wHAX+nxhxcUjYlfNSFHzdojCohtdncZoLyF9UWGJ+A+3BB2jLshSl21AUZTpnhFSp0
YAkBsQRMJ3dYoXh3t05rbTdvxxjp/7yIv0cuFWAer/KgpjAklk6+Oexj9+xlmyqtsntaS+ntmd5Y
0N83jRHPlr8y4QzgPd+TFRYDl71edMqYEie9f5Q/wYC+NM8PZ9TdzaVOoDhwR6Z6HyVH21hOFtzc
UKacVtgWcgG2OAdMKqfeLpbquAQbI/g4s8I4Yr0g6xU9BZQiSdu8G4xBIVzj/Wg/MhOqZcxSyzdE
uFMk5Yh120PH2WLY9P25vRUbxA1Txq38sjbuzikj/CIRKw1LcDmPZ6WhECR5Cm6Doi4knm4U6mt4
+X3sbVDHvRhFHCEqAQlzOUx8JBDi8/IEAfiFgYV2lpVAhspgAQzbYBrIxd/Ch/Zp1m5uCigpmFyg
yLVcUPp3B5/Z+SBXFITzuXkCi7tITVZ6sE67hIvyoC30Oqjgv1feM0Y1EnS29BQ6/d4W0ejpeiG2
v+7v+XdyKyob5l45RDopYr5vmNvMxbatcQw9dhGBEJjl8Qzk3zHsHiCK08UQHEdG2uCvI7WtoDqu
kMPISzHsgeGwC4zO3DBYTRhmDMV0342PacvGwS3lkFlJpctMko2fD1TEX/RLK9dtTIPRZlRUkpzw
kZxVkZWhZEh4wts4Cf9BwoAvfCMaZiJ9H1wGqxwr5w2EuklGSBGe6IHbl4PbHAWZLzFN1muAxuS7
rIVNueXJ/hNmbOpCYXSvV1JxYHd+z1TgG3RmUqF6VvkYytvJ1viMuC8oWg5F5+Z8gPYUOv4O8fFp
0CFAthzogKlunN1WifJiciRCXZTEod6Oc2VqfJJODskJULr027hwNwg5b0QjX+cssHVx0BrJm9OT
WQpZlrkBr2CkG/wBWfr5Pjmj6YyDmv26LicC87e+jAVTpj8Ku8jFAj8euJSlXSSL9GW91cY9p9Fn
LjuyLIl0uU6Yf7InoWciDnhyALngZpPtguIlAiLhPSyNAN5b6JTOeUIS/0ENDaOpmjCJPFVBHPwR
+KDgWK6hX7NI0Sc8S6VtTOAvpw7QqlijeVdBQu6CKoXbXxdYYHBn/bEwqLukkRa82c0SSfehOPpr
JxmBwZ0JaNorS0a7zV5OFjJF4yWH1Szkx3VbZpdE44WX8Z5XE3kJi0gXV+ssbZXOjncMq8A5UrWP
IM0ZIF0Jaq2Q6KKH/CapDsnbZGQgCmrmVOuMcG+hAIBKhSIsc+UqBr5b+VlvTo2EcuS2F8CzqOH6
D5nHybZlQ7J5u0V4WmjrbHvfQU+ver88maBvX07yXbBPqVxUCW78wdcpAD2ZBZGwsUd0Hypy0I9z
gGGPmG3du+Qn2SmT3cf+80q5/Pgj3GBeIbn6nOu2kEtIPN0FCwfmWovxx4rXHRatr2T3IMhHldRJ
Ks6bGl7Yyp/2SjeKLbc65s9zHN8uFzabavvFjdtLZ9pHJ4OPVeGwIsllMFkq2aAoD47bQs7Y7Vd4
GD45NEZmboF2hWmhOWcZpiBE4eWdl9evnhqkvzOHF1tNlxmIOF22hyefkI5Tnvf7XN0m75C+fDk7
zszSZyDa+IXPERvlq6RhGsi3dwj34B039hl2dFAzsV679M24IG+7puvojNpV9b+3K6f7zchMu3Fj
9G3gGIF/FSPGL+xfg1/w/nAcsfKiv6bkUFKwoHHkD2akZHBRC8Z1qd309kdr27UoI1+jKS+plTf+
02D23MhNmeMj5eK11fCChU1SRHVQ907jGiMDobHrK85A+flGYVMwYkeYY1FaribWASgYWArdtj2D
BQ2FO2Zzzczkq9RlolXY/XIEE4rX603hylxo1xO5NHmFXBqQRPVCl7ws5I7z+Q0sROadUgwTtxwg
BfloYm8kXykb95S0J0imb848ObCowvixcoWG5514zIjkxCc4/5OS0jmwXUqFA1ItDnblIOmUCKhQ
na/t/m54G2uFjugVg5eiRsMTevB+nr+DbH6lER4wYv7peFipDDp8OIfeeA/GTEsutpSGyih954eq
Ip6FZX268fwBspXrx8jcZIwrswQnlWOXsd2ivTPsSodwYrlHGjR4KmdMR+2MnF4fr083WkH/wkyT
cqqxmyo23Wlsa3c9lzmFFrnlFrb5LOW9bdXVpWFEJ/mQAaInSS0X/jXTCwjYqX7Y2vmema4m+e5m
H6tbgxUvUtROt3thAATLEZB6G5iaDpBLneLizur6N0MZoRMQ9Y2viuhXOv8qoe6jsOD+GHAXR7Xs
tSzXoVut/lCv63aO+7PRZG3akIlNR8miqvk8oh4v6p8Q9qaqyOW1PVjIa8qZDMIAIN40cewlMoI5
4GlzT4Bz8yYZEBpue7PSKYWg1Q3nmVfEDapYneVL+QZwv2eDMGlyPtQ1XLarFRY/AMFa0MRPyjaM
l4R2wo02kwg4f9wZtNEVR7k94MEag5XmncpMO9wGuDbAIu7uEovMn36eBo8BGOM8NzpZI8DgQkGP
VCXETebG2HoI8P0ZvrCn0kIKtqJl6HXKPTbi+mWUSZeLSu4kLQl58bcCl2JyxcgWFd3WSuGLATF+
gmJSKaituOhmuLSZZA4xuQZzDRbfmyWGwyP8oE1lNiDStFV6CNf1KqhLT2Wy/d3ZdgSVZ3mCeO/2
RZnC+pjypc22F9bEBQAq0xFRZR0lSmcZQnLDneJ3ZxBz6JqAEoOh1gWrbfw4Jy8+i1OJqsNmp1G9
7PgTuGrW8QNlq5ZHK5ad2lsWxrF2BMOEf/p8ufR2gQZjnV7YTUl5gCITgR0hDeViiSFGMuOjUt2j
/MvT2dr4mKJZjf6tuvnfsC2Wb+bzO/4f4eDW0rJ5pBtm5tGL3gwxQ0dHtbwLmbBc8lzD20IU/9B5
oNELaSevb1VC1fbotMLSJpUXSOZJBZM3D2U8BkXIKUDeDUzm4ussfP9AjZSxTxyTHcp0yWrBX3z1
s0RH2JmyPgzOFaFuksiAO7tNvzTll2X379wTXb9IxxDhCNHNP6peqmyVBj+iHnTYl1cGUxXRN22/
3+CojE0WpGXX179sL06/cjlLFX+8k8HM9i2+YZAzVST6lTD1nhV/lE0rq/MXorGDl+FNht8rdfL9
HcetklA9Myqj1Ug9C/ZurLK4LGUgm8WRsHwcjRegbmeYFrB9SSoVWuHZ+25b3khUYP3nZyw1huRv
Mt5KuFp2MxTjY4ncoA+YMT3lgKHtecxBLc7qGTOx+ieCMpV4BBU42wl0EzfLipBEJzI1gvphqmF7
fUKs9bJuLQFUkwIk6BrFORQWt00Gaeq1VJyjgEfTMQgUWNmmNj24HqsJpnKFWlo+DP7utcxQepd3
8K9DgqjdXDnLSiuKIsIY4sMOQocEAGvcekw9KEBNw5zlqSnYaeFvEoYrYm8GQ3bh4xqaXF9Xg/y1
3hgd4NNsDaFueYUPyJ0KukZ/w5dR46cjMxa3KFxnQvx2iEoKHgw8kYVs7kKz7f7u/fXques2FRn9
q3P8jWW7qqjtDbCP2LrLKfFNIE3hr5C4T9bIJ/Ww/c2rx2Fn/FIX8zO6CwLhY5sK/DGYJYCqFUXS
jT1aREFamtHOorRIp6jcyyFibcgIkPT/y6Zu0s71h6o8fnjQJdUIo3eRXZrM8qqkNBTSmiStxJiL
0W+Z/1MLEfW2dRV2U1eW97jYKopRvw37lqyirz18/lhYFBnOiRySc+jU47qiv1T59+MfIGL0Ngwn
O41p4cIa4pMN5cPscYOXqXeSVLrZypq6WazNttojp6LTRH4X6nkUDHSd97nOFDe4SnOwtcgkgRg4
w0312Ub1tFotDEJ1lNB6CNq3w8raESQoj0I11grjUDgwSpDg1834pw+V4eTH5Djj9O+PtBTORETI
3zKykakOwu380ut67/3iuyYMl2xACpWYZ+Y8UOQpg5X5Jmo5C1zO3RFG5r2c9CGJ/F7ra3ez/NN3
1zJBvCrZIpy+e8vNm6vdIxEe+1K2+OSPp+sDxzQIJFIkHQJk2qKmpHVv+gtpONRUKiUDV60lKVYr
LOUURlO6PrbuA/To7dkol22PXw8lWlq6tQ4OECkmyPmxPS3m795njXMy2GVJhJkdOOIcJNabbv96
ISdaSaoryf9cz+l680dCubgk8P/gwrS2oNdqjQjtHGSZLqEz3Kx7RlJ8H7pGg4GbHDRRq+G2zePm
ecy8auIPv1S2YDb0Arqkw5EGkZzLkIap0g5J4VrOC3yf+6dkoBdlcXN76pylCfP6jlrpcYtgHapM
syo/tnoh5ZeHQlI57ngAWG/+2G8IqhjMjBUdioawBliKKS7eFyVpqSkTQ/rGwWqAf944iMUkqVw5
POCAAfFdHAFcKh065w6oxCz6f7N+RRa9vFdRkt1bIcoHrA0w1nPcUag8SNJqwPbShR2H/qXDyAYa
RjDkkIVjwkrJlm7KB1lnAjm30oWr6AitBl+paC0c3mtGP+OddnJV86KU5Hn0xncxk5arhUJBMK1Q
xWYETdkOYoKvLZeqgp+ogJL8feJmKVc8I1L6XMCKRF3DBfmPPpXzKzWPG/wJHZVX8YkWOz0OlAhl
+v4uDJQ26VYVemypNwGGW7Ud+F+C69eVHJiXpaxmegkqSKc4Bt81vsej7Yq+6TKkZoXGaXxHjwo1
7YIKW7Qb04yxCmMEy8gDX9xyiXShqidoR/iyTwiieCoIFItbRXYnpbWD2gALM8Au+Tlw0ce2K4mQ
bwR2ew7XdGDeG5l24V6ZJEUOkExBD6fu/VLn1lYhsredGPeSGOhreN6SM2P83JIC/CxpO4VyFyl4
zzA02x0H1pjiIuXGhFH9sQCUse+zM5QQ4fdNFW8SZd+mlfUx122w2VguVqsg+F+QI2Og5y0n9cDb
nGKpIle5w3daCtQBglL0M/jk/EMGos8eeDaysPbYLP5AKzhBo8jWxzoH3n02Cxi24WoNBzOfrP4z
cs9CKg9pFMhB1XZy3phNlnnJgQOkeJLlUlCasQEbomey91Zu2hRiMs3xMKay7Rs4KqmamB634RGS
4BXCjosXlZatUYfqE1iT+h3KtsbIyNikFu3SHdR+cRMq6GrTrrHo4qmAPwdfiRfHrhUEE5DZ1z2u
3lCPn+Nms9siJls1WPuZEl6Xd9qdbZ0io8Wfc1D+L+tqleXc3cuC7ag9MXF8fHuucQG0aLslpOaV
QZ4Fqjk2ec33iPZfLgrQG7dffYTvPDKfnKT1eVGt/8aqTiDxA4sBOUzcbg7266McPXB0ITWIziA7
Yx6JhIf4gDOoXN8rK371IzBINvaoLRuFjirhipGkvBrbEJuDUYPkghl077lKyBMpl/dLxMzRglo9
LFHQknw4F5UO/e8OMvGfOceXXz1Bpkfb1LylDmpcI7cdw3scpPgldQKw/scheR7i6bZEbU0fPhOu
MDiZdR/JWoFhpBVXYn6UCjQJvHNMO5yVgx3OkjwCzBaamDXOKJwmQaNp92uh+PS4e2yCuDXgbuaZ
UYqOV2Il8qXeJSLJfciJtQpWdmG6NQuhJHSYTnnn+nQLfi8HqUHFW56O6QOrqSK9g6es8cou9wH3
hUvMf9pxJ9/RRSY0/RSHIxJhq51kUwg5IFyA6AjBpYVU23j8q5AlwsvRoekJ2qbAKbiTFok2GJ3e
QtkO6akP7dcKQuiOLArdAaRVlvcEXFVjWHNHY5NwEBcsLQX4BPnfnLq2qcR2rhOIjV59L6w963MT
lXHu9AIjovgUrCY79sTZw0UrXdOxNtIdJEQ5HZkx32KXTYz27BHzD9qEaNjtHUaPW+TTb+WU/LuC
cgv4O09HhwnLo+H/8b+Hg7CCWTz+EwxCG3SGpC5xtQxHYJHNUJAe2PH4VO2V50jdLH7HBC8urNZP
e4w6R5MICNhmo+UG90T0R+Gh4GZxMTvYhD+uUTTjxgLtBFBrdsAz/VsD6zw2N9aZCwMWoSj5CKfB
zEp/WDAF9U/8+44e4T4aep87giWcLGPyQ1EiHh4+CRCgCLJIfFOliYZ8H5Y40Dkuuw+iEfMly3DU
ZoRhSHEnXdJabe0kQp92pK4Vi4z8T0jXG9v2HhxqXI/a8gJdeG3oqcxLhvIirXp/szi8qBouQ/Tc
1z4Nx0uyozMtWsWBOvZsvzJ6Rxy8fKah98m1nCxcERvskS0VCc0fLioXaVVHLUfD27H8bJ1kuzR3
W9tSF1Sb3weKr4ACuBIoFWvmznIdcxN1DO0rjws+0G06WsS2hOPvmZBVKTGivDzG9cDd8XVttiH6
H1EhZkqEEU89BTKNpNFzVYr5EucaRKKh3SOMINaoAN9q2NHiNuPhwf42qu+cB/u/Qz6oBrzk4qwq
TWASEYud7IUV8gKlTNeIzplGBW1nlVB3wAjDpl9lRwpPY7nssgNbUZtjLRSZeiNKRLyaUD9NU29P
88yCl94Vw8P/39W/C0+k6XZImGbgtKVAhui9o1xzhb0d79+7N8jpNrVvaesAf2/WrCIVOjcWGlZt
iNJAwY7zo9PO5Nt0N6YBUsyxfHjJhpiACexe6uybSMfAgEqL+zCP1R0WEn74hUI0MAR9jBY5WZ4V
Vyg2lFR0TfgetAh6Yedd7142viqa3NuPVHBA9MvOUe2FYImWv+N62wOEcQTT9zw3QDCCUUtqP5z4
knaSeYoH7eV39SdoPdABtVggpmVhIyyOxdro5jUKNIYt5kT6v1c7bkSzUOAq2Xmsk1Lr4m/056L1
Wvs209n/eIS8snpNln2N9U7JsZyIJn1GvIdBq2TF6Xf+CfXQwjuBLXxF0wj+7FjhfxH1bA8/svgW
OtMwiskm+GeXBno8iFSwDJWwtItxVNmzaYepwZTT6Kb2HTMUyRuJismhxRLP37NMvV9DcDeDnCCQ
hNdPaGBMoUzTUISdxlEfQUKWyyWM/6c5QU2XAiZD5djweLita89SCVUnUOjs7/lV5lrXYijSCDUp
K1wSjyicbzWie83IKgd5plZFh3OvYXemxdCFtrnIl0Kry0rH4DOCCjpJuFfa67k/RhEb3bpevymO
EswP+ACDwfA0DaNMvSDbptRLAicZNC4ddzsnBw8prIduZDPQAEHNVe8TjNaZfQ6gLmpjQJkdKXdL
3jr5ByqALV2kdHdJ4zLJ68hi3535fF352euhERGM15A0JiKbr2CZ7u9weTs7hZ2NYhJP/HNrQfPU
gw+Exxlt1z8smHuc0maTVw62eZZ5rm+XXFzOYCFnxTyq83/YIXja9BntMofL+WSaaTG32l2bx3zq
4u2doysXIVmdgVQQyy2MneqdjerheO6ekx8aRHE+klG81jaVwnKF92x+hOC79LC/z+Yo7IOiVDfm
Cc9ES/AzE+MKeUNKcoLvv4ap793uEEjaGLsCQBzl29fFPz65w6woo06QGgayijNUCZdZFrn6FDm3
O5KHC1BTAof8YqJigCtnLU7I38FuIIBzaN9HKO+N+FPhEHTRqxa/kcebjfqB45IogQy/pWprIyfJ
kCmuPXqzDoZww8xXVXm+GPC7KtZ+0JHDFvGm5L2Z0aM8KFvEDnw81Wc2Qwp06oxPsnuC6K9R6mE4
wsX3hkdS1M1D6YEhdUXzdzxHmgrt6XenLxYApXe3G5pyStTJIZG2ibjbFCMLaunC3yat+XIP272K
ZvKKXCXq0uba8BHT0FhIDoAnAqAQxzdoizJSInvnMwXAUx8JBOD3S1gFC1ntNRvT26dSE0X4aEgY
8etzlqEKspRV6gpe1Pc5TvXWnmfGDotI+R8H0IA2B7KG6mDW7FRoTQIFZhh5Wd7EP/3oUHMBfIE3
OgHZ+s+umTUQ+Ap5PPjJki6cDW+OxR/sy2BlgZGv0YQSkeC/2eUH6MNoW6z3BJ9N46fxmsE6Ktcm
mZyleEG5nC/LqpzN1471EKHQ9fM785PZvVLx6AYh/7IyXHtrfv/l88slUcpio9Of87DcEsFKSTMO
59oW+rmG9S9joC0+79JZV9VHwM5fkZxDpJDb1v3Fl7+WxLWRYGFgj1nEoxdrZ5E2S8nw56nF9vev
VE+KomXcmd7gRe7uzrPmSGptGhOCS39ORwgAdlJoeNChnmIJ5Wxg1xICx5XEXhjzt+OTdMZh0rM9
rBSUaIKXx3y2wC7RiJIrOXl9TYLfpuIJw4VTZrbRY/Hx/gJTdzZX6nrxgzn4oFLCN66PIj2JlUTg
mMwTVrYeY81QfMFv2Z+aNOx6fiC7RRwqAZUFCl2Jmggfoot5yk4BCBnRu/GFZ1pWg3y9Q1B488ub
0ObvdvetC1ifnsaDg1PuVGW7rdNeldmVz30Yzs6y+3C3YDmCAnlEV0LVfBYXGUIcK3G04iehFFHv
N6UwfXbwj0h80Uy9aNUBfRhBjDrAjYGMbWqmYzZRJOtTaBhcuWImxUJIu0i8fA6/ChNpRRDAMOlL
SVXR9qB53vR2LMq7SKV8QIOomtnCBywkfAHqzILMMi1YjTTDoD55HsGzASYOEZBsR4BBK4y3YEh5
iB0BIy/U4GppTmoqvx06w1vtZeGoxMzr/bXZfnC5CQoU44LCmCc+Td4chFmKwbg/+54jXBJcaZnB
mpm3IkfXYkrVItZEtHkRk9gM0EftPSIKxzY5zy135osRzskeE+t1JSGaVUMyQz5/pgZdgOO9UsGQ
7p7raOHCNM3zCH43ajetNijA3ETFJzAUkN3cII/DAyqaAJI5C5WSqAdtFiv9pKPC2ip+iTslA5eF
/Bgfxld7jAP7z4LpbAGZZIyXV8zXVgGTXsQOTqAO3LaDxdNtSlGdpHqfEmbbMHbkZ9fmEAgMwj9F
ZxQe0dSNL7FtHUXpNZnZh0MQYwxbzqQJ0akrNcyM8mNdNyF2pBqQvlLQyCY6QpcB+0sJWpQ3VmB+
O19ZK4gPQgu/6zLw4D5inhvsStjSFv0tpsPeJ3KtOrQYgeo2RrLc51ddGWvnOWM8uow97PmxON6N
NIR5sZiu8M1HmN7DaHSFwqtWGydZDbrOLxJ0639mdY4Iy2iYNTuHEs1XO6nPt6u5h7lak9L5vI2Q
fI8pgwPf7QN45ac33U9UCs5yVKJtYl/ZuUcgPAOMaP658KdwnooWjLskKe48cUEDQ+ovC3oGnZmD
XUSYPq11y+wLuiTLqaVRNu1Y5blvOXDy/3ANH1BW4ImReCuoD+KLJmBfA2F/DfXnUh9mOSFQI0KM
jl3c+rsnl7c2a3aVIXOhw8lmE2HnOP20Bscet2TIzL5D0kH3CPRU+/TH708XgCMU/J8Rz8ZwNgJb
c6ateHiE0b6cdWLhf4wNTOEnUwQ1i/4niGMB7n+KXd6kU0JTNvB5GctHefTQCP7NzwM8taLKxbEo
/3Pirx8GS/Cg3BLH0QRA1LyWMXKL/MahDS7CgEksIjogsv4B3JlvK4Jo8N/R/wnEKMNZrdvcNxJY
PTDPcPIQIou+dthfHTXi4eeMEUxXeWbK9LlFfaQmu70H2FBU6hZojfX1ywGKjW/3boOniVzVVenx
2XJf1RKmHRs9OVnVWwj+1hinf/4vE6qXREIxXX62Ew2++A6jSA09752S5+pCGi18whpEi0B5+M2c
S7qzEuOA0Vol4JPxva2NbxkyF3UBxQEle/ZiPX7JBNaHxmHckDa0gDSfdptHr+IeLd0ENmytPmEI
YUgp290+imAaCRGE3W7X19GLaD2zxCzqulCZLtK43KNx0qz/j76QVdi26zcaW+UwZt/iyi3aviyp
LdV3NTY8eRmUQ1g2WMZNR0tJTDotLkNhj0GDzbKn9CBCOzOPY7HVfTn2tV1UxsdRtabuANscEDGU
iSUILQ6SW7gjMVybH5RB/m1CSMGp/xRaUmrXBNxEuOMG6fwPy0bFCJffO8l3mvYK+1CGzDJ3pWdw
wPfdfdkUC8f05hUnly72ZV0E1ygxW+fx6Ttm4QhfZBbUJNsLk93LgME2TsI7SSzrIPkKRZy4y6mH
6Ss+lQDiQ4X6uWOcJlT2f+CjBF8JWW8F9+s/5JNWvqB9t25pVi6g4gXJQ88/Vn4GsjNeKMTbx304
vHUr/C7Io2NZYCu14z5Q8fDSavq+6qKlFw5FOf+WtELbM4+LRDH7EcQZrjwufbD8zz9p/8LdJxsB
aFgl/GG5Ki0ITiVFZIntz9TMXcizq19PVvouCuexjJdOYonovw+4BBjJYoun4HIN7v0S7Rs0Q07q
ZdzrxYxeFsNHyAQHM+23qtlZV5bcKcW+EO16GfgzlP6flP+MoNTnKah/lGEuSNpyKaG9rC/fRBpA
/NQtufcmzI0FkhFv583q80dq4FFu3/HnscNLfLNrv5W8tTQtu7CHfzylo3eBf0ej606mYVsXGY9W
xBfblZ329DNN4QEKLgCVFths2hhP3NtRW9AaNH+IjER2jbm9xiO+pQqOjrbp+xgL2tRamymkg3O6
eZ+XjYYN/fjn09UXmGTMDpYO3htTMJQP7kXC5b03xhYNwtUXwAxltr3C5Mh2tuzGxVvvt/4vR4g6
IbkLMw5KsjYx9YIM9amM4yF3FGwVrdOWvNHttrLA74fiKX4jDchy2f8wWbTrwfawopJHIZContTo
cI/bELC166TBMtDM33IsazU2fsRyNVvK43WkiMNS4u/ClubYlwQpHyth9fmQAfRkaGHbASnJFqpP
bJcE71n/EX/FLeySD/KSGNG1b/8SZq8jlgyvaoAOvtypFcfzZRjlTXb3H0aTzbZ9y4e6Gof3BtZV
40ttS6xJjBRmB/MiWUn38xdGNn4lPmrVQEKkNTZf4w+APWIFCmYDTVtEIzPWEp7SGmh0mIYPsbsi
YgWOLQ4zjHn0Rvc2evvMPkYkni030S7pi6x4pC4Uq8mD6OYu3vXoBuhPSmoKObjPNHB9bG//HOz3
4AXoki4M6OZEwM275RXIVs0T9foxb4kOPwVL+12I1EGxJnF+etYgrtpZ1W9ewD9ePGDcUCp2gyGZ
fZzU3wVtPH6/QHnipwcu7DOCMkw5cZEodVCAOeFkGmDxfSpWeQhElxiWqm9bRSXc1M9y2T/Pc79F
yclaFQJ5NWLO/kAjo7PDNDbYjlgvOkpwBFqyRR6R58EFZ2oRDt5CBGFWoKHnGbCm5wpDa7oIsBJO
0mvSuzIUSeCxHy+QtdpNuXYZC2vD+Flds7Ccx1DcmmIFWL5OZ7t3g04Gxw8LJy+ERLNswkZkM/Tl
YT3cCI1BtugliOPFm9meYINgDrRRE8uAXKPpXwKBt5GFDv7h0I05cqiB5l74CBxdTnGlp4+Zvlv5
L1tMYoLTHznFYR9fc77rhhmzMRUVSBWGR0kt53qRH4O2PdfGK/cewLqa5mC4qpz6AROfO7PdUlVs
5zjlwU6qVWPjJ8gy6F4bqFXYf/iQkvy1b3V1f3a0xKHZtAdp9wYEBe14zEe3ymdUHITuf1qhD4HN
NrLBwlKtnKJDpu7ZpffzTj/9JoXI/xkZsfsAVzTquDPXOl8TmY9zMlJ8HHtNCH6h0EAiRguoF5LD
HGb1Zj/9vvnuFQc5ZRD7/PaJtHAJ1r600cubQrJl53KLQnVlLEDeYDBzLCbYTWJgkpE5ss62H0re
aXHQVuc2jPQ4Tzfpt+u9+UbkJhz6kCG/QD7Z+k/QVYK09l9UZg5jFXr5fxiWaOCk9uJB0o6HdRU5
vxnYmqr0Be3WCU4CYWdFbbj496VgI9UgtubhgoSBFxQAMY918flQ6IRViavtfYVCgg2lzaAy1RX1
1vRGGnlS0jc4tSF5azLAGUjZuP0GeEMby4qRuJ9a/DNIDw2acDBo7xH49QRSgab33GK/v8pHrYn8
AHpBl52GMrpr2UxoD8XKjHD0VEmGzWbGleLR5f2vzAkjaEIOAJot5ABw6IFKCoFmI9foed1Kyvyo
Ad9F6EJ/Glo5EqkZeIUjr2RdNAXkNdDZj7XJQWjhPggGjL8TvrZtzLJP9AQH524E1Lp60RWTqbip
6rBVLy86LZu280IXKgrAVi7fs720nPeyNImHjYtTLQWC5NHvoJW44/akwve2k97qgg7a/d3+lhI/
DSlUww9Jahx7SOndqpENl36C6Q2s+AGwPC9IdVM2ZP9CRmi3LJoSJdG9yS6M8Mv3dfBE6r4d0G61
vpxN2hqQpATIWbgD0uqXtYHixxmlYfliISjXbXnO51atK3PRmFa+ET+nhVWWmxJQDwRSk4y5LG3L
+cIUrlzf6YeESIFxWSQn7XyRAy3jFS4MBeFZ/fAHFbqlnLiZLt2USzyP47CtX6tQWJJxfMNjYwkL
DayS903onJaOI70+0KQ9Cp1uZHuUUpf1LYWTiy/JbS+aKigtjmAcWTt3fTJlAUg/kJMCaMYv6RPA
5w7BXXnf4MtvznhW3AnQnPmN1J4HY5CA4vDonR+WZzgUXg3JYG6dxKXcaCm8WHzTLt/5v01CKwxE
vfAEOikFvMUkL1jzy8jPoJjRJWx39oSVQNWti11zJOLzKdiP2weQc47SdSBiN2xoOegXKEIXizlh
8bp8o39pvLkWQBU7FebX/5GWPxOipPYooKhJ7ylAH45eEzT8UP32rT4EG6paqV2Ae365AYiXQ1lj
LGw4wLDV0GgTdBK4Q3EewguvWf2HUk6ICYzoPCHJUXSIXHOlPUIcIFkcLQ/5/5uqqdDfukAy9086
A6J0o/EEpxUL5AH0VD9//XAwxRpDxLz3/rkmgmkWwD0gZqAD/pqura2EEMxWaR4//H1jUgK0moEk
jByFJhfV9ocmJ0aIDsm/3S0hvmw8eKSbsiYl2QUeqvJD80T6kU9EXlBiLk8O/xw4kGBHjWCr4DSJ
FNdi+Ta6rC81hBJcmy8QtljAtw1ySUScbLM6avh/dIfSKlgwy2/Cfr8A3k7ndBPF+Om3Ul9Evj/3
JZGxrYtVmXIg9ZHj9zh6CZmWuqfvZV4YI9SIent5vNQ7lqoW/S3ILpLCK6ZrWQeLh7ZcZ8MUlrhH
sbfJxAoII6XTefIV7O/NRiP9DpNhPtJ1+de49WcFl44eWhV7T1dTlJT1vQ1pdFZuA9eRrCdMZoIW
74ybh3vYLiIPYjc7cM3+xlhalcVx+AJ3M3ksz5wMI/wSuQg3VyEseF+EZqies5xmjCwaXrDmwYwk
FqnG3031hFr+aHusAOaDqqzTHsBvFGLQeBuUPw1w61eBaqhX/2EgAvMVXNm26tY9HGz5L4e+24pn
SljiVAblv1eCGBGThfQhmAp07RyMFVofxPJnbTcFgml2MsbsyeNVnCLz1LFCfAZFo8L5R/wfePjm
U7286RdUe4tb839ZogsPe8zzxmGRzkFcKhnQudqR5L5UU7S060xlC94FpTPWBeAvA9Ke6wQbRD6e
1q/48YGx+jZrYPHznUretPloUwSKpNtpnVCL60Rrikc/FL3DR58PnFvyOozLWn8WPkZepVGptFzG
a3Bd3Cq2LlpysALDDtnO2D+F3MnPsKsgB/f8LKEw1DMplepLNpTX5cUlb5hMTVj8TAyZa3rRPa3z
BCUCI2Mdpw/iqv0BqotLrsnGTpYx6cvEJDO1EOXOjXjKfGF9rC1Ji9+Z+pErvL6LlF91UbVsK2Ro
9enmmDBi8NgSSfzVnqQPV7ZilOChgHx+sPIvU63eXujTnQP+go8F+DNboY5Pm7oQesXE5r+tg4pM
ZFoLXY9/jDLifBRbYYyrMFCKpQtvxzfinK/Q425ibfl1y7ogJGVWRkmefFAamikZmwsDFYwKdVkJ
07SQ7ZuYgrrIVnj4ngWA0uzS8IRRmNQVkW2pGnOvQ7tmWUOXsf8hAJq231loPxPOxVpObA5zo6lC
1NbYmhyQmYiLilGeUzaGKHi3fk+lzSwhmtekSNzvNvsrp5wFEFZa2lrnGhBPwJd8gMllnMPiqsLm
Pb2XzZ/zDRUWFP+5Q6wnvpsIqFiL2iuSjvWB8OzBE2PZLRCmzeu+QHs+lYvwTJu49KBU4wm5r3QL
bHG1K7zQ6C+7Pe0aghro83SNcaKyOYQrijuvaJvneQZT0FEvj9qaf0zUPmyM7u+uA2fELno7OfuE
fqRp+C+JJvlYvBntOSz7PqL4QJP83HlC4WCyWMow1dLp+gY5Z3lpWzH0a25OrKIBTqPHppJdJkKB
etctZsysmg8r9KCUqtGFc6hSjYfP7yEvTaX+bQLULYFAKegWgyb4WHl98MYq+gqlBl8OO9wlDUya
GtB4pUM/4o6kLcsaBzJ5yM0q4zkrvVbF9WJKlwZgnbh+X2Hw+GEvFZTur+RazA9/YsNBuuGAQ45C
nXOdxzLIdlbGulUSs3qBtxfkbRPLhFQ6WeWF5tDt4Jnq9xs2SZr3x52X/aYAqTYuMDK9G598MJit
xbLcrbZFzkppAIkCITA+YaJWv9zIXdLbsgoBfrAGaii52vUE+vjJkvp7rGrCMgxqezbDK9YrY6Eg
iJKjts/SPnmsDApzSli6bVJxMO+HwU0jpW/ibQ+qACUM9okTaw5zQKrSzsqgPyIoHbM+kI27OhJz
CiUM2tGcf6VfFbaRdDnYtpBEWRPS3JbLnTa20gSO+yech39eQanf2k28j9n9xs30C06Bkv1hK9qS
iNJUM2HtMYWUWFBBpLWPKBQVWGXqKnb17BRlxfSLpDQrq5Fwejg7o8FmXEaGbaH8d9QPvZuELUJd
v4+lRDG8+riihNEqO08tRlB/Er3C3p+3iBRGt8XZSy1/JAd5S0uodNZ1LbTJifdu0dck2r1Uf8Ha
CIVT0x1rJ8iDGwYWc8ELnndpZj1oJfz9NcKs13TyK7ti4aroQlFMNGydUrtaLnPoZ7mEa5C+ras7
DT9ebOj/Nnk7OEpNhpJ/DWDl2wGp1f8hV6stVOxNUWLUjwpXfOCh0RjXQTYTqJtBEsdDlhmlwYBD
4F08baylbAiSuV64tLHFlYNS7mMJy1/ZzoiYd3HIlRXje7goGb2knV4trOvcNDFzp8Z+E42ksFZd
ZfiNNz31dYeJV1M5iym2YuxB0rForqLYcJ5RJtxkFmD2WG7sqStZft3yvRpms9ctY26rsb9xnGms
BpR44HwItMxfQ9fJxioCehbnu20Vj2YIqoVB/UBKAmRfsMMbEdDDwKXEsWtkuonLcGOsauT587S8
WRp7ePArXOxO7bMHh3OROMbh38BohV+4dpkUYlwFe4RPXjZPuksOoeyeGIa9ibLp4CHlUHpIE7K8
Dk3ApApflgF5iaOBCQFGFYs4cn65FE9S/HvjQli9m8BHgrKwLisfn0kdOKArTqMy1OF9fKl9Kyou
kwMVFF7TssheQ/6DEqLlaLa0bq27UiSq3TebhtCe+eeEHXiCXAO6blX6gq/W5OF2b9ReXJ9cGTly
3goFb3UNX05HHzQUjKT7Zn0x+W/R/MQcChh5Wwk4XP2cJDY/YehT3x5Rtx8ENOAfNBC8v5qo2cpr
JJxETA08JlJuFYNGQnzsdqfZGK1axRn0mNYXw2ozhIZ4tz+w0PSILGH4eD5ZlDe9tRh57WMY78JJ
v+47l+Il0GmU2ZmXvTOyImk87myxzICIvHQYXdOcxBBAXnRi2B1J/cx4Vf1ffsLFDs/SUGjKlJAC
pu2rhvHKGTwIaYxY5FPdNvtyGV4obTGlCgVyyK9CYVoN/En3LyJtNVorY4bY6Do3CxgWOUca0Lp1
KOvunNOJq2Y82cLMY0I/8WyJ2TFZX0Q+qHpvEJaP4XTfJgshEIZOvVbddYmmoibXBdwPChd1Yni8
esDw9SF0qbdiYWRh+6Mpyfolt+T5wUNRkAb1Lr+u8OmfuNLqbCcPTyOXbWmAWUa07hRMIxP0n+jc
W7m0QYXb5GiVe5htSrtDRgbiWyCrDYP9iZ0kq4941JH5NTENqb5d/AgjS/j0qpQ0IcVVu2gWfYQr
TJFd1ckzDtfoz68NJBqtjKroP1c3SVi1HwrAkGw8lrDKDVvQmTEx8fWvympnvbx5mTbn8Q13GgaT
1WRC781HitpMkwEy7FdgJRvgq2Si13/uoeGCqhcpuHx2WNKICuBe/0Q/byK9Vz+clndqjAru1dlf
QINTMHqJQIHisGCaDGoPqLcph9nq7PsTgHBv55qVvgfqo3wh1drpuBVGrLKZQ5Zy5BSWKjdyyfkt
mxy744t88YNYz1K+uan4P3gmIQGJ9vtXcAENNQ2X/D/zuRSmSLnNAd3H9aHnuyZawDDqXHCNk+dc
6NS/o0p1sisZmRPtJ6TdaPt1Quk4+6jAUHFAxbf2b04cu/JPK23TN9w7NfmpDLy5VxfEmUF3Jvu9
K91dBH4vWe92XYC4ocaBX2MRHvUUN4rEMpyGVhu98Yln0dqWB1zQ7PMvqmjJ2/1citxsxOc8mP3T
chklp9WYA6pQuxRuhWcpYZkik7x2zmLQBVl7Ee2v9arZvFJJF1OSJDQl4RVPcC7ug2RFG4u1TMaP
OqmRBRcZ8ZIzWTHBCnatzd1sQTmqxAhmXlsJsikLdzuHrAy9smSZ8YXB0EeX9LQxtPDo8memyRgT
8x2DThCyMrWmtQOjzLQHRM3u1iEiyqmBnE5lPJN/B5rd3QHaPetFp0bEgdkNetGJQmV/AMGrVjZN
YZuQ3hN0/Zg1NotH5XsanHldoKCcjzYOBz83eOLVAE4BMOiAYphktydqu2sVPKCSs1CWEota4Jwl
Aeh22uPl0uDnPSMnYDW3Z4PWtbR3lK5ffB0oY1CB3St27gdeHJ1mpIJpbrR9GxTSl28F+VKklGI8
Y7iRm1DnpZrKLTOHIvYBASxCVrN9k/yxGjnHzyPiu/Z1NDq+DcasOUlmpm3Ogkt8aV+xl0UI/zok
jXXj6LJ7m52zSgOpjBBvr5+e1tYrITuFKMuAe4Db8iPEx/Q9/tpr7ZX0UP1R0OKweYwwh3T4TOHj
z6EtUwvF14rkZ/JEjlEtL3nGtCtwVohEF2H6pyshi1eb3xOGBTheKoCnFvsHTWFlU+tiZgsMB0Fl
WrOQzxgJ8GwXcxoJhrDcLomZ9+sXOWqAjFYfJlok6Js6KbsajvDn0HuKiwCFMM6HPV/CU2iCO9b6
c/9hFjD6j0BNIz1FFd2sdjTfMzrbufy/VuZKThr84i5Xzz+t1gPCB2V1c6MkjJoiSQ9hNoTmY+qi
L2R/W7Mx7n7ZLFSxHkEMTd387SViAvC1SQFhrZIJoTbIshsD2qgjPwrrB8BaxOmDhDWqQFdIo7vb
IU4Pwb/QgJQhIKX1OHvt7/0M5VARNsO09Uw4PeEvk1ugoBqz/iy4vDEmgX7t90lwhQc+rJ3WxwiV
KH8Y+m7jsnWpcMrL7iLJdSLQJVozo/TrtrWeqzQLsG+ONAt8BOPxzhY4WfcMeAMx7dralkCVGpb5
XUyAzezyQO+nSx2mVb2AOi/6QdZGn3TylBb+LUFo7m3cb61JIPOZVviRJYSl2PUF/F+wRVm0igtP
TEUmNq2BOQH/dS93m63eBOk0GZ++YwqnndSC8l9pjmfr5gGPhobiXELfaDeVhPk5lu+GPkmJLQEf
hwoPpNJ16we4vZKBmu/VJaJuhwEwn0n80R6uCuv0pwOlViOlNXTZz8EBXFaDZT0QuV8ptZZyWPG+
40mHBLC0teGpFXMCxpFCT/xZby7LlBjzO7QHM6OtprqdJ18/vp/PNrojbUltOg4QsR6IFLEm+Fk4
RHhAxYByZiMRA0GwsnVIfALa0AnLln4WWmnvE3McxcVlhLL7LWApeiOi7Kvh40JUm6dVzp70F6zL
XEossq4njB0Z+eoJu8OyYcqNledP4bQJC5P9jC6GpDytk6VteggExXRMjGjL7bQp91rqFw58XPct
IMcdpjkK372oKphePCYH8TKrM+T3sFi2kl5hQuxG386XrdUEY8kPWEPpl04BsFhvHNjJzKI7IsBo
cSvFtpcisMvbGbde/tebHUsu+x4H1Kd4IZt0eQVzf2KurJhU+cTWwLQlvRsCHJxuM4zWt6QTNN9f
8gExw0sfRgOXXzocdfv+d3cy+bGiPFDkNwTMYtz3CTmdKmiu6LoVRtRKh5oeW6rfvblXkDztgj4W
0S0tyHrYhPsOCkmYLiG1NZvgaXSBha06rHUApNac1eXedumlmgUqbs3nHUObDwZ7cH1PGzdx6nNg
BTbEmHuGstQmWQjVuQesztFN4quZk59YL8YKpIo5/8vnhrCNgm86HT3cpF3Hk0BFpjPlqWujLTS2
JwQgsMqalEuUXH8dBL1WOnIebLDXnbapN5jCRVulKZjMgVHOOQs6Apn9bnFYZVwshicCnSq+7CYa
IWm21FtpWqtGosgOIfTj2G/AeaxGIc+/x6TZmBcqWBWUiw2SYal5dURjtox/kcanKcSBr1Edn5wk
JvFnGkjRn2iKE1OOmuXnNBm6PvMG31UQS+41z4JfnApIspzw5Y076cWtaZfOS6bM/FF1yNptKYPx
AYWFMug5fUSjWD7HhxGWTtIdpptbo5wW18RNIsDCGF2E3r6MPm2A6OrTNhWNMtJwBQYNF7MCush+
yJGKO3cRCkiBnkXpnR6pSdzOPGrYltAVXykpjHRnYV5kT2oTvuFw0cgUgvqIh1lLNjvQrGMxx+BF
Xd2TzuRrFD2vLzzUK0CVVDEzGAPhrksPY6k6oEuqaywWyTri+2Ei8H8/o8AYBDWd6R/QUjj2lqzZ
dpvtsIX8k2hHYsRMp2epKlQAsnXlpC4EUplhLD5qHAgxDboeU/Vcqw3SAOkI22kfghOcpH7o61wV
nJ+/9mF565wIcrlAFYmWNtsuUtSuq8z3qTyonIreibQOnuhw/QS2wdRdlhtyY8m9eatmhgQGVC7P
QYAAFWXlcCHTB5Hl+17aGlOqb/xmOYEoBVxzoorSd/mbLxAzsBdK0DCjBCYgaGDEf1mHG+VZtmop
ol6W6tAqfbSs79b2vW1QRJZ5bxI4lcqgCI6AV7Ee3XEtPxhYvCr06DDUnzOkK3l8ClwLQx4rgcz0
a5RNP++Qmg8V9eciq24d1AaEessJ1mLoMnnJ+MsshT/u7lTVY3uYoXnneqv/XCYMzPNGP2IT0gW9
cu8NwNEpHDGk5HfQv23l7vM+xOqT71KEOV9Gx+ZN6yj/HcT2Hj2CgbIxRsSoYr3O/WvTZ4gUrDyt
hzwHQYxELei8nalOIUyDjYFqi5Dhg2N/6iDXlCdZXtqwXZi1D1A7CaevpFPNyUeNeSJ7sTb62inC
wu9mCBGGc30ZMR3eeK3PTAhECrO+Iv+F2+p0JVBcYn4+P/tMBAVWnNMzjQN0jI3ktOsxjc8POtL5
HMfEToiUvuEG0tdFkOygw81JYnqP91Uy4FzRG+IYQdG778gexX1/ASwiPJsecEp6V2D/zCQ/PAaK
fVCep9d7TbUL+I8GjY20x0BOQT2e6Xjmmbki/qJpdrUpIl/7E2RZgeNToUAjCquAUFhMUsj6T3qC
IoNMEKDwGvOqyKhF347oXPpctLYagEIAbrZK2ZQAVbxRUAQJO7hRsSHCRwV9KozNLSsS4aNQBZvx
qQwS0nmsS30Vz7POTcHBjLuqIbvrlRr2VBiygSXlUY4ANjYS2c40rmJ+RIaSdTuQoUNZG+Iv7bZq
6lLj/eBM2HpthAk92ZOmwsMMrL2IiiSHIRIJd062PdAoV6QVtkao9JyONjSzX4HHKy2WMFlmPwbq
BmPk3E9a+e8sqn19obc6EsE74zNjVV4o6laDnVHzp83ysRDFq9q0qDYmotgHCsApjQMcJb81Ks7O
q9iKBzBtS7saNpwApvIujPgTqQ9Pm0usGWNMlo2nyd3Bhz+2wjWkMlFWOwdDuqIyJOOnCk2ibRJ4
w5Ysq09361hDSPUoATJYDHkdtQWOizReLG9TP9Y/N7YqpCoEgrzot1Gss69+/MOFOK0d69iTwLAY
FQoRZX034OitE+eVpKz0A8XQUWCgKFen5gVrvBAE34X/mMqm7uwzgexTDRzfA5mh54z8QRkXDz+c
2WNuBVpDJsvEAybkQ1nU3Qqj/hVJD1s1j1iWHYEprc+gE8s0XSooox4JEMJqOQ80sFbHNkzp8zef
+G3YzFBFIIQOa3SMoG2rkEbOcqqZua3PV/Vn+3XlNfWWyFzegLzKgGBAt9Yj78QQxQpv9hC8WHtq
Af/wncXIRzQh+Gns0N2Ia9ZhxO00ytuv55G/o2Sj7VWn5gPfBHxv82r8E7gbxcJHnUNAKAyK5Hbt
Dy79LuCwUX+cWOYR2O3iNPMjYRHvr51aSl2e3V68ECnXNH9fT6UawhXIIlsXDjM4XGLcB4sFqWS2
d+o+U4bJ7hJhTC6zO+yOZgPLB7mWRTkktDqaO/+Uv88xyJi9dDsZqX2IKPYxYhn8F2wLxXvZKVgc
cKLY9I/D6pU2hrepUJ1RADsjbgIAe7rTkJcpVjQY5OJAMifKvx+OxTSKp5LMKKY9zUtAtZdHcYcz
vv0ysyp27b9OLM5rSCRmvf/NJUbTx0IyFWyy/zu8dE6CaDeHvyPmb6hUUP6Z3GLr3EhT8B3ggBhq
0AbY7fdnyCajx34p5uu3j0xiahU/4Njw/YYtttSesvjIA5gtbmMLabita3C7Mg0cFgLAPIuJ1cLX
+Gw6+h3oFwkT26TOvJtPsvVTFZlBjux3gDN3fsp5YRiFbFieuzljpVzvQ4SmJmmYGHj2uMA6iabC
XR040E5EGuPNkV0u487i1ofhNw+9UBJRLhwrdz0yq0ZeW9Gw/MlgpMZyNvwqM/vQ0MvYa6NBMus8
yfcsitkvPjD/XXZf2Z2OZ3eC6bkh1fHtzUe4cH/XhJJrR+2c/NKtHfueovy+YkmlGZlSoEGp4Pqc
ipFsyqcdCWrimILsLUyvtQnBllmTFtibMYEWqEOlYahC0GBRBPZf+HDwrKgwtnju2VUbB/tLll2G
QyBtZC3of1BRxPoHkaRAFoVLPS3tK/gexd+reB55ze8uBqrXauhyzUQUwifK5/vDJBAHmRl/vQBB
4Rl5eVtE/GEi51X+94gHtCjfadNufWTZFzIpcGSN1HkBm2yUVQRDp0XBmCTiRSZs05aWEx5/+pDr
7ZbUXha6TJcnT/xpvDVM03TLBMNal+qB4He/MY/qq/KDro/ngO8RGngv4MAkQU+nZVHL9mKb1Cv/
SsS1KDlduYMEIPQmuZxMuaqTrfiGfeUP7x3q5A9AH5VALZrhq08Kt7TODxJHAeDORAYDy0WJ7C6w
a4wl2cHOXQs83lLOjZOI2RXtD6b2AhLyO077qUTKvj8sJXc/SkXAi/TkjladGTML71RJ+zgzrA4s
2HJX/fEZBnAeyY9msrKWonkNEl3oee9jjT0mts1dFlyxSSkimKEiafIcHWuwi2dtAm/tIt7YekQS
oy1TmA5+vFStABd/K/X8VknAr9wzGi6tNCw9051fxsVocds7eb7NJYsmg0vCMA1dQUutmfE60IEV
P8zrevI/eznIvv3N9WURtEyX617u11fafNMaFIb1iVXOI7dXxvrUTjQbj/EJ0l3kF43IP0MZsj49
DhrBYgCoALQ1/ILKs6l1hUTX9QTZwDd+zMbTU25Ry+KQ+xIsAhTX4gzfb2Sx0s1EadFTRaT++XQK
aTKM9IetL/tDPzZJBWBakYaZtFmelXO7quvs9WOXVaCtsfp9fitsJtxPDgghuxcd5ebjmvjCBV/7
0L8P5Wp7UHIYftqbmxJ3DEfJB5Y0SaltbknUtFNyp8jxsBN/vfdWSkKKUDgk2Rr6okKCSPfgaMtc
bMvph720AxMAI50gMynsYQXvu/BnwLlDTvlJVAUuG/9+Fe1tAzZveNuGxBUEFJDXETnKvP8ATF7H
GEHJJrJ6hgJQoxE48iiTKEhKBTZ4G6EzAM7sMA5OWDfSAaAK2KoT32n52h6OWkysJd+rYmSdCxm6
wLNnzQ/Foe9kGJ3bVRgwXChcrF8vl6FVu6EGSo6nrDmmy8V/EQUcBi1XRpLKF5FDAFWjJUR5KQAQ
goIdpZo9As9kT4UBGO/E5BJhIktywClHqNNQp9wzlnAlsO5UUoHzju6bVYBRlasFrN7OwojJqh+x
sX/HEWKyK2x+Qb9GFLLqexIf2IUZAH9HgFd7G/fYC84KxvH6LiS4RtFZsAnfVi/puvJT0BQI0565
xaUkas5Ol6Zg/whuPcEAVvDoJsmSjBO9/u8NsfJsg/fpgjpGhifkxpjcuY8mJgIJophlVBDD9lUv
4IE6t+xgzhyzgRTakJCxaWQh4AIOw/Aa2uEUgSksB5v9S87E8O8o2Mu8O/PcRPGE/RfjHVg0118Y
TRwddS+l7UWIDRciaKv7gfzXRNCuMLg95xKMMjxw6O3oYeRtcWpqsoREqkcvNdRnr0497oASdoGr
qN1L8TCTPxleEwyLJAUXZkCDUPJ3DTgS4uz0D+BE20joEWE64elxKXX9oUogfCztlmJ1CKlETdNU
ffnku0cE2RIXOItbm8t3syjoHt88BTgfTeErocBJWOdiYbyI4w+QdeSJxtTg7RebOrrfGB9mwKLY
fY7zssTPSKxBC+t3WU5Ww5ll12aHr+R5LLam+xUamkKLRHZ8xRM7LPL6hAqq51tetmH8jKS9MaXC
VJash/p8FWKvwCtzbE9EHoMWfnPr8hYh2AWcEBx8xEbkeODkyQsqUvD1aUZE6oT0aqTXLxyE6pZy
tWdlYqx3xtapAVRtVRjnqYg/s2IQ88UV9dU5mCgaJcDruIq/lFq2Bwu4t0yDdrntPf39T9LEil71
t/jAWQphLNAhJJh6bE44dFMNICFblymWoSULfdxOrzroKH5VjWpc5PM3PETKzS++TJxWKkM9Z8lp
djEr9cWi8JsyRMSvKfZtxPVJblq5IfN+8f4HZLCtiP0/T4ZkU5dNzi10p/79pLu1sOVwbb8Th6ZS
fOYv9jFTOwpaIi8q25hCTFAN7zZeQAoa18VnrXq5twIHhkAfvrauu0kk9DiiekkLbqZqPXG32iyF
xXaWsd0LtW1zigTP1iZnkWJPVN3tv6aNGwMTtM6H82xsZ9M8PYukFncVVeJCSV2nGXKT/0pc15j0
v8DwJkfbsZy93fcJtsRJB/ncRtzxC3E0XeXKBFjJqClcfbgxX+P2jCYGBERw8aBIwPnL/GFBWlyK
85F8zPJ0dY9RXXpx8YZIM35NpqazYdLbe7ELDQvCDdQm7KUHqZR/eQYJ8pP+sq0wpB4Y5FmlQF68
W5kGty4nYUu2iYu4jiJ1rpxioVyF5hqesYqxLRjRkUI2tnU2RJXxuh3fNzWMaKEvXoVZdNh6gy8H
EoFsuWJcxzP3M/NmFi9jMK3ZqgpHlf61KPNioSsM6GZCCHG60Lsm4Y9IU+7u1xlt09gxYTbCKuC1
ULzDCXt7+NzKQR1t4YH6y5TGdTkhTEB2hVcXWq5pVSQaFWfS+KimbTK4EztuAVEJrVMvVD9GalGm
pWJVRlkcY2DknN7817l44/JfNRkmVzZqrUtwSnsQ+vZO6nqcLOnHZqEtRAe/L2+4gzKUGyaXt0rZ
rFjLk0SRB8OYv+kyC9ZZUtdwBs9f+pIa8Is3/1MFirUbsT1q/CIYzTWYEiYA+sSHv7mDrXmqNPLD
bibfQJl6z6eMr033xP4/k5MRTHDYJPV5uoET2gJCXzCODPhgBHybd7pYZpNJXcBzqacOXl85EtPC
hjczOpKxxok2IVci0BqZ351TI7es3AEX44iHdD2Yo0Xh3fK7m3eqsU6Wnjg6FejVDiio9SdiFYJ8
YPlrUWTNcgh5qUVVTDmlw3zcvq5IU01GUbplc/I5VYi2rtK/One2zKu+K/iXrhrKGb4gc6FrO8SL
B6FkTE49TaEnIqURr4kKoUXI1Sw3QwcbSpiMv4NNaPPHtBqFC/9oCWE7SDamsukubBV/zB+p2gE+
hZuPvW7uvj9qgs9cIU2vFx0fJMAa8ZttQUwxacciOo5vFD0bMM51LR1nUYWonadxE8E3qL37pK2y
elkX11FGL/uQck0jhBFOWpRU0oKZPwSMGvm+JmSU3439Frbo7NGdmJSusvOfMQJ331WiRJzyZ9o0
azzU56g8U7AQPN8FjT0/Mk1Mw1Uf1/2yPd/UNZGjSzJbk7mEYbCdfWTL+1HZlkZCKOaST4PWWEuh
vQDr7xYtWai/EOSR1qOSG1rUVbFRd37V9WDN6S4+rCKj9vU4Frgx4tbiFQiVPvtW2eDbqy/MULrD
OXYeMU4qzZQaIJhcwRd6tDPZUB/8A9O+CWOHl84d1AfpZRX+4a6FmpoWtnwVH/FRTtEWoccDjR4Q
c3PIv9X4P8eJD70CfYHxCgXd7SNhKUigfU4yoF4YHS/KYEtdfY2Ez+PNBYLe70Tw5MyQhbe6bpKd
SE7B76+6o0h+Mq2yaLK7yWBgrtMqQlevQxw0DO6KUBrfjL2QAsy6YLuqgS5MBagVFAIpOJd7jORs
vliYVjXeUtKrntANnoZrUt+qKz+eoIz5SQxhU/z561xVRbNgQgRDP1uT6wLUNZkllSNE8y3xqV2W
qjSbvO+254dDeeusNG4qa6uMvFYXHqMy7Ms4JtPRgqoUiL/ckvjyORtJ/Le/4z52Vu3YNa8bt5r8
iu4WBKup9zcZCLT/fOR/QXRejylXpYbxCzQiacs42PZZEqDvBzgHpXzFPJtYQxTFaUzSbIw9+UqT
yay28iSzRShnTjV+zzmXNiY5iSlfiDxZ1/YbFl5QGKdgkPli+2hC2H0L1RpEnx9srqls8nxleI0p
kvuuJqGeXIkKEDhkqgp5h1yd2NCFG5bzXYwihOcmaPfe4CIYBXuzuuU6hRCUFuty4ZYcbSoR/NeB
WZ1Ca1iY7BEGZzDkO0pY21J9pcKIUj99Dnxbc045mlZYWqabFVIDWgwaLnEJHdbFo2lwBWpW4PbS
4dgxAgVTm+R9cYGwFJHVRsDqarMiU6BGoR07DSm7TGJSFUCUECM0Iq9n2VxdATa49tjffojQwsTJ
x/qkvevBAXUEXNVCLEfOo8JlO/9+e+9O7NEcCEGBNpgLuNE0HcIM2UPJ2/t9PonGCRmII3sKztfY
24oqPszyE5sok6WIqPDQIcjmZrWbAJCMOopYn4cpVzONfBCAvDxRnSUWwzMqx91FGSRMm/jAXIqO
8jdU6If5o5MMsfgAGBaJlBy/ON12NhWXi7uSEk38+1v9+gwGcUN9QR+gjO12ZG8ZXlsqGO96qHX3
5pQUCi7fI+ZkqvRnEMZwVrQ5wRn2hfhnnOq+tazr0AqqhFZ//hMQoDJPf4531GDh72R/n1Tza3Te
e7VOJ97mqsu5fOQDK6odyt/5F+xlIqeN+akN3MrvUNuQRZJ+kvr+YVmwAvyVnG/oa3uKg4LPxwt/
fZIEZuRJpAJMD22zdjh+aCZXiAiITDrEJ4ANaTSTbZTLBry57Pafhf2RGIrfOAkEZzNXYx3Qxyh6
WoTlpxDrFP0wY9hUz5goOxFkm0yPJQRbGa5+KHuXxswuB0gWLEOzPZXTH6Vql5yzqk0TUheWL67r
OlXoJRXg9j5fEGOV6FDWpzyqhKIxk9tiBli+FATlck02GjOxQMQgPDRqxJU7RP7KeuGuJSNg0thr
OjT5OlWbxNLAL2Hfjjq4XU2pxqGyUHRMy9ITF32pa3vF+r7IYfmcMw9/flsodXaeOgkg6wXO501G
UszFJSWdTYH6dkINivmtxgkoTIIzwiDMEzzVAElR5hV2zny4hqZ/aNFroDePOO/figNwBCfFCPSu
qYZJrDLbLMh4aAaci2lvvi4ur/OuoHlhDSYcqbGhgSAWo4EEjR4Ay8K6Ti+Auf2bnjqLT8SrIVmb
Lv8iL2FvnHQKDmUffKhq9elYt4c7m7tBPJvla4lT5eGphpPmFuXOKGWRZx1BjcJiveEygy9CTbbU
tDHId5xU0IsLhAGnXl7Uzn+HkGBCjiuF3FXuphz3Xo5Klj28vEXOywaziT1Kc7a3+EsMT4eQM8+Z
WCZEO4k8/a+1mM+QiRLxxOh9NovnK1dLu+XOWFhau3vlhU23eY2D0y6I0OBsJwLB6PcAOt7c5Mod
humxU4zPpjCEgxTuYW+HtUP9IPTqZiXHzi4qfFK1sZMHGqGpQ7xrV3oJUJMh8idR2pfBi6JkVLGb
6kmebc8EuAxU+6Uyjrm9OAaq3v1wGa3Lredwp+Eo0VXe6FMRw5R1fysYLTf3nN+L0u6SAqHtjPNG
Vi3p4gU+C2v45ohprh2EbiakhO8tKEC3w2F2Kvx2eD0pbfRmRGEgl6vYqp4NYWwxn7ppYtXIlkT+
YrNhtMuZujthvHvbG0EyDpUkIL/dvtFyG6ElUkm0hlSw25uWbfiAu2ZNwviHQ6EoHikfXiHJfyIM
ppq5LSfV6KPl1Cwy12KTlL2sUrbq5PUPYJSVKTTcQCpq4V7BsM9Tmnhio0uh1T1Zb9nTCiEpR2nw
i2nnobDCH2BOuBFeVSzIjK0/ggPlcG06TVBkiGQhZfEBTORppDkbwlvSdkqWNIE/gH+A+0bby+uJ
9BbfX2BqW+lkErgDgjl95+6MTHivhjsnQa0VjZgDQlZP4VdygcgNOkczP7fU/oILkD2Qif7KWR5F
+jtdLi0dlC7neCabybPL4zg9pcz8w8kVOJU793mjQnt3H80N93wZtKTpqOzSgjRxA5fPkqrniIUw
FIwWUG7t9J6Q0wEFU0B3MFX86lndAu/X/5aevr9hnk7dk+S4mhHS/DYqgNsgfWf8DU3ey5XTW6oN
r9Tkfl0TbgL1yZnW/qLBwrLmLkTWYe+zag8AdKXRc1YYBsrugHL0jdvaPRNmG44VSw4XXIjELJT6
R04EpFsumMbTNZj4MESDz4PodckT9hFp/gcclxDNoCkc3hofHyi8XwTq36v8pgFd11eNnxlP62pi
ZwjdVJ1hOk2xMlbbnpolwz8kKx1w6Q44shhAEXwoq+adQPOLvfw+jf2Qph9dnJqHycMS2ZCd1E/K
1XRf6Z/iemyymrwBW8VExK/MUksHuoVcMIKlUFAECESdZTkCqel5d2vBSVr7nfNak3gAVbkuVATQ
ZC0D/PUG1PrDy6UcSR9gxBEKAA2hOByL5sae9HGXUpLkg/1+v0vbDX5pUq5q280xq5q61X7mP2wV
Uptt0u7iwhrMVVivOh2a4uDk1EXKN4QiA7MmUPc4CM7hpHqCvsMyVZHOE+aJkFQ/71qUEgg+lSUR
tgYcHKe1NVwtDZQClQ/7X02ZfeEqkeEdYQnY1TDojjxSYCR+GtQwEhtY5V47VseLZ/zNCq3aK8lO
cFujOXmDdQJX/MpuvBlo6AL0P0Q3ziak652gdcZWPDb4BE39ksOiEY8+bGFT1CE8nKjoeLw7SAEY
e4UdyZvTj5oPD/NtY+W4sR4ko+fERlNH6pQgzkNXUjEJgV3NvesB+tLqDchiGyRLoOsKAKxHdRCD
5IpeyCE7AnSidtbp4laPpsu1yIej2X2rTjgtuGppqVa3dM6rd066F4vEqhXNMO9G5p5P+hPdSoR8
845i9XPSJfBdSSnwvyjn570XkFG6o2FmDq+2ojJ2KeXl9d07gbxfHRWr50PHItdnpje3YEyJb31i
CDhmlmd6EOL8kRCeJjg1XcgTqPyugpcJ1ZgRoMhz1gf9Rp3Xs2DXDckwdNpXhYZoJSA6jvWEBUIG
p8S8UcUxkiFMsya1KInoq5efBGYnl3wDaUv5iNFLCvqwqliiBf5T4bAgpFSjnwgqTh44/UmMtcwE
onPL5ZaZQIyKzQcbjBzYW4DrODlF1DyoL4NgEn5f3uDPztstk0bbYhInIf26o7X9BDwipeBc2rFI
J7uiuSU5AbZ7NqYy/QO4b86GtQHQxy2/KCetq/X9xMDiL+2fY/yF0wHRxGs37085VdYJsj4fXwRV
Y3N9JZPiQoouL5786Wyt/1vU1E3PxuEPk5NlXN4mAf529d3ciOU8wdZWyYcc/zrf3VzI9Ez5O48g
1egaeNvSGcaR5ilXpKFR0qjqBw7zWeGDKWAicIo/puuTroyK6LHUaHujLv1IFXj12zNH3uccmkQe
d+calV6dMObyXzdZHpYxg2Lfno3BUjWpl1sdf91a0G5D5q79d16hxY2Fr3BngQc0zGHe+kN5itfA
KihFef9grRBpEl4FNUYKNkZp2duEzftGA7zBMLrg8Sfltcgmt6q7hIPxx6QSi/cNJGCQMYMOw0GY
4m8k2hcxBPeP9hTPnDZgKD7fBhjB1bbUrWYwjDeSzahEc522D7J/8NJtnoUdxQjVf1ZbppaRGnIB
PqyL14wsBYcPxWMHdm+mgA1FB/YbJNfTU8WqH6P6xCqU6nFYqJ2LVXkrx+ryFjlFFwZxfWcdQqO3
tRjRaROtL7y2THvoQa7HUofgBhUGbTd4b0kpVVjO66pKuniqgoUxz5vo5b0m18MmK0fLcPEFPIO7
7fJ8w8C/2E44WY2fFappXpyHe+m4rEEEjNiNKBHkUYoPoM9y1yzj+YT1VrZFUs5z1FbMWuVFxSSt
ZrBwVvQwUaTTZhQ4lO4id95kZlt9sjSaMZP2vea3SjXBmmsv/Ked1vCOTblZlUwwAzKyQ9p0e6VQ
QN7CWVj47q24naT1XjlVjjCvMbgXLzTmDumf0Q0N4UJGquHXZZgHndPV6aSdvDcGebrnWZOL7OFJ
a6vH5hXSpSE8WWHcpPKUyesvifhKi+r+fm+f7YoBueA9/hPg5g88FF/Y68qWyNdglCkBofo5RJtN
rplpd0M5Jw/b9xgEuKl/DPMpVUM0a6e4uQ8VkIsDGskpLRTW4i+r4PbwEpaDdFA3mOW0GbJJQYys
MOWYV/apFKN1NjSsWJuqqJGL/Fe5zqgR/jT0seZrXAzNO3z8nWDOpIuF+w8U0krBx2iBVHJ6KP1x
WOQxnFX8sUyjsZ9b46rjC3j8AHELZYlS/auD4yfhq5EwH9ItzRitC4cntR9m410iH1e74y47v501
fYTycuUbofTk3wNBCDgbPbXHDvvLF420EVEYQYImh7fOTQfLabZz9LlxB7qfOTUatMrMCeQpHC6k
nLtkxfuUA2u1/XGW94NgEc8NUUy4fRSkYgXFOqfCyqxPIWM4wcti6aO9dMZqddoHvWjXLBoBipxu
XgB2JgmeM0O3muPXhdtk8CcRi7R+NX9W7krnFEx6IEc2Zuf46Q/ol/dSbGAWaaqKd5XLwbvv9txH
B0ny2PiRzu3DNv3KbpXD/bCFqal2tc7Mx/n2PrnTxY/ahV11gvfxbb3zhglf6mfm/sceTRaF7vZA
fv1GM3HYGhPWpBjog55Hdh4eAQLFJieHpKt5cmDAnMv4a1ui1cncgP78OgHBU7OCI+BlL3zzuwa3
ZB2CAJvCu8kq07DR6Br5XJy+9ql82+rbVx+pscGqtp9YP1evF+RMXuCQfxUXgH3G23H50JvvaEkB
fJ0GOd2RzO4GNLq0jkQ2gmE0/ObPAIIxKk7LtOgasl89zbaKXAxLn8KzSj/oW8umyY0SF2NGFJOB
kCa11Uf+vgCLJQZx+vubRNhpXNOVZ1vs8TQW6oWmeJCYUBgV3KDegtbPuLmdfzCVsHViicbKYXgM
ecMhi2Qx8QgJN+pWWz9TvgaPsxtTkPGTfdCWUUC61QlwDPNuQarFa3RQsX12ZixXbGDwoUD2lnfv
iLphHjoW8SVqZN+Px3TB2kxMu3gJMDDuj/RdaN8HZBnSKENWYX3IcVzu2d7vORLH6676AG1HK7q0
GI42Jy2gzG/EyU6lXsr+N0N+w62jK8BTx/OtUm+Pq5TzyzyQ92KEXlW3ECov7FAOu8i97k6mTmu0
oBXl/rnGuzAjzvmEV/BhYOvF7c4Ur4ND/KHc4nzw53gnTBmzFXjPkeyP3tS8ZzBB5cm60un3d1dE
KUqaC5N261StBqOWsLRHwYTiJpNM0/ECvlen7Pi3JiHrMZbhDAlNQSBS2+MXERz4xgK8iUoW1Cun
xk++pPwJws4Eunq2oy0JH0AYKit+sD/R7Fb3YAPiYOVJuLxrUZtiHFk5lPOQY0Hf0PE2dEXxKYir
Go0A8vVLIM67/JnuCA/Uog3JSyZ86A56p0mw0Asw4tMUvHDBrwDYpav8sPmi02XW+Ge/TLAuOU1G
3vynQW7BiNix4+VYLsnv+ZEc0KxFaMZyIUJxFeSXY68FljPy+bwgWL6WF7fwKU4ZGj6uMrS88wf6
+vh0Zg1b4K7JeNAQfngBEk++vbz2LX88jfxypKTMy3hhHykBOIH5Kgp2pl+W1cJqZ1gxvx3Xc0/w
Ou0cCjedrPRiMptjZ4OmhPNmoKZg6mG5PO/3e5rRLFEETAFafJDcGg5mrDmi6EilSKIJdRdFpXNI
METkyRfgNM5JCxFyStgCAcmzEwQnKWFUwqmqz8TzKrUILZVwIYw7ht0KPb5kQ04dFbyw2BsmIxBq
hnBwU6zhguTN6+vEPyeNCxjeFC7BZ9gvCLg1N2g7KrRY0VsRCh6ctiK/kOqvpSp5E0gmW6iFweGK
zsvWvXKRu20cde1Q/K+T1wZO4lzq/x3gi9o/oamozbtgQI5uGFhvtPj4Y5R250YkcQ7cOZjJ5fYo
ADI0+xT5oFwjHXvqVtsF4ZmeBy/tqcTBnNqvzi55x4OD4sqJDCw8aYnMleo7J95l8MWxFQ4lK5TH
ms4EJx+Izlw3AcdARrLNON4gdqjTWbyR55X/dsWehD78f9JJECYTzeYNLhiwoWRNsvDCAk6GCTuD
vLunp6/ukgkcrTZFZyqdjJVHtrA83N1fr81AeepgIwlSWCfZ1C5VqIoYl54IirbCypCs+SL/KgFe
wLvfsw3QHlFd7lpnyPdKBNHxLpgMOoTPohnn4hSpg6+bKPBQ8oNiQBVMqC/cXP68Ij+TLzaPAYHg
gjreq5xVz59Ds22yg53it+Dqk6CFzR4cYsOjgu7hd6T274yFd8cwy+4v+BmrlnD++PafaeN5350t
jdWngvqEfFB5olzOVgd8dCCCj6gaZFskkE/Px+w8yViHjmQtYmDShXTQbcwPIpaxYEAcvErfgi9+
s0uI2iR81lJZM32E/bocaZagxP+nSh+Fp6NC2muO6JTXL0KEgjlKs1kWS6y8oywEsH9jfBNjuDcz
QRXSzwQDYAcBqb2ueLdP3mvWHmKNkC4DF4/KmzCABjqGu8YcRMdT8B4wLvsd/wyAG67g07mou0WH
oe9sBSpLfmujkjNuCRS7aaayezeXZEW2CEYdIXFxcUD3SN3iYUdnfUCK82DA+T8TpzCQE4XvdhqU
l+PVL+HR1DbhY2ZzDkfOdz7DXHujverTYIYzgw7D8AtoC7qUKwh5+T6kSEjqTJ3PgEoEfnaAb2E7
D9DrKT0o4X/5MVvR+CFtRUdYwmoq3uEfs/eAZGFT/UXbb4SCuXc9FquUuF/UPRkE7H9U1z9536/b
lXWfn0Jkpri1EQoi3w+JCHyoMn4TADecX8bWKcXs5lClPbST8KKrOa6vuuTDWa+TJfLevu96t3R+
oWUTxMK55gFcAUutl5UzVV3Mi3N89P5zWqnv8nDVg6ufXG16g/f6YcmHGHLdYXXdi0UNKEUoSVBI
uYBCbiUo6btyFiDO9xBYYZURh1fcmq1seLSU34Hdl/SKNFWhuwYbuY7OyX3v9x25Rs7wxyipLLip
v6F1UYmDAtyQIEMCvbUyglIO+SNbtIBYE6cN8eSOirsk7nzvMRuaWAi1QNhg3qdzOY8DamApbcLS
ID1uVhUmvosVrv2GaD4zVbrcPanvwAL6iJGgdRLpBYMGKsZe6On0WF89Mpg5h5ASBZmvlcOHvLop
BjJvscVYhQy6VVpJ0vgap4ekSiusYRg6jDIcpO+121wGmc74FIvReCtQkk2DrdhUXuTkOM/qxSEw
hqlQS0OPiQqMJ8ck/AHDFP7IsDP1NqiS+zZgM8ysShTpKlz9hMeNvueAmMpZ2dJQzpbXTfklyJ/J
OVSOfv/oIyhIKCidw5qkqOQtBB0HizMmmLAuLnGQlwIu44Po4qmD+tAuS+Tvfg9fHMzG6HO+X8m1
033NpRLJ8wDmahKDintFSqfVExfKc6/oK0YzeJOuVlE9cwOFKPIAFXoC0gEbWZKMaR4cZ3Ad9RAF
o/Eo+ep5ceOg5GWxPKZr4bishBvUqdD32KrkUPrnz75MNODxIITFevn91v0KvqKQTiIU2TynMX5B
CAQJ4287oVrgSBoZdXBAwtpGUsR0t2zlr8GjLju5kJFfp3zK9bXtDb8ZH+v41lHLlQAVPHG5daDX
yAj5+JMYnlwBKlm0otGtz0YZCKo/fzry/mK35JhMTSowK3Pdk0hXp5Uq19+Lx5z0gfnDjYL/6CKD
5SaxQLkH4PmzdUOv3j7JIzXPRWHszt6Ahvnrv+lEsm/zW0qmNXmONqPucotmkRmRKZupMU2MVHuP
nniG7ifT1z6CcunC+IdicfXOK5SNoGIMkZtm0mX/uxlwuO+sSYktTqhj4WMID8FjOTNnvI0286ui
OuJN8P5Xs112aOxcqtPptR3LdiI+FCRH1kvlbTVtaTsGtJTRiBF59jQ9igjubl/yTv4IwfiLicAD
S1BjERr+EZUJ7Wrj9Z/HwPj5IxTZmDI1q8N0hbHBgqVRvVpaLoMs98qyD/+sKT1XHoNyd7D5F89E
R3lTX0CZFbPLntIyrS0vD5ED+QlRBYUUvFpI07EmFnuVvGUCNdoG9WFRl4o1UPgNzbV3OBNhVSSJ
/YtCuLy98VtYVl1w99GJek9I5rJaLj5We5jO+xife+hds22QXZEA+xnN5Y6Dgtwd23jvcsI2hQ1e
mD9tjTTiXSC/AdKQ3HlUD1fHPgAzTihwxBPYIJz3ZU0Zpy3yWrRoTd9NlobQ7j5rn0s0pGB46UB7
FC0pzFBXbM7I5qJnNxv6cMi5uFvPo6S+pB2hLcE+Azm8Qm8VBbvaZssrAfeXIYscauCBOAp8tPu2
QdNuSKNyIdmMdplMzDUfqlGwlTGnIA4T8sGa2Ww+KsKYj7sS5JTaAvBC97wkFT0s5ZzLnErkjTa6
KyU8D/tdsN7h0f+eBJQU4QtrRumX/rHizG614wRWqPD6VcRhStF3cPKYMx3ujwujz4sw65a0qwTs
yqZbY4f208lvAK/3DpGKR1U8lPH3BQCSDU5auOPWE8BhE1ZFb/Ijdc5jf0gPmlIzdJtFnN8qJhal
+f//+Hli5GBjST89uSE3PBWrNja7pRYT9Y2369CnFCfiP8hkJpAizwFLgA+lim7PP3fkyCStGptO
SBDJWm+gDURhjN4jlC1xPwW+BdPHDoI0siTobf5AB6r0wRKsdmv2xOVE4qflcXgYdTGp91FGcObm
DvLE7oowt61EHmWgER9ECIk5KHBhgBbVbRTTzIpQ0+shI+UvZJqHorCDB4byOoHF1fvF+4ksnX5e
fPTlmQCgkA6nfHOWaljsY99cmyessURPAcakzeI49Wh0z7FWWeeY9eq1uHgExl1ziqIZBkFXhwGJ
H0WEfaE+AgN/teK9zONPnfa+ibeRP38IZQcE98ep833J+qOe0lMJFhMg6/rcTUQUmzGv1fmJG0hu
tGEp/J9Gs0C2Mdaxn0OKbDMjeP85+MKsQyupPx2zdMdeai47SboEMI2Yy5gs87AOSTsOH9Gg8PLv
Im2tDuGT8aeUKdFQQWs4xy8NtAflDbW1ecoPYhOD9/PT8WgYXELVaqB0TkhONShllwYXpoLitkqq
gZbYX2xbrS5JnDzqXUJsprz7zA7cfBzOyEoQaLNUQF+6neEq0pfTgAs3OucIS9rpOSoGMwcu29Ce
rcdVRU6s4+YTDIGsVEQOQx7z6RP6N+n+8ImsxXgMr+F2tRNwVR0AV/f01okC1po+boVBO9u7OCub
7Q7rAWM0ms9cfVvHebmD5zQAgJGCP+WIuzkx8TxDhXtwz0APcGVy6L/UTBmrxgk9SuHY0Vlj1pwc
mq0uG5O1g4gvOyYlZOuz7AI1yKTAjyGZdo39ZqilGuZbmV+DgzwzJMUwr8ZZSqTWgnyMfavwOQbz
7ExK3rpTE2K/2C/983Ob7zns21ilW3GYgCXCeus0JgGb0FkKlJJE2ThFtyFlouYByUNoN7Qkl88q
ffOchtceoNPFp31M910E1qEBJw/IJfJIAUJRryZ0LQJuD0eT9cuK4MtacmLgBPBKsXtlibLxWyde
gN0p9MyR2YEMoYh/jdNlT3GF7lPivQsCLG9FjQVzIQ9aJKHnnJPamMrNfevEtro9MTFowWMTYtwZ
PPsigMkUUnT3QEuVkdW8aIf6qS1GehQlougnQ73/V3SMKsS75nPGcVDvOQxM4Yd6fw94Y1aElHJW
n+o0p5UwcCLOCGpCmqfM5eIC/iIVoijqLx+HixCJ37ysNi4tA2x5IZPhCmGQfmNzJ559H0zsG4GZ
aMNPdwkO1nkEbU7dDyBCX/X4CQ0cHnyxX89iM+7uaSRFd4bX9kcs3YUlVZ8W2sIRlfvhSmU2e8k6
FH4fUIPwsb46IGvaLLfXvD1M3wFulj7O60RvUSQqX5f2Y1GaL1s3k00ElFbbCVwwjpIOf8uR3w/u
xjxBHAmYpN0SwaHympoAl+KilrKIGrB7tmSse90C378Y5x8b76doKrDE5++yY2YZgTQbbzWq0Pim
UPlNG3U395GHOTToo76++++ezAbYtYHUpR8KBZ4/uFyfzv4reLMEYYNUD6HmakbwMS7LYLRkCNYP
qfdTNCEhiepmCiMlpt04mxjTzMIG7t1Mmg68S64N4pQ87fJnbZ0XdsmtfyGcfgPjg2eC3HKwMuEn
mZ1RzjHF8ZO99vNw2H6sDEYUL07rM2Susjzix3ZTzifKambqyPjXPDght4Faj8+VPss9a6a7MA9U
acnL0opX1lnK5dIVjkVT3FPMdGucjaPTdHyPErrdQc8pmFBcCUUi3PxYppnf/BbHMwR0nkawKgaF
mQS7fBLCqZ8qCUE8eGzQyE9QMHvUmRslIcg9zhgVulv/uaENGgpR7dJV2pwvqxH2vcOAvb1ZAkKD
CpTbJ6qCb9Ioa3xm3HE1AVy2fbgLaQ8YW8x5JtpDviW+wkpK3VhObEW9HwJq3YX6iAxVxbXxlHl7
BWyu+hOxM3uog7ClAYxgdcWb50uO++IN68766SyBNbv0H+KTy2AwoWRRi9ieYcpATYmEPFcF7rSk
bng5JA9w9/9oenUVtVtSaI9nZTxpoTQl68W6Y3+W5WzFRbErf7JZ7jE01y+T7V82oLLKY+GhcAB4
tgA0tj+L+b0KPARahTyKli517i+Xfv2NE0dJncrXaI4TrqtypXwl899JHktrFEr8XBtQl4zDboD/
sjyizO7Upa6lywnTuLLmhKr7ubJZaaLxkl4NC3+BS5Vtz0yWRtaJelPG63sMIbhkYCI0Qlwk8UKe
in4/n63/fKpgQSdb87SlAqhh/wmy5yIs7fte8ZaiDUjs4zm/mjdwC4js5BmkdIfm5NfDLuwjZlsx
4iDqenBc06uUz3m2tnXQo4/pjEA5s0sEqPAJSf87kJdvq5KbqfMSCoDo0ovN1/yx9dW70xuwaFLR
Ddn9iGZ9ZX0HSZjSHDXEJGyYsB2GTIl3y5GCLCRjBx5fGbeU9skGW2KIG1ffO5ysm/5dc3NdU/Of
nLZYGIcB+oCsSUsZH/t3N2geyXaytsSTUBl/fd7WYUg2bEWaRcIJTxGVpNth52/O3mtlOTcCX1yp
wf1DRmvKy3as4/CBxfpNlf3uChNa022DE9F3x7ox8FUDo9EAUvCtc46wVmcHsKxrzcpZsYqNJo7y
Xkc4tsv614Q9wLwF5NSo7XltQfNK81vXeuwHvE/IEDNnXOCMOLPYpD9uh3nGeIOXYxTr/Wbc62Wy
HOimtUqYjGw+iapRMlEFe1OLKfbhsTdJp0EARmhgGEqCocA+PEWvs/hf7uK/jKmLE/sF/Yw+VnqR
F59HdeHW0/DVHN2eLQ0bV+ubkUiIaJRotfotWeU3ItvHADpSdJefV8aqeOSURAs02+rGJ3qmteYg
aufUai8ppWm7hK58BLBOylveWDuIjMUjB82FMtohVOB4JyZquPcNgLHz1coYZqJTdjs+daT2RxmN
sXfGPEq6me3g85Q6IoJR2UrEExgQIYPxuG+C24fFwAZKETyl3PiLLzvKsQmQ0df0m9AIB0mmLaBB
m49ThTZCNVRBVj3EQKMNWP7S8CPDLkTjaZQM7cdi6A/Tdd+TDdzd2+zjnVK2b3k4nQJQ8DIydj2x
RcLlvGTsbN9/H7iGQ0XjnfRdRKQoYEM8ZcGvOeTDN3eguwUOTWvNe2J/MJlytO7wP7q4hm9D/+Jf
C6VEwYvTy6hOaH1Rl0tKKWr6jLHonodrQdzfXd50FLcMAWOPT8Nhfkx64yaZrirngPD6baPKv3Sg
gQeEeiSj7C+qb4tYg4jIv15LrSCbHhMbqVZ9BkWuu7aRBgQqy0YMBrNDiAfU6Ew7oxy3t1hyvLMV
IPhfcYSNEeW8bmbxIwDSYhbJCBpNZGAznZBUR9qUCqJdTIjkVQM5NWDEvEr4hyg7P9KRv7/nAe9r
Lm3t0ezZ2whP6bSc7scFF/uYUpMvAhapHCcFp5Twg3huq4fAD2GdY+WOgGegs1fe2DgIjnGbRBYK
PZ4qw/bhP4BQD+1Lpfbhovr1+AHbj8Sin7LERzrZbwkXl6/iOuxEiGOzMcdaWM+DhVuP4iMOg0/y
nrZf763ibV1241kcdTDRPNnrWfPjk7ZQPN80GuyNMsyQ1ENoby/pd14ifxtlpgx1POpbdt44X/ZW
TufyVXs3EYi5FtcLADS/xy2007Ovt7SIu00jOnKbCtH7/DSWBSNTOohKKM7AG0ExOUF5B5FCoKZq
jVFXmSoJmorvuMHvuJuzmzxlonSMtCtWJ33jHNtxLgeHDbUspURoUFfa8qdw0sWnNrNd/b2NmwaE
QAS0F8TkDk8IazyeqeJm3eiPj/3HKIYG2/ptwFhmc6ZrcQshRx+7n+pqxq0h4CBizdj4XkhAr+GT
rXGaYiQqFhF0sbAlvRt7v/7wVw5RVAu/JGfGxOZRb6ONDlfuGeafO/pCNHsjCFbhQnm5uFMJN4z9
fRWM6Losfzc12/bhUeqUvN+cKAqhdEJ7/RsFJKzL/1IXquwg/rTzLTUPOCrJ6AcQtS8CniZEwZfJ
zN2F25V83ubOzAoSr5gvx62F/48H+9GNrIrFrvA1kunMa/8Z62l0e9fvfzLAkYk9eakSk38jqbQh
Kpdfj1KbDgvyQIADSK9spZ6bKIWx8NR8PMoNiDxH1q9Yd23uayl7isf7w/2BCCQQx2fO7HiDTjyd
xWGhx/SA6qBc9Xw9TLjw6CSSTXs2wgtAdCXKzEH3/rJqsk9kWbxwBMmVpWLGbZ6/GQBhwegMU0+O
EAJ0RVglp6ItA6sxZY8tQcUujc1dYzrd7oU4WGalJLSaw9pJ5sOjJaEDI649hMCYjvOaDu0iykIn
JHMiFYrh30Nlvrap3Zwb3ApwTVXO1YrQQdCUIoG9Kr6wwqgluWWy9Fr96X1Xrc4Uce6qOTTO+Ixe
lN173uZPk8ZnHhIa+FelrFOmz0c0wk1JnImHhCHjnpvIMv24Jf2x3Gb9SixwG4bHUL9GWNeTUxq8
I9AfWdet9ttlCYQvF11crFu8t8gJR758Bo3PeDvcafrYn6t1syOs461bYo7Mi7WKDKVD43376HBv
X1BS1jasmNNzlZq6fsLzOhQ08dKi/gLxzgTkAlqHUG74OHd0iDcsHLtH72V4EWnIQbm71ckh1kYf
3SJbtguwhL3SDmvjwo9ZE3vfaVLMdY0q4adDtQzvUIgekBCVzSYuQj4bgaqYSWEb98eSaOaTSo2R
trElKc/a7T57zfqT/HlhQTbaCa5ttqgiOOaHW0oXAREJW3rMwbHNUPJCp44ZsuZTL3D8imN52fDu
pz2iQyzFHi3LxXY8EZ6sQFCPGHE8+VFF0qjiOnYbl9/C488l9vw+FlRwQrIVyyF1t1y4WzswSzbx
31iCRKVaunUIEaa/lj/aCgGqBx1GpBWj+I0ueVUtSbpm7ZFsA1c1hqFltKgoKXaM5On5h/AaAVKN
OLOURSH8/Cy4oYBrbxxg4WAcXhLRLyHs0x4bdBYsiMU8XfdjBAQkwgmWy8ghEKAk+cw7p/UlLenO
FENQswFXfAlWZBk6pGmmnkvjI/GGqmW/D5fj/t4IE8wBrbioYVZ2jWNuMO0xtkYXFNcCnWcu4esF
NZVgPXp0eXg393Hg4B9HIJ5IpLOaCrsTxMFCoD7eI3xDHz5efkTkOf3HMb0P7WZHE0LrRvayCQzJ
bmDzwPSq+E+htmM3K73Qrw99qO8fJwMwYSZ8eUoQaf0zXCgxMesxzt4mkQWAqzKsMB+eE5vzpOgQ
3XZjXvNU1v5W99SX66qB/PRrKpW1pdtn2cXzquCiLAKZxyDWO647D/afqPMUFvmGovYRLcxzrcH+
LVh2NUSsshniXLc0uPXqFibwCG5iWk91a9gsr/aJdZo6JDGv9lEHK6oBn9I7jpgVjQCW0wm4d5/6
/jBqdn1L+uFp1W6KQFQoeBKAuC0C1kyX3DSt4qAQx2k0qY+Jgo9WMcXBdNqS5NqKOIL400GmbDPn
J2Yqrl21RmrWFf4mC7jHkcuBp2e+NC9cGv92HLrCiiqNb6jbneCP+Ii9Tj5OvhGUbGM6cpr/LVUK
NdW+vE0YqC8DHfOhBb7Z/gFiIbhTzzqw8a64DdtSYI8aUncyt0K7kBQ1+6t6eM6hjVyho6XJZwZH
NLuMjXZkdj+ihncjO5AC7H4PZUuN2fdOizppZTQ8KEXcvtPgKYMIeFCswvRhTZTzGag4BGbeG2uC
NAfHqLUbqcUmHx3hy9Q2+69W9LjcTY+GnOS4qL91zZD7et5iP+aPicsy9WW/h0g9NLGj5WimfAjm
oOU6w//e/N4lfYi+kYuD/r7bSuwOwPVLkUOWAx1I0svyalMAR/BkNdv4rj2kS2/p3z/6VU59Oq/0
caia5gAXWuviUGlLSgNAftotZKj13lkvZ0Pxl+NG4Aiy07hwzgyNF7txQq1KjlIS8/xkTL7kytUw
UzuHKS8zpSBc0raMpwwTsMXzuXqY6I2F0PgKe2+Mzqg1QADk2B5wrJ+cC8QwSVAC4i1KMBJp0lO9
T100HNlL+ago83AShApZEoY1IMnthoeBu9hJyupNk1WIVwhM+UARS6Wh5DaXZljRdY10I0VptCFm
Km8ZKpiZP89McuYonmxhrv34gBnHokv0+K1ZSgTvTYEHHer1HtOM+AUJup3Jl8B390XivhkshDBm
6069PaXilsJfTtRyvgMRJQDbQedBrdN1KmlO2xQaHfX+lVVbZsUQv2fNZTaxISsu/PxXt8qM3ojd
o9YnpoJkT5DDEBKu1DkQdHYNVh2DXQ3mTj3H6hIDZVu6lSzxSLjabCSH8jUFkfveF/9I2rQxc399
Y2D+oEj5yMnaa4FX9Zl1tlq213e0oFqP3O3T4dOryRHsSVfflE5o07VY9qiytOyKWaHWxxb1PAaU
GHzhjG/TK4BKWfTRncOdd4ogOiE2TDJP+lGTpzPyK5L6FPBQm0IsZLU4Ap+NHf3NdSDik3qrAQjF
jsWTLDstX54n2tV+DU9aCSwgiPYSgS+vpF9BvOBq02zc2KDlLr4WZ/6lG+Simmnsf+/fXhRARE7P
8GVOSNDIWqnnZbGl7A5MI3nCY5SK9/kDp22rr3WXdPMmJ4pBg1pWF8GithiOckswlAIzYhr9u/wJ
x77qzgACDvFD3FJlr49gsst1wYIeqfgg3P4Sjh3NKCPT0LVymVKNhuxh4PP+SMzlKNmHQZ4LOtIg
kskjJmYGqa8M20ry/s4RsQNNveKjO2hY5V1ARfNoqdcC9kNkfejZj3O0jBK+E7Bm0v+D5RCexxMU
LPAa/MgPLi2peGSnL2uG1yOX6qy2ooJLGxFb+w+7QSrj/U1MR/gdWfMzYLj38OVPqtuv/9VLGJpY
PWUXi6RP8LSa7h8SRmnLckyxSdoGj4S7Oy1S3ZKhvPzTKE/NbrugIj7WPootn4MVDDxJ7IOUVp8z
jimj5kzoRbAoTuFHpTUCl1ej+brKijrSNOs117QSTqUMP8XsP6ZnP4cAf30mkzB8zgD5Fx8+qMhW
5qs1amgB13KrUeYwb9d4xUF8ldIXYb7FGHPSArbmUg6OvVDUSB2fIuTsEc201Z5b0ZVqCGIdD0PG
6c6gjiPPuzfP7UIq926oXvZOh7nAwGTdWp/dVYmtKdBX5vOBHiaekUy/6AIGNI8OjqpshN/QurSM
Va1D/bDUaIHZJLYoEiknh0+QsV5rhDW8Hj6n6DgSGlfG6eXAgHhKWcT4E0K/Auz2ub+RwqbMeEOg
QrIYrAOxmKwX69MD7Byh91atshJDWE7qeqDXgUt3H67N0WKMI48nf6WDv1GEO2JRgJqiayEFTayO
qkisrm64O5FIIXtky2X6Vc0lWVB9OENNjUU/XYr/IEgMCDp2+S/+e2oaZKTGDBv0NjenL8NGTsfx
/7LbHT+NFCTiVmRPt39JzAm6w814k90RACylgkzE3XZtYqJH1lKPoRyClZkoHq4RtGmnXJAIpe5a
dLAua9BaRG2Ci7jkTmvg8yjRuseu85Pw9BqnD1p+gpU7BgL1CXkfOz1CerqpymKYZ++QvzRvyUM1
YcC0Rq0tBmuPu+ktrUOn0TreYzUvNBkMysUCLJrPjWcK/ehERBwBCEolATCLsUDEc1DyjS/Sbriu
E2UGoA+8zoGejCNM8SVjE5f6r3LZ2CT50Y3AftXSBwIaiVmDQRim199ltv3Qj1UELeXCz09V3I8Z
4SoOdowzD5goJZxu5XfXJt/6CK1XCHb4os7LYFtiCiH8di2v8KQg5wTi/P26oBTed3fkBhNlOZv7
QmuXL7cJSPsIqJLWz607KqEVQ0smvBfao69C2RB3UhyRttQTV6gAmxRTn3jlZeR08IaoV7z24RY9
d7LvYqyqYXWa296EO9nP5miHy7nTf2l3bXlXrWduITfwlSAC+0AgPTHyG1GvWHiR/r4exSTOoeOq
DT9bi6JyGGFlh9K3Qm7RCW5zindEW7GSf24LHvaUUhKr1X06yGDC3K085E4S3k9xMUyVQgOdS4A+
4rK9LEaG4cnx72ygQN862ijR76ceayi2QiasxD8CEjjxkG2ZAnyUjVgADbpwS8WEr2K+9ApdzprX
BfoSkAnOtgIYKW8wb2U81yM8RPh1eYniYcOKcbLnHMppO7B9TSNwuMuIBch3gTb5KtvJCn+H1EJ4
YCkrHG9d/V1BPnChEGFaRK7C5r13KIgzv0SaJ5ELZxWiGWohuK6LVR/NJyUYcRsoxa+OC+eO1KP/
mTA4HuOOYwCzh5At5LneZ5kqDP3Y+rMBKy0YB/YMZXnE+5M24gjROXUfqkxeLgEaPykkEBo+6jOd
mE9R5iruJQ5aqtLbwl+CtswMgZx5MHIzAZaOdeX5F7gPMAl4/P3x+M6c2TJgifiFXQ7us0cCc81j
nq6JverDKeGQffUbLgJhqKrN08OrsEDND2empBX4A8oGgWmvtabC/xf64N3j1l94QQ4oL+LEosD+
gUCI7dXaARfmJiVfPRjp/C+4YNCL5n9ywXbX0y6iX4M+LUvUpcOrFfztItllNGWWsJ/JfFJKyUm/
rojwJ2K9CDWCCdoet+Oc/qlY0djowGVV8y1sEJ1sGyk17de4IZYrNdznc53R9Fb15hQXi2DiuamZ
MbIwsOdRp5mRf5yr3AACa3VsaogmEKDnVvti+o0TBtm8is7WiOKIeWHSS4x/LWzPIJsRkfQMzTGE
H8/wrk/PM3R7H55gqUKaomZQHrwGAQfv71DwHj4uC3XjkKbvatTyXtMmcqwAxvV58/R0RlVnmU3a
KlFDd3BGWelulQCRMa3NWkxgymownjcR0VVMuvvmNnMGFEQ+WzqVAxPKXPjz42K/nLqiC5KXDjCH
6JOJCX34Aj+ZCYz78EWSvk1vQWlq+gHhw9S9jQjQwMoqxBAFluLt4HfEkIObOv7omE8WYjThxW6O
AxoRCf4zv5+hwWudmj94smqojnRqStsMLTbqSmjIQhU63rkl68rgl3F5EsrUuPUkQ8TsDL3n8XBM
89JvTxgElaIstbcKiVMJL1bthzLF+GY27fzjrEHjXyHcZbNm9r625UCbUxErERJEPKnQX2leF0l5
04FUznDraGNPmM2HowUNWE59QgccVEU1EucY6oWdm7jPgA4qQUnZAGGtadDMgyIjsScQ+Mb2ITvy
XVrGpGTsPNy5XdDXCvNW1p+0Uw+uPyXt38YiZYVmrecSfFyhbhctGXpYAi1SJIIqmS7oGk0x5eQa
frX68d1ghJVI4F4lJb1FBszuSWS2dMmgjPChfbPYOJ+mgKNHVeTxRQ/2d05kNRKtId0TXDvhi0qD
FCFwYZSJt/4r1TKivPiSe8768lhynHXfVjtOlYvdF/rqPiuY6c1dldZpZCSKsMS1jEgLpO7UTEtQ
S5P3wBBfx4F0ZPXAuiESNkmGNWME8TUGWpnrkyqCi9xYCT85uBOM8KBWgNeeFlVnCgH9zRLb2eeJ
y5ccBUl6XDsHxMrP4fG09Rs1nNOgDJgDVidnngFixxAOg2fvX0orTNz6wXdYzpm7ISHL5koeR1j3
59wypSJcYzFnTY35Y3Ys60eGNarSQF/CuiVpMwyyvgdxOLRCjoSv69UWbL+wr17VtgV6x2g3q5gT
7qKVhv5fuqkLla6N2sOPnERVLW0Slgx7VPVhfSgcuheWGkFel6XNvsctRydlaS9WcWl801SQJzMb
F6gtvqoXFZthMNUf4TbruX9vZbYWCcHSTMGGr25SnzBzTMFIvvrkQGm5Fwnuey0MWOFaBpxN6EG8
Rdp556ZIy2JDJ07k+xMPKSQImWSyL/xZRpvkj+CfHp/8sVOJM+6UeXzhUI+VVMCwPffCqATdcVR7
xV+oRG5v6sEw/GtvoyNvEQzig4avl0IpQumHVCZkK8H91o2oOmfvZtW0uKKWonLkqJNSgauAmXa/
PB9P8qNkKtClcdmUKysAb6+hk3xrkUdhjEGjCHs9nmR+wLfxKTYCXmjNNHY14Mizqa8aTFFOND2v
RB+KuNXmJmlFXZkGMVlH7CHE4sWmlH1AcTeKLQGqcIMszU2mukF+Ye5EESEM4kTdcGsnHMTCo7Z3
NxQClxZ9ae53MTN3FbebRbAfGgWq7OBJlEiy2zPFAQhdTI/ptWEVHGmcpyBXt2m73IwXOBg8FU4V
lNumfEIKx/CnsvGmy4/BElhi+GmwTCKTdKgGmZLJeYqC7yd3tZBeGPTJ4hEPoOZhUEgOZJrrPr9R
KUZ/rffFrNYHtQK05x1IxUpQv+ZCe7En/ZMsMh5/DZlogts/Anya4MEMu3F+NXtpzHHUF5h/F6Pe
sqVj7G17SHXiaEfW59F5EH3yJalPy73Ks1HJYCOA3/fH0CMu+aH7cxOfdyXmpwwYyG8ibQikPBXM
OWu+UslKwqnNUwe6kPEJM2AALOp2RNMHk/RGufKkyG50qsfxNOwl7ooMuTVVd+QE+HM9+yMTo+uO
tgmno2I6wGT/fx9shJkNsMK3+dHq4PM9bQyk/vIQt6lAEHg6HFyyOkqUG2SQbQsmy67nMRl4IIlA
LU4P9VQ5zxRJL2YyuL7lEh31iHldG4H/7AGp/RGqF1bW0+2VGXXLWe9nzWjZ7+PTbYsQbmyJU7lr
om9wzyEyBU0+fPjzxye3w3Z3MbjG9XFPrTlolmfEChoAAiR6YR3XpzvC37NJvQWTD0kurw7P/Njk
fXQ1TdJtTb4Z72WoHuCWcOXpBXCl+bgNxbbwTXOiKr9pGNOl0mAEbIWE+CACaImJn4Itm2H/95zw
N/ND3iJg/doYcSn04F7VF77oixO79WdDoFD5OjWHAUa+ISrppOGqaooyLOvV0tCRTzbMvl0D2h65
HFzVkivfz8hlAA8C2UpEVlAkjEbxXNe+mwixRoM6uLXAAl0WNt3hib0oFlBr4fyyz+6nvilNzNgY
FFyICFQfqBQ+Hds5Dpx4DMC84p4FL+ss0tQsQPZOrFL1E1HYPPrttcwT7+HET7gA9QEYCYa9OB8b
KsI+0lPl56YjnOAUYUNDk+YAtWWOP5HlJgjDTHUBFb0HULgJHsw1WXBF1jTDMZAz5W88CAK2nNJo
NHFRdTszktxcKRLlNc0yakI7jKod5uFufnp2OVm8YqD36tW56b+G/nCEgQAILLyikPOTz1NBrRoQ
ac1NRNKPsandzQpFrVwY2ZU/iwHOtzWe+2CsweidKpu0mBnqBKEJhdeG26Tzb2mF0e61L6zrQ/2O
nQuPn66FiAvB4OYv7mC5AcgMlkXmlBiHI80Fos2GHKqiBM6Ar4yjn/kiBV7wieW9ULlJuCAV/pDK
Ls6ugHcVg7ITNSTOTKPJYKOibIjRu+lNhCe7cLxfH68UxlPI5r0tmHhdxuxOHQE7uNxa7GzOsdYk
3rBG3Z3R0l+e63NCFCHl7SQlhGA1VI46hNTvttiwxFdnRQdlWwr0f0MAr7iPqh2vzu0lrzrzyTZW
n6gdkUKGLm20ycGaS1mofAea0ykE/02zeqXWf2yiGBWti4j/a1IoRMbzUCoYpqx161tUjeHTkvxG
BJK6rTg6/dDN0a30yWqLbAaVAMbq2aKyuVqqLYlpTe37s3FJY5or2rB1/RgaKxezdrR1MqaqsqMj
KG6QY4BC8LWvWn5s717wBXDGxTPhFHIks8xnN00/9YyOSKHAhKCZpv/PWiMqljjIvxs4auhnpY7f
isjmpq4bVujbkfecgtdpcsOCrsxSHL0cuxpkf8IaT2kHyEMsF19rXOzXQNBOD0ci/9iH+ID1odBc
27PzyjEV/mWrvGbdBE7pBp8d28znH4qJmxITkgL+SnHyLVqkiXy9IlnpuhluNecImsr6l547xdjg
7t1aWMb7zHB7UONi6/SzdHq/u5Esjw0cXpa+LmokLUMxzfHPbcIIQ4ibSbb18SeUlH2m0DfX8hbf
O56jBYz2tVGPr/7TWVoBaGR5g+HEsCid26LZfiP4jD9ua8tvXewNnwCmp9xupQk9j6NH2nztpmNG
jtwwi9OGSWYoRtaUx8ovgb6YFs1jEH21AQgnAB5ynJZKH7wE4Fse8UAH0j8z28Eu+Fyy6p2Oqpag
/esK9Bbmdf6BwNauswpfbpBp9X0Lc8lCH2j56LlBMy3X6+KbVmJjAjmF7CttTooX2AkridRWspH4
Ruvhl3UOWU3cwuX/DsqTaqQB4Nvbuy6DX/Jv0A7d2IFznx53QTcdwWT4d+TWcnL5njtudTMrp7CQ
Izubmzh3tE9a6e7d3VWP3oB3woU3wgcps+J4qkLIuerQMHnc8YSHF3JVe2ZgwvX8EbuvOLmZxZMN
002YDMjRM06OdVZcyktl8uFQU94y6p4+D80CRorCbwE4D96XlAcLSVsuDkPSper49ErLfgB6fkAh
3bYLsKs3fJxSD+BBrxJHihGF04SU+b7A3dyXuqt1b2p8vmfmm5Zyngv1hHmG4WEFITp+A9L4Gy4L
p2gEB3I5xjz4HncwFiEqp9GGgC6ILH6oka8iVqdYnu3c5XBoNo8jN4zCS0nslQc8UwKfT9SILycj
3l3XJZ8k6MhAubVJv9dWkv343E5MCwpzun7oBHAMVzUys7oZTbKpfXdiIvgAyO2ixR1w4Ah30WWS
/pZbzpB3+vDsNFdoOGmOiHj9Kcr7kSAkcW0YaX1VEE0tQ16fKox1vUMTmPL9oI8BQnJQh9360SJK
XyL6PQMJO5v9w97JQ773b367V5WF4TDtDhXmuy0l3+1TGlyBdKHViVV3X5U/BX6Cr/bzFSzzKrM5
HOoOFq/WbBMCmCl0/BFjNSNw68ZcEt6enDbsvgttIfUQRoJfiQ6WPXQhAX9L2Hh6x589xS1dznmG
yfsW3m0Mw12ZquNIKcadXoJYdhmDyF7UO4v1BiS/yiBF7aqlHUs3Se1d8cySiF3cVQhpuQx+mRNa
EzfXl0KeDBTKbtRnyrYXRmR3RJ+a8krkgqxNI81C45uMaxcvdzPZ3LKQvPwMLZhphX7Bih6xVoh0
1JmfznkL/3Vo/LvQBfw99uI9ZhSG7KPKDyMfMKNz8YKksEE0FPsKLkiyIY3pOD4DbLpiTqGvJ8eK
cYDO5m9lAF9FmfZLumVCYqLzaIYF4ml8HsjCCkEX0fDfFS/d2QCutA9O96Wjfjufo+lWW2I87nCP
qG8svdqUI9epI5c7M1FEx4BY9Gf2y6dDYH5hcM15pZXejYk3xUIN38TxhtDhoELB8rBA05QaX+R3
SzlWF931q0marLfI9DUICRxpUwxMw3PAGlaerqxxUZQg/NmmtC9raocdzjszn6qcxCqaXKjzeG6B
mBKOm4H6rPCF8LCyjnp1oLbhaOuBhz+6aXjDKczAT5YmceqZ85CoFbIdSX3pTuKR8ztESc+r/uDj
wDrFLVsuOzDNUo7tXKWZDk3hB042E4NuYIsiblSRfFCulILdDvRqOrMy398ayTfA59Q4rzMQ3h8f
611xrV3sHinMRMEg7EzdXmabqJkJ6kLoJiiDQnpBMJqqELsMvKS+GCfQapgyxOnqdnYqtOQuu28n
ruLWGL4/LrDI4pwpu56bqQdfFQNffhntJWi3nZQTFLayA4J6KsHrz9BxCGR0uLr9HAMfrQt/YO9h
3/4PZgUMmqWMiqrBoJhZO7cJFIDYaouZr2CqdZqZ1112/u5Tor7U/GJgHGKH7xAeDpaQzNQYeWac
SO55LLBrvUGxpCBAS9bJFZaDfgWmR96sUMD2JkU+uYW03KTZOD/63CMZTWd4NX/hKM8wgV7IE4iG
55dsJpiuWTdmvsaIHAY2ax/rtoSQicQPkmmAdY1euXxbTL/vN9uHITDY/buO/WEu9GkY6lu/lIIu
oQ5T1Ctjb/15Usx7V/4ds9Q8fJmonT9/a3gFjwgW6mhsQlxx+O+oH9yAmmcYhGrXVecRY/D/7wjs
eE4YJcXli3TQHMqyMjE1uhuh3rpUI5HeecIza0VofOncsFJEHFg3Ve+YxXaubbNYCdUiNsF3TTP9
nZaUEDN5rQFFRGvboTRsLk15HtMOV040DQczC7/Rhiclk9nItAk66zMOYUgNAy4wdXO3qzZLyAOJ
CoXrVRXrkn51YI3Ad6q31wLb4zm4B0RkKDJaPpyKhfDProCfKMgut6GPTbnRhsqu/JQelgSV829I
dqeWEOxegAXPBkJsKBZQATEknN0R4NQh7TvStYA8zVOzbSu/awQYmVMy1gM/w17aLLcStPQIHzg8
wZAiQgmAPmBV726yd469QBoWHybAwvkJBkIhXwYWcAB6IIHe/e6Yx0uH9swkr8IsVTKCqL4MvbUd
Mv+PifM1P2zNwkejUsbEOe2jsYJ3Y32z0MFHWL1/hJ2sjcQAWeVqtVQpYuaYRXpZVuaDQRnxIZYI
HQJAesyoD38q1OY8b2tzXtxDhfI/5YEblzdlCUkbYwv+gnfr3YJQzazJYI13H3e4hjI7IZuera8c
N1j3t5JOlhvwraYacdHKvU9nm90xT+8X+hX/paovqV2+z9S3f4HxMJGQLQ5hLnixshkrWFtjlhlX
IzfgANJmlXLhkddJRR6MWpDmikbIHLwCnmW3mRBco53V8BT3Il+Dk8ATXWOCFFDybc/RqDHxR/ss
WvEAG7TCs9SphcJWp9JiXMtxQXgq++IDHSxeaRbTu3n86/QathruZht7a7jOB9oDQUyI5Frt7ZJZ
aovx05zwKiA6qbFfwV61MqevnNH8t8KC62OSjbRvH4O90RKbh3UQw73JsdqeZWIGfKWrHw5nP5+7
eJAcxsIsSd9PqpfAB4AVGk7kwQIaWsMYlv1Nc3TQTbXFG0DZZtwrN5+b2JlMuqpkqjK3cHvZ8zBP
63R8vowNSPCWERuYuxjD4t67HJZZS0a1OPqBMry/R+xxDvTQ1azPnhPcyZ91xIhsQkjmQnuE4CLE
jPmkSCzlXBX7aBlY+I/PdXDWM2y1ep1ftCJqdjw5i1CT84BrmE8RRRA2AcFnKSAMTkd7til0L707
GGo9jftB/0NPagXq7IAbQ88SUhjOy3lZuzE4n7NZurrF4nf/6fJk5hexGc3kRZ4umbSGB2wKCf6Z
K6GOYOh5DFcf7QczogH2Kse+wd07wW/vefXx9rJMwHZqVxQNnjer3awQoDV1eNMRVTy6GyRpic/G
Yc85QNWIG0KQVp/LNwSJ+jZxo+WMSY2MgoTAvsj78wjqivn3wVmUVn7K8fxFfBFYWu3BXbzkVQ0s
ymK402C8Z1th+qdcIWvgsrUNziycTbXuaRg5cRhKVkpR4uIhUyavwSbnLjQQlHnH2IAquFOAl9n/
dtvGiHM5kutndZ9yTBpn1+2wHopGAOVKHZlJhsEwgv+uH2feCgFKnSSQe3BIo2gqyGq1DPPNr53h
3s/kPopJo+92tjicuKxgk8FnvSxbSryWXPmkK86mHX+nzvd/f7VvvNmMuaYw3wW+YxOrTtJ4RWxb
oiSqq8xGE6J3/JhWg8joamWYCi/MRYJVY3JSCm2KaNEwqdloHomQ5rxYZDSt636yoiUMkiN6Fgne
c5LiCEUpBwKDErq7OG+8ZbF6suWGgS13uT2eVcEAUV5K0lzVcLxlGTob1Bck94wdEoKAAc44InGE
ghxKyV9CDWCr0/ZKXR74WKX6oppo9QoJ5YROA9u7KiFmmVTa24GDw6Fe9JEOyVX4SYnpGPNAlGdT
1pAPsXBYTX6kN0nEfeFcfWeb5aU9yS7R7O8D9sWbmLPo7tXuHKVx2UHJ6q9N0Pey7WHnOAkrh+Bl
+b0pSnPo49d0yj8Y5C9jyfjkWm/zjJJpJMhWyfU3DiOwuawjrM9I6rjnncpziuShqJtmlessF9FX
KXWuY9wontGKFoRTkcbfM/qHadqOCfWYlvooSD5hEvuaHttB2sIYTuLic5BykqTdkEZHaDfnzQ+N
Ofm/pnPlQZBGuvjC2l6/IKyYK+UMRQ+1+NjQvRIb9TC8fCs8f3pO/d8mL8YvDf/GA4xONc9C33jx
U91r8iPZhw/zwoHZrEl6TWqm4NRCD7tT8t7CzRSftx2xekXo++ygxFVUAV8xqM8MMQ6CReXDpU6q
elQNEF/op31gburG710z+McOVgmq94GzzL4o3k82Y/YaWUYAPJ+SAt+VMl5sPqMed/IrG6sh9U0Q
dvtHn4sBg+FSlv8eEb9MLn2D/mK9UJpcW9EWZH6+EUb/anujToEulf4J3BlUTfK+aUaeaGez2rJL
a/lHK/ddtRLzIjFKhV/QmcZ0gQtrVtByLq/OiLcfBka5fCSHJvH+TVjfsAtYMk7Qu9wvzI/6zrYQ
WfL2FhyHhS8O9pjuGdOLNvvMbaKAEb7ZtSnjzwqPrbb637J3JvWD9+tiBHmQEAfw6cr7U2DkncCJ
KvcS+C8DdLoLlSe9TS7l5nC6TEt2mr8azMNxSEtP2vS6doVa0D1zRp4IdvuOL8yfOf+R6dAcZNAV
EFTdISYilAhKS8LneKSlqwH8KpiPbjB/NsBhbd7Kp3OgEAvCI3zYncdDDaG+ihbzSQXXGLkPG2B/
aVgYIZHRRjUG2Wno4qL+SQWNKNWQaiRFbfoLkaBirElRLh4+ml6qnN9LInppBvgSrCCDrboq41CQ
PsyF+SRBAFaQHY2NKxMe8dHnM4hK77Z+gUd/kbdSTT/y/Rm26rXmg2HHIEDSjcbIGY3Y5dkbNzOM
PZeaz4LN4rii8PuaQfpgZDgoxDrl8MnvX0feAE0fcWi/q4aYVfP2vevoFe3p4vdOntZc1sJF5UMF
gfCXeCyvgmH8exPPnbWhTPiQLTsFNvSYmAWnYVKjpBDv5z0pWxTdLP5iRIbJljdTnquVaX8EZ3Zk
/CY5VRdgzuwxDJD4WLk4bPtozHr8PPQlipDK7fxdDKmz0iI1LVc9C/lf7EDw0LMXKgzOSrBBUbf4
nbGew3zosOXYU8qGNexWjbYvyQZzF1UqcnuDSCttogkdpupA4vnoZet/OctLgSKIEvS+O9ZTb70R
ziiJ/g3eRtiHpT63Pp0TmHqax7RMR83PJ+8k4oxYP4coC6BJIgt3ZHnDICj5iJ7Rd5TNFxMhlvbW
2MAB2uYutDPeyK2iV/aUUweNxuatwhFZnSD0ToWYzuBCAEMy6ua71iTqgxSUya84aAvDnZuk1QAZ
+hwqJ28jeeZG9+92emlC9fkN8/IIBPe8Ti7A58vn2KuAZEe6rRwNGc5pWveW59m6CorqB0fyJexa
sni8dwh3hH7gfm7/TuBKurcN2wgzgLO9ThrBArk46Uqr60z7ISU2pMrIoKAcJlo9IyjsbzAOjOfk
UzQKAOq4elMBjuPBnPNvcpPrw5f9tDLXLmSJ7d0zcAYjNo3Enniip16Q8yZa9ojRGsra77VbMkt7
DVoFxdJztLMXp3MPdwVcW0U5TtU/Tbxz3Kw2vkaM62YziEmjgBqjhBpsrrTB5nghpVeTH7mr8d6A
C4IFEK+ybZctSjkhbKVKd0fFMBGJIx/nRMXwKB1gMLeVoR6mn0HPYi8xERxt7VuSHYoj2vARQP+M
ZrmZhO7y5lSviV36d9aTfwJt75haPWfrTan+NOAct+anOQtnLswh5oy++YEfgZN8bl4tGKkx91T4
XzDPqk2DJcJoZtbC8o4iBx27N9GqFZM0Oq479uvOkJJ3Bz9MsdnaxQ7wbZWTCS2YRKFe1UvMSyVF
be0bb+6Rd+8vz2E7WT1ejhWpS0ZUAhxtdfGTXdOjg7Ki+bvz2TSAk8sD8L7kQXwrTLLfaPD7jCUN
gdqVxzN7hqw46Yy8Rme4Up9CUNEL3na3mExTllpvnSwS6RWyNP5QxFDCUiQmX5ku8qQnImT1htfd
SjovjYeV0avZVQj3L/UMk6MM8kR205WQydjogYt1zb8zCg6UJ9hoILHrYywyp91op/b5adGYk395
wJkzPYeZtOGNJrN9XAhjmyW4GC5ofy2exvtxWLhrwkLPsseyFwLHxN0OPiiWzBVDMZ+QiOvNfii/
uC0tLUd9R214v3myEAV2p1i7cWnYFNwPI2evaEvUl/WDQQkQcrNkJkbYm2NyAXe3Madne8Bx5il2
mukUcK4qnR9Ic+TpZ+VlkCGTR9QhgJFcZVJR2FGu3cZoXoOLBuH8lBfEONmufzn9+kdEtWhwQ+6/
MY64kJkP2cHCAblu2prMtBy10qLsOpxR4Mx0WBhNnSYPKd/nNPqT7Dnf5hbgbkG1MDv7hgQjd0Qw
w3inr8DZmUzDPoPKpwtsqtrrGRJ87yL0D+Shq+zGeJ9djZ1Xvqk7rz+OBUf05BPHRlZO6FeCREjY
CXcBER54h5CODJnYXlz674f9H/j/BKhwS7qXcP9mCnuC9mRrDtMHrFDv0cQLKLkh513b0netUk/H
ql2HZpa//3PpDzdfLMJKACYPZKNACiqdE7FjJ69DpG7YWwfsx0aaiifWZvCvCAapiT/S0OI6X6Ph
v/mL3pYkn0gQLtHppP8Jw/x5ps7VgnADShkkxPDxOxv9v58zkCFI6XQymurE+XhqtztQHkRbMQJG
H2gxHRtz60Aw6FX+78Y1i5lfdQswxTe/OKCKXPyirPKOXzfdzHRUJ5Jr8pFaUpZh28SbM8VaMw2t
TYJ1zXb81jJ08mswps3NQCDvbGIDcw3xFq4FueA8rvuPYf+GqUGf37bYC5P+LPMT5TdpR3SkK8ko
ZOUxz7FkSZeHvUuzKC0GH+W+3zaCGVq1eKe0o8iAIkPl1UIGH2/5lcQ+3Qhswdtns+r2aIkIRJXH
FRLMdQ9iJHA4txJveeUu608G4b+/mllI/92jnSGHxVyYHGZ7V9SnQUO/QMK8yMPE/jlcxqvInpyt
CxoYyVLaPK01lwqbZKWmC0AaTTORFZ+HsVJqLVP7J3Od98vDZx5clnhdApPRsh+Y9CLoe+0LZwir
ZqWuve16yIiwOyxgFzArgO+yJRRX7HFRAfyNtGGYlqQJrEqlZgYUIkJu36KqgP6aVT6QpFhptbls
A6wa6bDTlivegwtOHEjuTN/PvFdL1fbeqTywf820MYstEWRziYZWHA3sJNL6GNJs1rV+tyrEUOdz
7Fi4j9FkqyMJ8OL/5tmaR8v5NoHb0njZL7bILenUZPs2m0NvzVuoNu67hz/Cuy8v9Byc41VUr1Hj
nQApmlCVFPQF4+cxO+Dh3aduWKyKc71nTJQWX4K0EPfmZgmFcYiVrfi5AUOfvdRC08/FlQm6Czmb
bilgg8cUmG6zlN5pN6L8LUsjXYArAk2ZX+xSAogQmvZ8IemlxGbrlYxuORW6kjaL/1+/+xHae+5+
YDvw+AzFZt4P7KgPxtN6imquUVWMQ8ej3v8gYjBA+fX6f/6uCpmWV9JHwV7rHy84OBDqIHYxFon0
9oQTCBS1DjDyvfqjsFOyG3AA/Lt0JrF3xHkFncOrdIn7ne4qIAvSbfn1LDgkclatgALn0IP9/cVS
0VNdDj2DQUTp+hmxZNwcGWxMKz9J05NDU/GB9RrTecabiOruQAx3jLiQAuqKuZLIAdpp7K4grzL8
IeTRw8UV14+tfzzwdUi1kGxMQc2bc2Ri9ICE/oQsg3sUpqkZnX0bdu9X5GBCz7R/aKuxIoUAAqw0
//AZiOkjRHAHnjhmzVw/B6ezw+6fSE4SDPN8zlUyVZSSdbKyg/SWvfF1ZogAj7c7xxw/M7qmbwzL
jtBb0Jmacj/yoMS7Rh4uXHrPrUW9AUDEEsgiIdEVFEt8zq3F87n9xRNe8sZEHyrRSH3dD8NhSSvj
7ldqVF2yD8/sfEKdIZeNqsiVTgv6PbZXLYy1P7NZz9+hd8Qu8+YknOnVTCS34dPkWO0QYuHOKMQb
zgNsHvfiu/lIeJHQR2BZR6bDP1OcSU3AWKObBhmIwt1vylx5cdwjusqxOK9+YE61E9ig0MmPpNCh
SMrJfua01WHN8xuMMZyzD+3lYDGasdRbqzKuy01ANX0gscS7ug1z1Zg+1ieB87pv0Dyn0HM6KvIU
Z9dPExw5RxgL1UulYVnxSgrBHPle5qjtogJmDZ/I5hDSvBFDX14mLfhRXF+WOv9C9OkrIyrcqEmM
QJz5lgyuWxQ0L+qyNLRzwjOXPpxM73BSitr5y6+NPaqDebA3fpk/INpAc5vT+OmzWhxLFUzwi9A3
acvLfMPn6HKcLaFJoJWUod07Dngl50vOYGquIG2BAtsX5S2NWkspUvwzm9juYiK00VSRs08OhBoN
mHmgV/toGdXzs/09qmfxEZnIPWPoMJk80tAxJBXc+sgXnebvFbBu6vnsfIQloOFmIYGWbKTb7qTI
7w1ve/fadFWz58N941xZ79jos/hO146IahYXF9U8Fkw+4U0WA0OS9y8xieXdxWuX2uctN5bN5TbS
yFM8wVqaz91wj95AZch3OfoIpiNnGwoBx0Ovf4hvaxDTouQ8BuUGsl/02n9tYu9QYzH+f0CA+sfF
JhtZkXgzLb1c1rWAUiVIVAAgfAU+PutnjWcsGTHFoy4ngSK0d8e63V3Vx3epsr93m1ekaijBypf9
/95GGosDLgVqMbIQJ1BWMlBIYJbVLgGJXInHnfY1ZmpxMb2pB8WaASQJcSHTdDJ8a5nm5JGmzrFm
vSIQYoLOEDLEWsjFBdgeqa9L1iZ1tG98lb+Oh7k4aSx/2fMSIIt1Acx7BWh7wT7ipmMIjSPorNOk
J60UXaIs4wBn70D0DzgIYt/1AwqTBz6jQO65ffZg15zIdu7mUJe7gpjAnhmtg333/XBK0BDpR+cC
Wb1Fp6cMNoNuXPdLmqAmIxFhpVFsA079zCM1BhQ7wtoT/DySRCoC7RDi8dh13BaAYsnfnCEA6RXR
NvcahcmWwHGKmx1n/ETODvDFi2uLiBbgfrrWT1F4DkmLxDt/ZGxb12IfEz82pHNz1PGAl8HisAxz
GlGyg2YfUnI/JSBy1J1MljuAOyMhLdrAY4uX3xJiPFUr+9rE02LIVjYl3Qk416/UFAlaPGI4XVAZ
YrOXHhiU6Q60/geh8bxV85wfdDKge9JPH6MhCxQwGPH5JUmgNtPtvkM2XoyxCvnVXE3TrvXxOwAE
C7/wGIAdIf/grYzAJZFgo5MEfauK3lJecoBwzelOnlfNAHarIJUHXF5L+I0EyvXHtgLgfm7J36Ma
7quVY1e81M/18p+KO39t323T5PW6Scoi9bFj9oDqauCjZuow8iqMAfDHIWRcWr24xzt6om0eRBAI
f76ltm/9P4b7vKaI87q6gH8H5GSwdzHw4VqSXfehHZiTQ49FkT8S8A0SPgWjvWLhAeK0JuY32Wr5
0okrJQraOCjG5FtO2IV+8xaRbYXMS8laU2m4WfETY8tje7HEVtF7HY6fnNjb5nzSqupuI+Mty/17
6uQHHOsCgFVCTUZ5GB+HJP6kNuXPX9U29VPUWWw8eGSq68pQ1UMulw25t+qAUYHiknxVXsFlHFbT
4APpiviwPewdLB5wASkYOlnbvkTAKCb2MOrMrkQOuuG8jltdLcmI3tLX+axsn86YJgI3XCs19LmE
gpgixtOiPaS7wamF+7r7WJxE3k6qf/hghFSearIMNU8OdezPhdP0tRQsBc64Jx/c+Ya6CUYffKvw
PUamMgEpQOk60nQ9wZRrvtTGDasUdCxCcdxtjlj9T6Kkk1+EWw1ma8Rag1RVTkn0Hn+mgK1hawYA
6xDNoBKaYjR+YoIsVF9dtc9g/ACZlpcZcJiIZLTgcQV97iuW4y4mk3ZQW3/31RbJaBfKZkyG7K1F
uEdFa4rOkDMRpxiPz+Mmtt9pLa41ZUFxbuYc1GsMfpsWikcMaGfokseVZEgPFIYUE2rgVU1ZqjPr
1v3QPOv7t5D+CAd0iPTuRPLgHNludwtABuufJ+hZBcErqT28M2YCjRvcB4gLAl21TzxNVaBfsB8B
eNxX2a89E0YjnJkogC/u1J6g+jxq2gvUHS0xz6xj2mVu5Tks+hWqfCR7HRVA0flBF3jIauud8S8t
RmzUAmjzV/2qGufCpjoLCyaawpQa3hp5beZ+DlH8ojNBzKLx4bOA96WNbeA4OiBhGJ/rZ0lGfoBL
7WR3Y3O5fzIyYjjuPtol7lxCB2GtX5yxuwvodgCaSJbli7ca+s8M0+gQkQNU+lJaXlzRYSUzl0hk
wbRhkDsf6I45gYX7jArJUwT/ymzvTsQGLm9siv9tyDBcyge2kZVpzJ2Jlnpkbux/O8v8HkhcIdPO
BNZ0rnZnTqpE8HzKljaN5QOC76J77iDfeVohW0RMz24/Ea4DJ+jNGGcra2L4FIFsE5PC1JhXjG2C
zhRwaFE+wrxhb+DXeYZLurUxMvnmtJsuu5P9Bw42h6Wke16xsbr/NBhKsC4ck4EOo/SBbpzTdZ1g
4wFyrhDsyArX5n67ribexhFUgk84h+Aiw6/GOQTi01Ih3QfG9WY19ChlcnYOjKgqsDqlJBgRFPOP
/Al4f4WocEk1yk7fYl/LF3J3I6OqN1Ls7sDNyOS6O377GVhsMrLCdUTYreBndsPPOjg0xijkP49Y
+s7/ifwykX5kov1HZomMTOr4V2YIFwCgh58Hg6i2ME4sK+S/Cc8BVKg0iKMzOMIX3aHrghuUmmfO
8D5K7mQJXoZR0qU5nryMFgokhZtj5ehRgZZXwT68M0C+i3syoYYDGhi4Bl4oXtKmtetYxbCJaZoZ
azFik4ZFbuabLqlTk9hWCg+AN4Sx81dglPIsHxpA01Bh3DqNQrccRwB661I3nWiIzeCFY8CwzQ1c
N3Y9gFpbx2RYd4mtxJ+LORr6exv6H5aBPvmQSDFRLbGVY5130FN/cQYLaEHQWtGkqvA7rXVDy+El
tPMuroQgNFqKf0KpHOD7AtVmxhf4gPfZGV3JUJcQ2oHzA/mxFoo+8SkdnH23x2wsaKzOWucVl/me
IZExWidxEKMozwKTdtbsf+yHiwrCxmlhFFQUUT3RQfbslAGpkC9xxuz9HwrQuJHTbbD9Btj3SL3S
3118LoeLvDq3cxgkCKzzkiOPXQjJUkWprYBzjiE4H4cOAldO1Z6xkePDx+yqqS9w/bwzZfGku0v1
hsrCS/ys791XiV7x1oWDBffAB3ekBFSXZ3RLwBcrjzcunlPhKJSCjrgS9rCqVC7zmo+1So2FX0Jh
md4upiQ7QJStz3ZZ0FVg9xF5yUmyknoZWi/p/Vk1lot/IOQCNrUwF8Zdh6APQx2ZeIP6/EASaTza
C5iiN+oFNoS2dtzZDoIj+9EBP+oI0T4ksFLp+3+nZNZ+5yF2y/PjDgfhRm/PaSBy/Mj+6ps6eBsV
0Tu/Fzxk1wG+16zhuTGNR4AWTDnSs+GeSHIE8V8N2Msbg+qfWiyRUwJco1+5Dfzzx9TcktCesWR3
228LTUKPOxdpDfdta3Cy56WOP1ROk0d7f+BnbqVIwAz1ecSX9f2JGbQRHFh5ZaCrvkvjh0UppRTn
iauNjGm1eJ45aduBfYG+qCKBjvvd0ZItaoQM76h5ZxDF/piew7UpfbUbzF04Hk7al+46zLFGbUwb
M2iub21paicRbEbmrTcbZiP+G6l0CM+SaPcL5bofQOJ/NFraRb30cRCQCySqz0FcW9syphvjsOzL
UkWnK3e0dIB5k4vcGtQz4nelSELCAQjC/EwjtLgIQQLs7hROgrPra85dIhVbo1CFdEf6LYwDT31a
JkjZ5qNoiGa4QBRRax5pZTpJS+Ndu/BhdQMtLn1hxMzpshMyDEFR6QLIhwSYWIXB9NK8fdNSXPEf
rdIu42RLx5ECZDzOrRWt5d56AWEE5kXYJi+BoCQpUy+/RNfsrHrrXS/wwD9SFr6h4PB2aKBm48YY
yveH00SH4+OVbsJ3+55IS9dYzAWlfVL6TWxMipMT2uKN7AomJnjyzXiA09lnhZVvWzpE9a72+UX+
fjRwjlFjHgiqHOpSOam1PcKYoUm14z6ADVOrhYWNJVZSJc+q5SqK6/CuBzdcTi5lOdN0FN+ZyO98
ozNnf3sjK4uaJN2XM86nqLJMiwE7W4KEHmkWhfgmDQ0iLxwXu6KYaMDUb9gZ5PeuHVVNwTjwipqB
h1m3Na0qC60P8VX1npN/QNZR2dVd2tUhjsnYNX6pRdrvBXs7x0PH/dfdZ6zEOJsu8PY3thxrNy7D
ERUr3ltcXAY0o+1tO309fA8kL08yNNcoF53n35LtUG2UVR/zMVWhtdVsHt66ikk2tZk3bW3+JrDZ
dIvap022P0RTGTuQYIH7eBs76biW4UQJCKn9kaXV4qJQhrIW1wPf2hFHuuZDAPnRpSSI/sdh6+Xk
SBvp3shWEVwNkeiOqoYHUYC5yEr1eUcNIARhfUSfRVduyOreQiBoGRy9sQFfVxfj2WVbCLyn/MQ9
hq9E6lvSmtR233yiw84iyOMvw1WKux8hzor7VKGUB5kLcm1+kO78oNRa5oJFH6gXdQGQICy1hdOw
3ElKPbQViuUQHTNeDfYuE6qo3v79CvPY0QSKYzUK69g4O7Cg3jm++cX0NCGoGmfYs6eAWGGlY2mm
IHqiog/a7DUixMmnWEdNB86tELdD1nhIPb656ebKcWbT5FGuq503U+vGW2G0n3UuHeYwUywfT3gy
XC1NOTrz3QH3m1jiTfcnb5lr4E8iq7hbMgEGm8Ggo8v7/orxFQCoaJHZxEbpHPE7NRWbUaXY8/kC
PUQ9gAxamqMlSqG2q/W0Jw3q7zpYANsm6aB9HNLDkwNFKBdwW28gy3w5cyXajJ0AvPC5yAUIHIbc
cjtc+Kkg2Di02GNcJqYHwsyxhmf9ao98QmMwhwR+8IXAy43gqcPJ2Ordhcvy72QEt0XWolNkV0fk
q2mibu9JFWThyIdRKDV9oeZ1Qn4wNolseUCZuklxdV+JksnZYTex7//rcqFv6RUAPRA4QK7//dYF
EhUkA1tSbxvpa6DXVB/r2m7ClqN7fiIxWyfVAIwicx++POMbp/K++6DkOUuqMytLUQX993ARKYfq
mG4YSjGCPsEGANBXRmdL4IJpV8nOKWWDI8Qgg+/P8xe+svb13+uj2KHdkemoXRZFG7kopZ8FcPSm
3c90mFF0E1/YFwimXzb5Q7l4F8zzEsqC0U9itieK2k4ubpKbuncGQ7x9oFq7Zky1gsiUxKJfSIzf
lrhRb1VFec/FvE0Bd7rjqy5dMZd4ipG4SNKSkZojwFKEwKprQW7tDhEO2OVtxbSKJ67LhcfZNX+j
Ku45J8lVFZke2deGVH2wNFZu47C0bAhuZ6zC6iNE8l4zy6+obnRnX7NFfBkDHLH2/2Zsvh/WH2+j
zdYYuFPoIJL3LHV0A7Q96iAXqTaMP4eM7RJq8KnZbjlRi9GFHCxHziAqFTVVyrJVIDz2k737hQqU
Sxf1rRmseU+OJ/0ElGGguYtGgda4fRtEZCMco7JLC/Z/TYf2HZoT1/2fB9c15UBxRqgECkEYOYbe
KXXGLUgifFT8OHcvxF7+AltJLRWKNkBjASzB2PsBll/f2ZfX1nCASUIYccE/D9dDBACgNChuOlaX
W0Z/A0h/kihhynOk79UekaFsnjLZm0DDRcNQnLFUrbygZiqWIPc5IoV1L0j7XII1DYnR73bGXRPm
RP5uB3FhuwrPL41Jo8F9+6KLhjKE1r48qRcLuJTcZGmLiKKyX6N9bkDPUXWCJfIfDhm1pt3PNVSB
PnduiWfGaXCiJ6Uvjt++1NLib0Ay9t5w96aQ9TYXzah0iTL1UkS+uI7lbF/Zt3Df8LKGra4IsbCV
SBScXBdaEcp+1HAoYBRGf9fw+FgKYDh60f+GZi9Z241nxwgP+A1GeUyem9DeiaD8WwzkAO0rJq2V
cW14EN8h2Cm5ea03kgxzT3KPf7coaX4mKyUTPPLyY0l98iFb40L/xzQF7y6q/ec0Cx/gQsY7111X
FvaAk2OzA60sKAnkrFZ4hex1AbmWub9dbTygIYpDRhY//KwGobMnoCfilrRvrcBcdanQWIHwjqxu
1ZVMGldehP75Dy9SLKENrpc8p9DFiBIV7cpmIPkHkODlhnFGyhGR+nssJx2BRI4JYw5ca+qDfdyI
JiCYl7ZbVRKEFR2zZzsY2iwsC0mayUbhNwrRpPkeKD/HqsXAAIrZK6W+ANE6MYMoDn0ZhWHkDAH0
Btwnw/jPbweXpqwQvfTmMAnjJZ2FUuSI3GHAd52ZHKEv5XGedW837egiP9xVy/QT90VXaCUbz3lW
EPsHe2Ko8nwmYbYkdqtLjeJeu0jbY6s7pQyI/CvhqG4SjsStt4EXoX8MXdKCOZ5RMaldKeAjwfgh
WTVW4wOhpUJlB5cgMy/GPi/n4D6+Srr7pXRcHwxOVETkVCUk71uIkDgMs9ZdoZkHcyfjlCkHzOCo
VCNu5tBVsjSEMGAs+/IZv33UOL8Zfu4piwbRts9CdZyAIXrgTa+3pPoWoOFKFnrlLobOC5XAoZmw
GI2f47IYObQ4tN5ko3rfgq6SUy46M9FRa9OofbtOcrRPWqkYdlDszz6d6tehk4PnMgFrKf9lvTi3
lvuFp48k5O1pYz2jvsPHdoDYvi23psBwutIxAoKTXPcwHzaRROxHY2dKnPriQxsWn5KOBcG9w+Og
+WpmsVz0tR5GaEWwwIPPRWZg0C1si+qLpDN7YHcNro8eERXHThcqEcd2iHMRgc+vyKVMbgGjfgcA
OKLugC3erJRYz+zWzj1AMLTQP8Av0j4PfaQSJsd+ywQBgR36k2SgT44Tgvp7rteaIGHR6yw0qLYa
rYZQ7aljEgQNq2fyoVXT+2cQBLLRgjEeqo5Pi6DLKzBSAd8MuWh+llllzQjDD6wpyfbpaGpLnFO3
U8LeSSk0YFKs6+ZlPUKFwj8osM4yAHUMjkM7DT+B2borRbZJ235IegcnTGDZM/lNsb4ikJUzt5uY
5AcN9Di6Po0zTZU0b8LGSX7diTzSprh+zv0Zl2R+Ff6np/X+V9c5Pt8Y8LTqiLc+1fZDMiyx4Wl7
7RcvmJZR9pZ34VnaagtwcbgS9PN5rgK7FqNKuadLazqWvTqMzmMYkXfgwc3DfUoEL1ofvuwz+mLu
aTr9vFQBwzkx7aG8WHq+DgB95vHrOGl53NAXA2KLb5Tbn6hU5ybQw/E9gmchMwL4+e7k+XucUjnk
wd1NmAN+TFpLpGncG7xZQxyVCJvJUJfvcMs1ZqBOQYE5jm3ScEY4IPFsAtO7SI1T0VmMC7CsF+Qj
NvQtHU5mXTSvSflHDfCwtXl5folth1x9z/63YKgxIr44KVQCAmKBwEAwy+7TdUZwtJ2bphknmYca
XogJqNc871Io4KL9w3B5GNcuIxiYe6eOSXzceQyqw4nsw2U05KtwtTZRMmEWTX1VmnzFrLo7O+s3
yO/rTQwiHsOw6A9eEQkg1yCdrcNavrK3uOAHYPqzG5Tu+7SEdYVPz+iM6dmGVT/FJSKAcererx/K
FkTkra4iMBfjVwmUS+abPOvsb1Y03+w06FxCNrISdyGwaxDWLu19o6gQoUO0QqdPUhJ499q84Lr5
m8KssXh8ChXtKDGNT1a899h41BsV4ePwb995CqlNzdwGT4SBrQn0UsiQWCJAk+ef0J4yFUfLFGSp
xm/gD7ZKAutneZwrugonCSkUhuBmF0gk7cCT71HUle+Wgy3XZGS8TAxYh+jW9tgNyTuLDsKAFFfz
sW0Wnmsbn+mEiUu1lCHe4OYd2pnfUquAgGzPUG8d9PmyHesQ7nkPOmbB4FOh5ugAKh1xFml0Jyet
VUCbpGDZoB9xUpJCSl+r1tYSW3TQrX3IJD8GtmJpUhnkc6OAySYdAxCGXdQWS6CF3NYkz95iKpCO
ldxE8iBBZ0kXO3XCiQRem+bLOHEfWFrJW9DmMuAZ/QZvegLd/vLXLTaFl0nQYk4U+m31ENiLX7u+
opEPQ4RGTONSboFBejJ2r+c0Mo49f2noH9Cj6KvLiW4CbgTpjEYCdNBU3CyicDhqCKE2I/b95jik
4PvTsQ5c0mCZ7Y19JUkX/kUVj46ZSrofXmmBvgHlYtZSudz18HZTPo2BByQGxhiNNNEHCWNpjmfS
gqsTinMlcI0dazJzp1tHraMiJf6zCdTSbgCLTiSBY07uWcOpHP6RgbpM6LQSmUgbE4FOX5vUfh6F
bDedm7HJ+a5RfimfVa14uerqSfis73H/Z3kn9U9wn6lPVWyHBr5tgfNkzrYLvSCM5IcfvLiCNXfw
3VTagRFSV1xgQGXP62Fy9rlYqrKGr/yzQtJ4QZZciKbdTsmvA0fcZ5cL/2b6T7zBhLiG8rcpq93s
BfFpR/zDQnTk+cqWQT9+WE5A1HLkNG0dGjqS2tMbRMMXOpjgrtXeFrgkxWds4q1ZMjk/glw67ZsI
eeGqJ8eCRPphGFu4+TD6AoIYX11VH8mN3tIdi7vrCMj0HWwRxLrcpivlrlyLHC+M4fE+IVNmdj1O
GGJTHHeV4iP5HYKwucPQZNgtFpNj/rliWhOlLo0m1iSNkDEk6Rwb/jehrpWFU8vNducyt+MULGsQ
PbaIDWSWbzvBQ7HEMLZc2Ex0itIAse+CVPkotclgJaJwH0YyVkOeLyfr/0p7UfvIykXuBzHYF0jJ
Kt39s1kOowwueKPHqwBrrr8x85MrCbf5mnTjCEbfuI/UAnKC6R2TT1pdXf7U7/yKyYJ8mI4Du2qi
/oqPdIFi7jl8E0cfPhKZS7VieClmBSxNrcOvtvob7RLM0L/heTaghbZ0PJYZyS4PqAyVlfOrIGSp
x9m1Sk6QEO+jLblcWxc8a7VCUS73vK1iRCAu4TvComFbKa0elCP0/O1J3KjBZ0ziYkvmeFKyA75Y
66VO+4svBGvv+R/vv0lgmA1Nr54SMlHYihvnVrLK/tmfsKUSw1NaKqs43kuisxxvzWFS5QUYttTK
b95OOItuXliRFdKvKxZWf/wbdgWcRhbWKl346xvJCzIEb2k/+8d0cWtxCj6DwZ1VgtdbVHl9KU3r
s26epHt3cggBaf0vyY2w3hmoO/OpHaxNYORXyxj4LTbOxhAbH5Oc9EIGjCYEh7c5UVDZ/u+3mAOz
YLJclCu6W4p5zwfniSrWlLqsvjfdH6XUkxHe7RotIxkRVjXTgvv+InYEgbc5ePXTW3C+qGgFcPrK
JSn2dXE7jpRCvnrKBoopTYw5eZ+CKoYhNw+Wq1qFzAvpaLleWGlGahMLpl56Lfu04er65ylgH53z
ZGeOV8wYk1VjHBFEUCXKJRrRPVSInUlbBlJewsx6+PG/YeWaATyAABiezYWtmio92qhkk5OMHNfb
KoJsfhjQq+ZcNesysST5duIht4n2gKhLMNUMkbTrPN1z+91/KKfGMgGMImhV7Y/fbrMS3oYHMWVu
xpDXjTnX9xsrZ/mSE9DE0j9spTP7hgNRiU1CD0kH4E3u1u1c+DgyLzNaITEAbFNh7Bm9OSq6t66+
FzxWSlHoq5P+RsBdoQ/asIYEb4to5B0ie+nqIccofumq0dLM6GjpESyA4cmtAMO+ewcktdHA5Ugm
l2ierfh5WzKv/wVTLuxZ7xjaCZoq/R1QzSEGrB0bJWzvRljzZ6E20+IaTx52f9bUGAayhap/V7Gz
lDsSxlkPAFFZWdsa6r48hYOH3cAdQ2TQL/w54B38r0r95geVzfZtDc8/wLLb6yRgV4e4A7eQA1fI
gSine1oFuiGvlEPkvz/s0ofZG4/mp529afGLwkX/UDkb4O/4EV5nDt2OCD1vEYD2VVe7lWKpfC5c
dauSo4BwzkWBP10TrAENYdeXeV/opP5C3EGZlNpbpZxaX2qQcofCOT3D7xuOSF9bC0PoSiPszo++
hyNppyYGfOOjFJdjkq1cufeZHUPcAoxKelb78jVvv5rjMSF5/IpumdGS3fyfIEbLiYGEru4jb0sz
KG2h1Y0JmOYM5iUaZ0KJxsTOLfW5NtHQn/WaG93fUpKydnD6HqwJ5LHRZi03ioA8H2a9nAbD0Qb4
WSyf21EFEcdGspexeKT9NBdij3zOoMUVLEa28VKC8JoNHoIBbxigRMQSCcmXKpv+YWpeh48MXH2F
hSqhJO1fe2R/GlYHTDwjP7xnx01vdnPQlbceINYNOimxYDAA6Pr8pWKmd3cijjJyvkdWVKlFh9Y8
4JXXsXpLs4Rrh0iX44lNQh1KhDdX7r5jX9i+FAxJYKw37YnSja4sDxhRuqsCV/fdOxiFkqFHktUH
dJQDJuwsyAHJWiLW05TCaSgDXDnx+k1hACLTrhZkcHtA1bj9KIB0J67jKmsbrbb6asr57eOgu2LO
mR8ELSRdrYrQA/qt8Wexz3BRQQfnd6d8nnA3Xh0RDXDvO7E/hTn/dUjn2NU9FJfhV4hm7DlrwG+j
OvuB+RBbrV38NsCI31B4OYGrmKQNTgcJlUQ0T7Wi2OjHr+cshHqegu2CSGrbd9Gh4GZ6Gyw45xsr
QJndutvnnYgbXrCRMSIvKwbbOyAq6mbFwPBo7jtaFQizARZsDL8XUe64Z81B3ufOBRoc+XAjXjBT
k7gaqe/ZbmkfJMCVAzLrI/djjWJtcFvq+Na3nE9eO+lbp8nZetf7RP20hFcZYvzr91h9NK3IoNhQ
s/cQ+q+3QiXk9fYemshWJFsStVQwLaO5vpeL3DBdpnoyy5UwmCV62ZQ55Ks7/8NWtWjdEeLKVr0R
T2GurX1RUGlDz7Ba2Ir1sOp1X9Vp9Jg/lqIcBQ462Sf6Qy4lwYEWe/6lMg2X9GplMRNkIFQCWweA
WI3kqAwEwDzqturH1MpeyJ6piZI37uWqUzPpsIgmFYDDWxr0KmoOCEomU6wMbOdszSrRALIMnWKq
fujmjbQY7t7m3uEnFyWDhvn3aLkHAfrQtXda4QPz8TvGcFkPpNz19NWFfgfqqNBwDf6VIy7jIoya
7OHGQTz3UyeALIgw4BR7siu7QIZrSZ+sUcs2DAyZ+ZJzF0dSUfa1hd1GM0CHX1GedBntomYJXe0u
I6Dwa5SMUjC1BTTe2jFTQx0Fkn3yi7EsHG2FVz7yJFhjp1o6NMJlUMWspyh9la97V3v3igIuOVim
5A2StjOhq1IhLgaZ9uLBAoQY9IZTLZci7MPaljG364Rj8yTSBVa3POZoNWa2Y7zPVhCBZf2mcCSg
QUJhWmlUjgd6QwdH20KKu2TwHC3wlxmXqjv3nRe4JnfV01bYdic1DecuI9Mfs99YcHjldBc1Pni9
sHQ312WSkZAobZui07WdL4+gCVMH1jZVsGOwp5ekmtDKerfXgUoflaEcA82DmnEVdTyxMCwzR1Qj
ytLq2Hi/xCidwrBnctuRruOIzyri3O5uHQW3rq29EReDQIMMFum6gI8FiUWvb8iPzDANTHE5Jk8f
/NVsFRCxwYYYSyldnLF9qWj1YAPn+M/543S+m9e+8Hj8os4xs4cHcDkVmSBh3K7rMLS1sBC1Y2m0
wfwesOyuDtvZa7eruJ/VHjW8Y4eNbmpdF27UGWGF/5LyI/vn94yfdhLLNivLa9d+yLd2zRxefxLb
0+WgxmbIMZrwCfD2HJ4B2fBcTedLZjKOyQ1cbcWj+6jIA5FA3V2HomEoRCHb9RVdR9wdpwThAfLT
3jVwHzwKyUOqtPToH4nXaE+YoRkXGo/al+w92jIacA2nQTNMECjLzTRaLrXelBSSU5jRSHa6NqVY
ioH045KwJd+2xsg6dIATZYxpG33p0FDEUh6b4vpiFlX1Rds+Jb4BxBlw6vOAjyi4mGvMzEIknLkN
wbShudfE/E2PRLoPUKiaZ/xCEyrREHZzP+/ah70CXqdlIkiXu/98l4bCOptIVczsp3XjklXzEoyZ
+HhvUk4qzjYDImCNMbn2C/pjWJ2Ous9FIZ2WGWHQeqq0Y7po4M9xzbOHkz4eq8/KZbWEKZwFp/Ss
DVHki7yWIw67E2tlqjRQgEWVtx0ramceSQ6VkjDdv21c2gko0o2gOFT4XkRTvKvGzaIUDEc72xa6
9mq6bjbKAEePFP66ezQamAio38m1nx088b1gDTlsENq0S2fIC7Z91OpSMH6j7PG48s8Cwd4VrwfP
ss8mPQRvLVjgpi2XMbgoyyymjKf7CcptzaACprQUUnLDv708GM9ZjHwSagIvYEErEEiwxFmjVGfZ
Hdfrpb7EvH5cX6d8FU8KXXyNd3mq+CX/CxHnoBgJ4cogRwa33rfU1lFS+2SlaS6rHIsK4YqA9Pu8
YOLnO9pOb3k7ctEpIsyztKEBE+gqs5nECkSkbBSVIv3X9qzsF0Qi+4P7k8pM7ibDOuk/5AUhcZKr
WqQTmvLjGz9cKWOe1cEVjYSc/cdydecM4nDQLCPT3X0v5KDeimyGQP1kTV563DSYBS8XwhFyjOM9
laURhi4DbbfFQ3Y3/GwP4uE0GZJP2ZtJALXmBYzdRSCp0oBRWIHbyhVaSiSMnX2hn8sARYC3f+jJ
UK7/MQcUp3GgbxRysGmD0M9SeVHgMT32Nl3RCSrRyW7JJc5zvwDAm7bK8/YQJpTGApkezavQv7K8
klEs0PBO8RKR7NTrTOcEdqBon7yRqmuOJJ/mhey33sC/SC7RjFDNZcxqMnLakevfapbBpowqoBi5
p1MO/vHDzD1gwFRwgO6AibEB2ZY1e2sphkeIYEoeWIuLzw6qYsh22fu0nOtLTk3bmkvTZKYnDTbL
cj3p8DwuZ5hZ1mHigPOLTo4lmVdn5IEAtFNqEsE7Pauco3axCuL4uLNMAiuGJWSvgUBAGz4KnLDd
SxKGdS2dtk5suamBmTOoTzoX7H6KxokC+6sEq78UZ68SIOApCTXT5JbdG2ItVrZVkXQQlk3pngFy
fJSc43ja1ccbcuv3Usv1QvrnZaKxxn929NBC6Pljw1uk+w5xtd+/5dQ4f37lh3LKrW2A5i0HMznQ
Q9n8VZx3pe8epW8jah3mbN/qocbwhFdDx5ITL35GNHcrK1yZcW2bXxSH3yIllj7ysx/uTTHQMHuy
0IpWncW6lFLa0UPovBbyZ/Z6HTed07hdIvJKc5Ue7fcWePasXQQnBG3kfNZFY+Vc1p9YzAnGsC3b
GMYxmMVzlu0cbcwyCRMWBo9GGVLtponciXcB3jj081YOOlXU1FB6C3X2a790bjQDNIJVlq7ybTHW
R0+cUCTvtyvlqaAs/CdjHAadQal3wiDs/Ra/DVoBniPikLtU+0cBKY0O4/+Wc71DwJ2l/iXFBVL0
r7dsB+7j+Z47c60XkB1XNFq2KDlSDFYM1qdknv2vIqtsIeQ/BrvXfsNsh1T9Uzkv/WU3gDK7sWx9
BrAKvtBbxiKbkE7cYWjpU53rfiXGxXSrTIo+ro6SuGAJce39Eim0xBnMjxZn16VKCq3rgNRUCrUf
KykKhRp0dSw2KxIwRovSb3LfoQnO8Qjh8ojbEbB03aeaAr6EQCcya0b+0KQdYg5lpVb1HLG0lKbM
lPKggElqlhjzSVPTYsGeHucPz27kGHbYDM5FAV6iBnTQoympmpykCCn3Mn9vwmYNp/zL+fiBr8ii
VSocxjxf4Qj7rP5VDZ6HmMRr+WQMCLHIUlb8VtdgwUGgZx+JoELY+X2P6bUmL+5ecLENbPo9cQn1
EtxWDxjRyoXUaueithHEViqHnMV8Vuo4YvbSmiR1VTSXT1PfyN88OgXSg41rUP2j/Oh1jtWHojiu
iFQHs8eF4u7L9YnkFVYiOpyO5kmj2W3G3D6a27Vmy9vxhu1AFv6H5tEdvw2jTvYvAvbFUBDt7Yjl
hkbHcgKDDf9QG6Gw4M8tvHRa9+21Shzz26JEpO3H1EYy6XnEmdPrkc1s9NDq6+kpAemQRtXUOjW7
trO3yyKjTiesGMR0ZZjawPBKxL66SaJp0lLxCHb1CWDrjgH/6OfmuX4JPycrMRKKub9KuK88BQvt
BmLSHKTmMvUOYK7ytXo+o3cFL1Sdu3ekmLD5O0nO54IbAEW5rMri6MK2JCtT9yvJTFm6vHhc58vT
VlOQISfpWU34Ip9vZi1gIkgt5mGxoCUY0XEJXfyll8co4SOX/888jZZhBGH4knSv5N3hZt7G7zI7
RgCMmRu9TeadF7+gnxJPV1eqO4ciBcfJrfQIYR0AcRtKuvxiZxFnUECd/6jg2VpvDDCQL/0PmM+G
IpflJjm3W2DgsuwzAAS3uDeo4vKh0BEFbcu06KKsj8ByEBvadh91cRUKFzuP/UqkhSKAI51n9wvi
yhtLLbQOL0P6jxRFd+ry+TWP722LkJB4v4ZRGaBY8v3zK4MZqCbLQavee8hDojYPCYLg/sARYBHF
ApGRn9sl4xWMBd8SACIYfNtI1MVtW4IJ3y2Yo7QCSIS5yhppDWI09kaDGc8sAuqDrHJIMCZHIm+5
ON4mZe13XOys9HDn39SABXyXV0cCehERsNDObfIf0RzJUTxZWeJbsj3Y/XQtvBAAybEglqcUC7nK
yaXIB50l4onH5MSTe69LQdGc0cFPu67SUpNimMDSc9YEnJCyFeCijr8JNtDVCsYOhsX6VKKRjHsy
k3G+nFrjKX4/ZbFTgwLT2MobAnrfuUB5CO57OhIr+OduKgcOHbfVh6s2K/ij0cVY4kgBCwkAFFw0
Qs3XCDudHkmM+n8lQrGZmexO5apIC7m2nltgUecsmrNmtmdnhoFm8NvymjsIStcA2cLDc/kiUOZ6
LW3gnF1mJpMfwIMYWfKSN1A4D7Vvp86NbGMnSP8IxbEuJBQT0WzjS/uN6E33PCe9pJjx7WyZVQQj
UGr7FFDpvqAI8Uw7Oi1nBUJz7xjsUsGxhcFiI0zczons7Fa1LZUtJubVOTKRPIB+1Z3Gc+4KXcxd
+OZErfpgj4Qoue9iVRo13ljjIXxTK42ia1IjsncTo3avgxtOwTp4kIJD0Znh8+ayHgz5AI+II3iC
fH64+T8RXzKJT/udaKXI3ydszzgQzE9YrtyeBP2VyHeUvmAdw4OuYSZYLvwCxR8REegU/Ue1qJZ1
ter7l+hvz/dDMqj9eH6iTfCCMihV7wiruVY0Qr3S1f6vzN5hEqiHQRv5r7uNqi+pgr9wqRZcQRMi
vdt0wGjq8voHpLNO4LKZNGgLXFeABrDpCthzEZIz7M9+wRmJXLqg2kH6WMCL2lU7yJ+nPToCFUPz
6tWy74un00CdwiaDgUbGioq3kodKX24vXLL8A6eDdec1QyRM7LfdfhWw+kSRM8jqoB0OiZTZBZHc
RgXOu35KmkbqzUi41tebpLY8Z6H9N3qkZkNL0BWLhbdCffAwdFU2IXMgsyTVmWhYooLLVnWag4l6
ijAJ4oAtbVHUrErWa/l4znSXORyysJ2NJy4usyAjNjFe6CXB0MUZA+Punnb0OfGYVd1BpcySwohv
uQFpCmC5sGhScHLcVuRulbXINl9lvMt3N0H7j41LsvlC/QjB5oI2G0Sc183yHssw7WRnCFQEJlw/
B/Kh30oOaEXicj4v6ID1F1iPS+6+uIuQbe/kEpweCXyJKqcxUWi7prUcmBgIZzZSltoDNpFz7AIz
JE66bOQFgjR5H/fjabGb0HQgEdlaqolxvuyM1f0/NJn83Fm+jYsg5daMzvWh/sD78E5Ogi/9WJYt
RmlQfKCQoYwMDX4cTDYf9PV3s4SVIgGXvmV287ysgYQEJeTAHcOP8atqH1lc0HA4LVDE0FLt1IcD
T7X0GtiucsSK6L9GOq6+jO8rJFsXjVTL/VYOdbPqGCmOBhb6suPfNSLaEUf7H73XBFuPXhnFkNg0
LRmmGB4V4D+mFRByKvvV3AOB90f0tB3LBvLnU0282PPG8844ctmmZePKhOpbfTQ36hJ8wV8ZCfZj
6qtxrRvBqeBuKbVAAO6ib5h5pYGc4f9sZ1rYwwf3DiM7aNUIp1JHMzIJzQtg8EMloZ/WTo+bUCPK
ogj3pblVgUsPD3OQFsrdVTsL9oefb4/LF94p+78b6GYqcnHqrX0R86ffwQA+c5fqUkXNP3ydHbZD
G64h1EuOAI1STvcL9muN1sDYqhDOZsDW/geYEuJ4vUeWceYpFjhMzQgIczBwJhkPjmlcy1QTO5HR
W0nKI09KlrTbRjm2MlFDIE5ODw6l1kkDh5nYMMkmaTak6dysWoHpElbrckhEwYGclF4Ra9rUrthY
sDz7uEpYb3XToJVs1/3ZNpkJFzv7Jxrhb1tysvwnBpfsVCQwZeSrUhEYpNNWRpEUPzXxcE+Dpziw
9PR0NWLcuNyubWGpOkbMOv9klibguWzvkWTkA+RlBAXnk8X/FDVRLQxnAqmZ9arW9o5Qfu9mEPpw
TN9CwVGNslnwQ2PYJP6eeJhIEEDNiKMhzzrWpEbBZJzyZR/XCaZS+fDODFRlyqXgNzJxXnzdKeci
gnk2BQX31pjxQJHgk82/rpqo8ylJ9Yz5387ejCTlGCcf9mdhL7+wavMDBO70i1lKkm930eC5xaQH
cTBoUNUoh7rRSkioVYlUR6jG4krP3dJDyLn/6atIV78czUel+FVHrnsFQpJTkl8pGwOHT1qzqh61
3W4PONofXIanHuKyMmHrEMzTzpxgVSVT5pCPRublJrWTmBH+xQG1oYhvoCeRVz97hG8aMV2OpZrq
0NLv1hrtxl1rZKQ+VgL85ig/GVEXudD3gZ8eqLynYXCQNa0v1dYyh0cZK6+OfhEqi1hvRrtVgYUP
qxwMrgAN1WalkDBiYzqbGziuxL5U1+okOwToo4/NtWmGsQKUK1k6JVp6rjx7YyfXLyXDV9wg7BLo
Sm/7ud8Ee2FCIPptNGAK95gf6hJqKmyrSjTKmhO7nN2ZsFvs44TBRX2nJ282Q6ylm8H1UwPZth1c
U0IGYnTUdiDETFBcUtiG3EiyaR/AzoNcQD8WxkXoU48+rdn7kQVQULyqJuGUhXh+UvUtCmNKVun6
eDOrjGhjvMsSRaASPD7HIgR2241fBBDpuY9r/kxl8VdfZRtJc5NvgA1xIWHh0VtHKAzlBQEJD3EV
VZG5opsakDRq75e8xufZyTVi6eQK0FO8ldl1Nn64nVYR7bg3Pv0/D5PhTmCoKx+9LNx+0qNCKJ9X
MYJ3Nc5oA7aqFd6/efr+JMoXL+5x68OjmcYYFg9+0kydlMiW1ByTCCnNAA66GtOBD4BC33Uud+QC
8j31E3uzqaofx7OZzWCpIgQl8Vv8mgh9C3/PcBSSN3zm6pH3AuEoND41sJs0pmvypuh2FNIirEwO
8RHowr4/FFkPWeA5/oJQLy11Qcv/2obvehCXQD6w1J3R35FM5Ccykz0bhHHhWlAuEWpQTW1XUHme
7EG52W9NVmliodTGWF+0Oczrb2hyL4HbNw6GH5s1PxthKAi+vqZaBYM0pNtzRnefDU53lY2vUzid
3CBbYyhSni/Ank/xYZGE530x0Xe/sqXxcHaLYSINnlrOowewClH//A9Qy/AiKPaO8v4zZcVCz1KK
gn2rCaLkOALTkCG9xpxabVSGM7B6t14DCLrL9ynq1ffhtPrViopbYWQQ0zPw5Ff9cDf+xbEzwMAS
mE3gPNgtXZXqSCgYqDU0d32PBiQeGESwtItaIn6QUOR3nky3Q9r/BCo3nPYIiigz0nrGjev/yRaT
ykzdadg7F7TuiGBYr9mQpbjQNi/1SSg6VMI7DkXX5HSEU7neR5Mu8Zh/ZURwG+5gJA8PrLK/ipfB
ey+1DlvOn25KVnjDksuhkA2nFd9TW7LCGYU3EVWWC0RaPH+XUTTXfjAdiBy4RpMVVRf8Lb8wkwol
Gq1Y3I493GRIwnDeQdNndNIqcBSeHxknkxjJi5eB7fXp2wXO7+sXHuzFwzv23LtbHUK3hX+t7rvS
Hyrpp3ySH9+BB208RG+aQ4XhIAFn5Gt9DTbip1khBpBljKo8DSOc2dFc01gvBgaO151X7dD7vb13
4NeZi7N3M06I4i6eTJLom18oegZnNx0Wq7S7wQVInN21jOzuUrsSc4z8XElrKuIkosh92I8rKmCB
tiRQCSVoQM7Ps+XyrZi8WIGyqQtobcCu85orBRgUr07O75t41mumZ+R2CnW50UjhE3Ct4YJe7VAL
8VVe5L40GusDTKWVsEDinVrhylsfs0h0jkuixo4wcqO3WB1+/tggLryp/bNwP5yTvr9bCPEOyrQ2
gH7XBzNg3evGVwxUffhm7beRol9tLXG1GX4Fibl5UF/QSXaUIkeWOM82TAoS6p8LJf5q6isK196n
+4N1wMg7D6o+Nr6GwpzWX3kbz4Hdio/XOjMCHU89uKTb4AynNnJ959ew8UGwnwG4gMqoRBddFKld
aDZ2D4wixHeMgIwun0LVQB9BUrbXRyhh3wl/hPhw7ng//3XJscnnm1Hq14UAwBwsf3h/68K6TqFe
t6dqZwpPij8msicrSiekzJ55LOo95Z2rEwYBq+S7UKUHf96woP+RB5Mf3XbcM/sno15CStfXqNqq
NQ0nj8PsR1Xf81ajCu5bicJMVp3SS4yvVWuiczY8pfbOtWToOvJb5jvGItsZqaTf9oow27xZrwFM
QyYq3C86ncwI/tKifcn2bxqePpIGw9cYEQoOVq4s6NvqMpsNh/RhR95TINNVNPyjGjE+Y8NsaL9G
E1ahpr8l7vuDApxCxUFlDsYbYxSvg6QP5+5w6b289EKx6cpGwAt8vKQkTkjOrREh2iK9hhp2tr9J
a/MtO1UqBxdsIvmTUZgNjzOELqyBJDHZWTTHy5fwv4AptWmcUoJWaol9IpQtwY506XwsO0ZwVugq
Mh/dZ9UhAoyJWnHySkKq5kYn2dW5jYvVSb+6P7j7YyurjfzWdsKXYYH55cQZuZKDHlSH92/G0oYU
Rda7tKhnShgqDJK6ckwmfuPYpNIrQFQn+Vq4CfnTr6DWMCLgdHMZSgINz8K1QlrCNbZtYE/qWj01
5lQ/uAG6jrBEV+UL4wpIP5b6A9Xkme7qMLeU5edsnbqdS6XIyfeTgfZf/dPuIGQWJRz2SiZQMZaT
eWzoH2aiIesaQxVgKixMJ5o0LwQ6TkvPN5JxC13Nyt0tvc6RcKu/PJSfvOSKuR83zNmwTuF85VoQ
zstUWGT72zSW2O8iB6+qoL/uhXswVKXH8Xq/SlGmDseuB4k0JcKV+inbCKnO6jpqc6MgWJAft0Zd
Ck6NIUufuXgP6/Yt5G4JQnXPzb5LnjPLL1t73+tBBB3Lkcz3hI0E6VcS25iRPfnWR0xjkxbgysTZ
PAnlXXFMmlVcZHcT8L5QDlIx6NbNCAJQ6jB2QZ3KLSSJwfAAVmsxthlvhJ7iKVByDPs5hVJwFxZb
VevIfaHocaG/1x0n5/ggo6K5RtbQ7+yZO8N4hH4UZbo7jGqrt1AAmiE+uJvD46A7rIpJaiSH7feg
sZ5TtO8V4axWR6/4GKuaKqBUQTSuVwLuU4LyHnBnj7WuOVYq8s+KUPl8dkTtzCo3P/M6EVraLjWq
ZocbQg2R2lAexP9yPtp3o7eGO7BwpKmQOTRjVFQGs0Hpxw5fRUAsUcL4IccuuafnAnl/P70gM6g1
cGeh+ayWo3xVzHGjXkE5I6uIGEaKud6RjK8pezOpMxTyQgtq6RPsk8hxK98yLzvLkQh8p3Dmq89R
9JNDeJsavUrPnJjhyT6j30NuhLo/tKqJrE5FCUfwBU3evDsinAf8Pf6zG0DRDWEjNWDbIojCLeQo
WPmxF48Egzt97eIzohFPZvQCgA2unkRGgnfUzppUlIEgWQV7PX4gwfK//lEO+m/EDlIuer2Tdkwa
uw311iBmPgeA6t34GBS6i4JjKmhA7MEEXQR2TSONWZHFnVvdAo9wFLr/y32n5I7BHmOw49oXhpH9
MyUpPC4dikAsiskwhjHAMiIFJY2ERAj1Un0jdUls4VM0oDLmUNhJ4O5HCcF5UtVpyY/oIsd5Khl2
yAk0NkGBN9gSlG8VZ3HepNeMRoUbJcH+rmATRioYBU4SIPiB+ZsMtMhq79y6JCm5YVTPCVVkk8Ck
VPnoS/qHd+bbdbPd5wHAmu88BImulKI1MSH+wGot4FySR8cSMXPPpJ/MQ8UvRrqfi4CAt9QucCmw
i1yuoy0OzO5SdPJgO7VzYGCTgFSvmq6uUI6/hrZldzm7J+k5RBpIZGT8j0vJKPIyX6RleWSBZT5x
phjAaHlFVITYbAxV0yeHz89oQC7x9udI160fcrCS0pkU4KgFumbOA1bZKrBPFw4V21zURXx1khe1
xhIzsUiKqxM73I7kaCASIpBbS0kuv5t6YqMisxKrBX+S778griKeOFm58giB6gF4taZPuXyVrgjL
guYmg2vjnuV0pRMQOMQle/wp+yr5gxgawnKq1mMOK9DfWP/ricmHtd7ocIqwGGNpOGHoVaExBka6
OvxgjRpTBoFa5kiVr551/Rk5ZD7f1jOOjXlE9+jqmGce1MdoSai1zzTEyaXcT/f5eB4ZpUuyD28w
ujCgfaFneJbTNP/x/CJQbhxl1/QrfcHRwyPI2z4fzb+fmToopVsw9mbWAhFRmup+/yx+PbgB1k11
Bpn+YbAyCaOwQFeMfj/8yniiCZrUskAYMsOqxuR6SLgvlLHathCUejpRKVAP+ZVauRsuF9gIoHli
ssbA1hshxohfqq9B1/I7W8A3KA4z3yHiaumF528GHADIx94XkYjfZbf9q22iTAioy6md277DEMB4
eqCu4MMjDautj2pTGRDoQvZ+zJwRyAZyLfjgUoKRdQFOCUl9/u/1CG+KzNTPdmEtPKWILboUXEJY
mArm5nqVkLoFn+f/YM0lRD1rR3gnn9FW0d4X89igXonY5FLU1jK1di83uJRf9RMwzF0yxRdD86GJ
q1CK5SGsSQWg4OIwpwBWveCAkFvN/GeGwDZ0Ps/GCY8yGss31541Sr9qpfdhtIswXlfsUm7XY9uN
0j+v/8Bk2J8zzurlEvS1c367lNOl2lDgwTR+rUwrLYCP968UaDSH0LD2VNMhLZBv7sdIIUyvJDs4
dSKt1vswGG8JUjsAzn1EdvKldzHZyXyr9qcwbrdDIrFHouRdkfws0hlhPkp1VjJf13t7qyt/Cb+m
JRU2jLCynDsF9lpkvcN8OlPWpp3m/nBwp3tt6PdeffmRiOM6kGNyd3vukeLyqddQmMaaZTwzzS3Y
XgE/nN/bi5F2F73TaTUrbMz5lHqSfsLW11Oj3Ev723Mc94osFxPXUYpMKDz2wuXoH1p031ioDdLx
/iKVWhA81GLc6XvkZ1JJmHIC3Bc4nNbhMK3Netr954//L3pKgjL2F+1h5dNhhSeGVFrr4armMYCO
qBnSV9cKxJ4GSF5DQffyKPSydG3SrW1aEGGyMviX7gCmsT3C4ZyJrDlmVDOLktiMFhVJ14ZCl6Kk
jcJwW/irGphI+iXQenOhFDAL1+cBrOW4KRyZ5t/chxtsIghv1o3pIEynZ4QHhRCld35bfNLaOkll
7GnRQ8kWnR7Aq7JQyBAm/nQe+WbI57GS+212bYEZVlHGgVctBc+nMJlQED+zO1sFFRBYSuWxeroi
I4n8Pc2Z1hr8WNxxFKWuwbMNOV6OOvh+pBUIBxw2sYK9SQRoG7dDtcwmaVRzYFys1syYa6uN/JJ1
YyxRT6/+0ToEyPN2fWKDcN8yu3fJShJhQ/jyx8Rd8O60bPi3How2Y5M0ZmgJS/sR6HSssKdLzbfK
VHU9kT9YhQw/7PhrjqKwZnCEv10/t7c4vpQPUmmvPIM37HUF58XgHTqw8ec96dXoahbw0z+sWUDi
QZqkIdILYxzSYPZm+ctmEiKsCEXvoaQI6lboq+g3rzVqnnCgCDmCanMhG24LvVl398+A4DeRVV0L
TRZHCKolA6iwGpXpErPCiC6WL/9EI+xP194wr60zFh4OQ04z2SPp7mlxJu3sDYB7LubD+GksSd7v
EI9/udq9LR89zdzK9MkghsLVfhsJQ8v8FKNGfXlcXmfgEbXiaOoQJ/v6XlDQM8X2z4zyBuKfssp2
m0SURPnlV3gJfIcWRp3uPsccQ9HR2JLTYdyPkYv2L5xJiGQ1LjnTWR19EfjTMrZxOHapYIZ9KAJ0
Ap5xBHz9676dl+8ZM4a28Qxp+SRBEPuZsV/QCkFz23yAMlqlnoJKBZ+t/MNdM+FsLEg9DJIlCiCu
XIDRyBaIJGtlJtQkFkPdr+ML4VJj4XhMA8+XFAWqiNh1zNZ0Ck4BpBeSNvd/SYhKW87IuvA2/qjV
XpF8ezFoeKTSrx3PCaAcG6UnGrJs4yq2+NEqrTqPHiEXtEMiqlq6WUhgNJyxGPdiL2UjWh6PqYre
szYkWK7fgjqU5BDx3ZWRhBsciMwtky3tVMNLQvtx8VBF5IXDJpxfpbV0knHi686WW1YiTBjdtjqU
P+EQ4ll+6hd8EXOdcvFungnNPIts019BC1WNKqAQIgj1cOhD5gakTcUj27TAoouN+XvHvq2bBa/9
YLtD3IYvI43mCpilUPEyzIS7ErlgjKmMLXPTma7Yn/R7z/c8BEClDMPma4j87rid8OeKcSiRe3jy
mzE37z8ud+6m/TVfzmgMZy6Eo4PndOiUPrUHgQMjhkvz7gn+sRyyOuSv7e7hYRRWHvr4Aujmfw1W
hxCQhYqDJSMc8TcXNnraWN5REG6IwnFJYIt0RyfvyHFfsH3VvWAcnE9PxTHOKvE/xnaEYIgwOayU
zuDCN/obkrUWvCvqZ5MVj6MGyIU6Ns8lv8nG/sfcFVrBKewBYHluJx2aY+FLuCSqG6zK0bOmlwSP
EiDIvjuW5Fx5gH/1WGSJ389tPqnD/luNXILhL4WUC/kB1lwNdS2A0fIT5mvdbqEElegYfdzfQl67
2IA0mk6KcyCk11pZGBLFFVgyIT3BPoBAZmfnYUuQkGHAvtY0wxD1BO+6Zk2Db4Ar9VZThGwCz7YL
Mmvr95d+stPoLP3adcKguU43q7BLSn/auImMp+8BqRaYI9ZZAlz/SN+EoATDdeaoSEdliRs3ESFe
OV0nfi2llUUIlbAyhHFfNz8QGaCFC555uYIKLGbInPweWpGMTr+LF9VicpLL2iVPxFy6p7XAdveY
94YEbn6+Hbd8rRLCDuYWQwUvJN6CRfqnrJ4T+d6TLV8ZllrMCoNJxyV3V39Y8islEx8BKZNNKlM8
uDPf7Q6QbdpZUK44ZWZHOELLsiE0CWrnahGL1OHJuMu3EeA9bZ2t1BkQzZhrcknhTXhawFuAuRNr
+zSc2YOHLbcTy1g2iVAMKpjYvu+uyawckFNwQgXf4n320GUkjLUbehnpZo3Ar5Gz5hotUVQQeRyk
IhTgHPyAKXvChz/r/bGAbyWYW3lH9eMXGgDZIROiPk/HRfalHXRxdKjiUVoQrUezOVL5ugArCJfA
mAMzdnNBHXNjwqMy+cTvad4wKBcJamLf1U2lhTvQfKh9rolzCz+oN2NRJOZyrXdF7Pta2YvbU2l/
5SvDsptYbA8uMwOI2XY46BQGXhQTJ8/CByMH0U0eU2zEjTgaoI1dslIJ6RjwoHCd+0UIqs05WK/A
i6vgQZ7NPCMY7h7Z6TP8hGqQVb4QGAkCD3Lfaug5JGuYy6gu4W11MhYEWVecBt6/VH3eF0eraw8Y
FI15pd5hH4dMP6IS7wPdhLBkKHjwAwyFkMmcz0gFTDPShXJ5X/hsRGrl6+z/qtFJX8AVMbclMhdU
9qvSZfMgD9H9Rh76NkBaxuF02jSsfnULPK0SANfaFlk+we9Es3k2ZIf945efEFGJTEao5PWUB5+b
hQ7iklBcrZdwP2ik5+ECpyU7wDsbYin6aIJ61e9NKceSsTUoIA/sDk13jpAUJ/c4Yu/WkAkElStg
LZQ5tJVfwqJbhOfX5da+8TdIInq0HhlSdVyEO/VBDiJ/0oryfK/2pm+qCsz8ZtNI3L9vZAKB5ADu
2sb04r9fO3VDSppH9jRbd54jqLRgSiQFht7ZjQ4Znc2DSzPKlozM3o7iDPHpUOYGxwLbXUpgSwbE
UF8Ig1xKBBEBeCcAjgr3zd4OuHXOX8I6k5cCfJ2Wf4vnV7tNJwavjBa58HgQ0lgqqe1zqPMwzoHk
ufXw6mBOhK5LArUB2HxkRh75WroXeqYSP7IPWEs0Td7gYmRJrw+jozu7mWiLcMiO9QShYOhxa/p+
f5OtyArAB/npWIZWpoj/2CpScC+EN1i9phWHhOSJK/Bo8aQlsL1K5a/BkERERB3BL7vQs977XLr4
L9nFcB8ErObWKVCqfvGCtgdy0N/hF7Jvwx7H1Tcpt7PzwtNA5YJyPOczcrm0EoKQeOQ37rBwrEIh
d9ZR+8ihZbv7RTgmo3CpZtafFZUo5mVMr9smtT3QTj5Y/n0aixrOeS/av/zxRwWfsxC2SB+fIFMD
CoY9Jy7SdHHOye1PoDICONzTKYgaBOtdL/U6oZ4BFkUKgi+2ZAModiAwOlnq/fPJtUb8jlNb1KOp
3cZAV7BBVYkVE9Kp4c8fJxn0lPymHOvkvACpGsmdAetAypORMsxMxD6YpvJKIpYQmnpb5nV0tHbC
alZCJ3jJJt2FHt9xbIAvdpNGU8fEjZmWMzyE+eEc3Rn08UfqJmBLokEfM8SS8Gm0et6PyOTP/xyD
n2Ru0vWDbzbzoFJJFCsMc49EkIWHZvKVV1ZPedUyGILQa8GmexuP4bb3DYkPh7lEvIMMws1ysFuZ
hbx7VQMD0QZGh6pPSYy5rmNMSXpeWLl1vi2l1MeZY09qjsURN3kLFtO2hpdqvTGMi4xSD+d+3/pH
4f4rPvzZMYBFRP1g2/erVEbdQ4pvA/JCieaIjSGc1nRccWlI+yDlDDWXC+8PcDfKAL4rm9ClFenH
Qg8JnFJDW6PiBIrk27/UsQ4uFLZ16L6JtFa53Bmdl4180AVBhF3NzUwSeJb7IDfIg2kmSg/ngG7z
qLXtjvKCWI73YIumad7ZIl73VcD91G9nUQmNsWPZUgOhgMTBTpFYdZLmcWhLZfAJ4S1/iD3Qugok
G1sJiQwEvFr9UNq+qKJ2mXP+8yrax/1NAXQfI35XHd8PvdYujtuEoJwpF4zSbMPVgD+xADGzd793
45giELzaweDCQ/fs2Jgjyaqp2mLjn8gF0gNyl7fYB7BtOOp4C8Q1NO16tu3W43qc+beXJ6r9MkXn
JKolp+7VrpR/ag88puOT0/OoO+s/hN8EyEzJ8r0X91yc+5Xl48yuFfhylAbVoM8KRwNThFa31xHa
glsfd6fTLqRHisOOv8fyv+dFWsdk5QEU8nO7r24MECRHIZpnX9iJ6dxgZnyyQxRFvsFa0ahDrExi
pW6aGpVbWYuPM+SGe5xwYD7/pojQPAwetNe4Y7N2xNEy/ihj/vIcBzmcZz9OmMaRBNSBCeeryv7r
R1wX8+Wa7nU0DWD84xE9OlvHVNVtUPxzhka5KEE828QD0QrmJBxHJyT8wSH9eVlhN//ZVDX8Qmd1
11GrIRCa8s8SCjVMynAJ0V36/g92ltMCVkyUXBV+LKL/MHvpN3hwWw0q66/W1QbnPPQzSgmtBFeC
xmRmC88fFq0GXMPfWI01ezDBUJ8DBk7DZmxnCyGE9W6khTdj5UoWt50wGFhKf760Tgfqo01nzGfX
r2Cm1+hcye47cJUEqieLLz83d5Xxc6TtQ6dkRRTOtAIrA16+EiL76u4rKifEUyPEhYK7s2WZeSaV
wRpnYo2qSKqqckO/e6fwDqWdr90p5qi2G0OZJMX/I8qtPShKYJyEr8JvyrM0BkMBdxRJdjue5D7n
xhlnHHw2/5tZzWkqek8RAzz9VDaIFpnV12OJckfQwlUjFaZDIJ3B7VypyCpT1lzTfxNJpBxZfAsZ
rI92tloidHDt/d9TrxFxwSBhNMBa8Il1kFqNKVi8B430Gx+c2kuP5lxPFoIkyroFuBc2NNKTqb1s
ck8Aiw9XDanU7Wll/2G708pirjg8CH6mmqmcROC1PzuDDjxz+NWpUtDl/aw37SVC1ZiMe6s1LM2+
w2cBfL/Zem5hzuSI/YjrtDWQxWGkcTPSOGXgCyxg7LzGC/RmZdfx/K/24FZ5/N3NNTpkc8J4ZBEh
5HMd2vCZIcRep6tfQ1VFBVqDBl48h1H5x82Vfqmuxvy4sIK98C4RlAyE924jsB1yZMA+CZD3dQol
iHlvMX+WIo/dxJTedf/FJXtEVfEkV3qkB3QznGNTPt35Fm0MkThaPm0pJrRauKRncevIT1nip5ul
mfcRHc3+CdE0keyT/lCvA7LEUUomPrsN3LDHGFrhYFV7KIloboUQ+y4cyasKNgTJ9WtWViQktlNI
yJLH0Y3mEC1QGslQABr+Q1G0v+4RwRw41GngSVFf7Hx2Ch/uWY5725OBBF8yxlXXx8CQWFz7xpgS
6QEBFzWv10gFgP7FyJKRoJF8bWzCOPvo1D2QcQV0UXpPKmvMPLhq9KD8tL62Hib9aI66mVVSysYg
Wlp23WYEAOO1UJtTPpKKRhnSf7C33PBAgBnsN728IAuqwuhZcgGUTE+LgUs8MmMa8B/DgkhrPlAP
c3RHoAeM9M6MbzsRx+BiY/5gdinBQV7dwODGjTFZwWznDmyNfD4cwWtND8XuV1YVqAunZ7pJbbIB
4m3whqgBEY8VQgeZcJtr9Ll6hILkXrNaowI4OWn1Tf3GDfjfa9eByfHcoN5mPw33EICXW9LoSe2R
WcVJx6sDjaEwFFCCW+krUDgLrTqawtPoMgHffe7JTnTenOb7kXguzp7ukFW0MruqrVpUgT22smup
WEg1PYYym+FjM5h+BKEOp00itkTkc0Bva9DZcW8jTXr9kSk5pn8otO7/V2A4eZaJerrCmpYL/zyG
CozfaqV0tUg8cguaK81gjPCDMvJqXearNwNXK8krj6yEGF9insQCu8HO6JMilrJiV/5bguFJ5fIU
P1PMIre4rLIhDvuHL3a9I15x5N+SmXx+ijphAoX/NqoZQuB2d/GPb8r3p5O2CHRAd6Ux0v3Oc3G3
BbSFE9U3zgg+AqCkZVUg6vyt/vkHBGLN+TiIR4KgFW0z5FtdHgE0/CVhoMBJgc7Z36jHSSM4BwZx
TD6Xij4TcS0zSHobVnburutDeeJEg7de4xFhfGZxAv8gAYH7PKurFGIX+GWVOVvamn0DWQhR1s3d
JZ4KzvObtcnCXzuGG9ySYcHwUfrogzzP7zioMF5RhLr87nmeHL41B2yf20O57tXyfSYHoij+2/DA
2K0pR6ObwazltyiYyt3Thy866DQeUsD2k/ZCvPIM2lSCcwtfjTT6FONKoeKA/XkKntr9lR9rdB14
rcmZylQshEY+gx6juRG/mzLCo9Vuh/gYwIZ8kR2XJrA2J7KfS6ZDcys2/curDQq1TvzHNAQ1Qdng
IJ1DGddxlmugirSIi1nARXUUiNdMN70WwaV/gJJcbWVTHtigpu/vrCRt2h/hQO/1M1mrLyDIvclo
xnWhs5SBEe6ndL9bd+OB8TRxc2i3dAz232RwIFiPX5/r22Gku/ZPOFGlAB2hvs5zETfJiclz3R+W
Ls1s02co6kF0/RQ1f8+GJ36KzA+Ypcqvswrfcp4NBP1bx3w0VCj9lEHJktlbb0As1VOUmCWRvjY+
ip05GVUVKpBXUdu26K6IqcGjddp7WcvPVdQsALp1n+68NoEYk9jCNndRC0ciVe0rh9ey3yPSdWCv
OKbEOQfZ2FmJ+/uXp1p9P9n4Md2rGK7nTjYLUDOIDZDU4BqfKLiwiepc+MXxnnQBuuZKuzDHTLY5
Uju6N8EmXsO3RGrbVKTGQvjgPgYgIf4C9LQmdia98Q606ee6pUIzcRYT+ENcE0aC4NMVnmLggxfh
Jf/erJwCz7bsu/qiUVPfmO5qveAeJzd7fM7pXkYhljdcZhm5T4qHuyyJr3ESejdmHr0+7zvTvAux
6Ci1nB9CMpra3CaQUpSCMopTf69JTVgD3UX3/vAuTmVucky/QK+rByocH4iCZAN1qwQReA4Vogxo
j8HINP/pf4UpAxXyxTRGDZ5yPChlZis1Z7r8eImNegG5x5C30gunnrbRY1+jMs7IUzVEgtXfpX80
hxX+OrJwOqmQ5T6BHGZsWC07Wd3PR6AWhg5IDIUHL84RC0Ler5x8ORgyZwzw62mGANXsiUQ2qPbO
AnpQi0Oe3r8zfeXZrKuZOXNQSWux3HIqDQg6Hwlz/7Czq79KedJQsWEuUtmn9S9Xkl1R7o9KVuwB
Y5WpJkLEnQJtQV5aflm8jLrZfiHH5+3UfJlxdDJQPtX1gJwZRQhKaKMeaGgTL0beJD0zN5AIqn0T
cMN4dUbuNCrAqyM2vSBJmJSJOFc7YgDlw+QXs6NTsfCc7rX/u0SlxECg7Ac1+zo5IIzUxW9pbBUE
DTaEmSnwf2Z523AIOWYCbqgdca8E5qp5AO5ZCjUoQIwcDZ3gKA8OWXsw3Nobf+ldNEJMDa4D7aYd
dy6ty4qMlWucWOV9UuFiq+vI1oENhxsrQOUtQnZDvY1JirTwMuHIDcWK8qCt6LuqTrkaJ2K8ib7Z
ByXUs7u5QW1DpVX4NywAz30EtNk37ygT5gvQpbobmcvO9jlPtl1dIXCQ3yrDJF5a3kjgHgz5NWC6
HUxVdA61vkhr2vz5T0xx6xp2RzSDSL64tb8zkK4HMItzYskHXOCpZcECijU/XP3iLLzxy6fTmtOk
EyTQflsr8zRfku7zTb1JNSW98Odrh3xqalAruumii/XR+9noSimQioGUJSolF3yX2hhipuIlQJ9J
z0wZ9QjQ2ImgKMBv+RNm6EztcH6F5wfRXa8SQhkMr/G+IMZTirxdaRr6kMaM+VmygVz+qK3bNG/o
WzNUgiX9tjy0VKwzbMbSxGzo53u65TylN7iR1gH7+OFtLjxTZEh88BVFMXk7acVym6UDZ4UAYKmk
q/uLQPjC1svnEuyj/0NLdCJWaLgEkVyBjLE/Ktu+6o1FVDffVDcLz9lkIgu72lyONqwsEN4CaOES
+vf3cw9vLA2FcGqKcu6BRDWRgnuFAsDzharysvDONG5r43R0lz67fR2Ht1pqqFJJ5FlbmgShhCJ5
YI/0Wp41Sfn/zkdXZYEEXGNawtDdQ/60AcE89qKNGreKxINjUg5XDNy8gE0ydsHgp8LsoLmf6Hr1
4HxPVY9XViRT6wubiDpkdNAvMBtaDCmLzwYM9rhtDWomJghj8opQ8bA7ki4rP9Mxjdmncrn975D9
wPQSvdVUvxIroitqoLQWUjAhI2TLsacN4+/nLiqYT05+2tuhvV9I+ec/TseTT1Hf1BBKeaetA1v0
NKC6NMwmvX8lHTa8uI2QrIWt3iJDrf+QPXkzbXkoM/fbS1tOqyvokyM7XKXnSLcvWva/23Ds5bG5
nEbyjxZBCXLY4cqYjsVFmQJ36uNyS6inRz66k56QKgF1GF5oYTOIdsH+l1tNPOUjQ2sLhrsXPjHm
nMu5+n087VZt2SMyROs9jdWtK1KSYUp2CfqEj/fe56uY/ySVn91WJMsK1oWBIwuNPXheE66IKF0F
uZbwLmZKnTqbXvISGL+AO0djJjE8DExWZ3rS2+yz+uUW3RQLUTrOYuYiu3HE1J7/DNBFhvmfSrBq
igURprvXkKqxd/q4tFUddgD8ImqFuem9NgazS26J9TIZ25KaLmcTm8NEcBmODXFhSMJdbldL28p4
Kk3okkkU1yNY9/1j83y1EbmyS6uVTWt3rwDAeERzzKSK+8bf7yn6WorXXFVoRRM7J9mZJcK8cqRS
Bk0P3e8Knl7PijciTxdZ8HyoT47vEAEm5UYTwMaKuIQBuKn+/PwHF1gsNrfIbIop5rfeIEg2dD+v
Xmck81NxEXd61cZRI1cL28n85JvBmNcz+YtzhDi8oHvBmx33Epiy97xC9Lp1Fm7pgmg8ReXG4kUy
527NSuS1GF1jPhP4MWV65xvSqBZxtnM5mpqodQaIW5RJzuIPEwmF2rJ07UqnkLTFemNQxk9VT4xU
BgtjNAylz9stczTPOf2hqGBlYuLNiH2Hcvtr7YibZ0upqYNFFJJSHvyXBNR9F5W+ur8YlTMcraWQ
uTQxBmORLMKvAtmRFuzKK1hFhz3sqqb15twb1vufS+gGmU5bDRxmcxys3HOBKMznxAuVJS+L0WIJ
KIg5A769M6f/lGAqvBEcYU91h78mBVzBvAevXdzU3GueaarKaF5ldP2zgDATF0JdbEQyMEVAgQW0
t6eRTCH0NjsJSmFFWImxz3dBPuALwge/nJXLXTlrwPwwxZ+6Xdy+IBMdjF8vuXld3oV8JfOpNlC+
77FoGxnH+kq+40FJ6j3k096aUozyA/x1fGa+WoyTKgR2WcovVCVqasuXzX5WEduQVaEEUbZHxnCZ
kdpmlkqAD8MzQ/YVuM65Pri3kieSxch7olfyuJY3f0ny1f1dUYtv8+xqF81fMpMhA434UbWGVRew
JW1nRSNKZsrynQ4r9k5LPr6k60/o6FrIgMAnaRZx1bRJCXgHtloiBnisMT7WiDsX88P82WVQpo4b
Avc5NZyGMlU+wz3vxM3hQZHHPSPsmo9LgzFXznQdcyE8YKE5ZJlOj32Xd2CLSSvmxd7HVeX1BgcM
uU/67LMRaquN9ETJhURqmR8kAtIBSDlCvXbBHB7MtQvUy4WCSorOk9ZAPRigAzewTbXAvq2cgl26
+rJnYXNc64EsfDCvaEbFj2yfdHfNIFKELQC4MGktBhb3mqTuGvJPoM7XNRp72cRWp6Z/Yp7jHKvn
bpimaz27uxr/jK+Am8S8+x2sQlKRHVsVlfuAog8NmP5rxscBR/+qOy0O3WhuERXZpUpm16vgm/g1
8tab60RIQeRWI1TxbXEncWbV1I8O/wV6L5C9qs9BbuTSyVS9eRkifU8HW7x6n396gfRElGu/SwML
aE8xoD2XwgQHr+BzcpLT18SCvtZSVzxASsCdD0oBoCB+QKTgqH69kwTkbRMtyHkDLbeWER56Bx5E
mF5Uq++SB/9yj/pkm/3XGiuHE9El0+WhkYa8k+5RKciaHwOpSO0rAc+a58t7BwGF7IqAaT7CViN6
tJfdLiWE/agR4JM5IlbwtSp6dawUuXem1GUKT7NUEJXGoxWsvxOBX30xQxVA2tBoYMvYie8n/uNW
19WQ2klJNHMwGlzmFvbs76X6nkzUGB+10C6wTvNRW4dSja5A0PVBjBCZaz0Yh5QaWW0S25GlAj4l
Uv2jFnKeb6De9slr2DSGvHg7l0tPoOoUpHhajRgW5f92x55WrtPz41GetTuSNgfJ7m6RZWkttDd4
sg3O9iib7Kqu6x2IvUh3dShFUJq/TBGryno6msXu0y3HIbhsXjFdePxhn2kEzvx4LBJpz1rW8GKb
xNsQXxAKBJBrLFT+tIwmKEBpqmjX4XO9w9WL1jxBzbvr/TZOMMboPlyNgSNPtvDIJWvZBUqMEXa0
xFP+EQRSrx7ex9gG3VXfVAMVBlGIiFiIrcBUgQtQd+zZYVVzkvZhNbIDTDTKQ6+pRZahhPT9rpc2
vdxQsX4QoKP0WK2NpmcGAN8vYdbodo95Msxjd4lcRVtKaHvkr+//I8LkcyD+b4rs67QoT/M43t7I
MjcjehWCWqBcg9M0gDHnuBeRkLzUA4kihbwtYhYgKO/kIBqarBsAz0AcyTnOgK/em/e4NgKdKeco
SCh7rPvuaMDmTYtLPQhWPQtvLRmis4/ie2NuB5PCWi2TWXI2z6z0ntsVuUDIyy3Tp7/i0UrmytNV
jWxkYZOHYIT1cw0eI2oiaCVZrQNvVl0R3bkfdEWOuhRK+5lIJiyFjvxRRJEe7drUEFqKDF35PSBP
vmgNJD7Np3IMA4lp3S3GnRn7p7nS/RDJNYGsAFfs56s5aIHSExCS2tiiccGHbg2r3s6Z1CNhP2Nf
U2g5ixAYhuChjICeajvOUZp8MGQU7DEjSpid6b491WHQwOXFKujXiCJq9tdu5RjvgYVXpqdtAw+Y
CuBqtk+zZLcsl9BhNWtBf8oZkmaZqLL268MJ3cHvmuGGfuxqngKNbqKXZ+mKxnR7qHKRBYDiFGPb
9vSaJd0md7vFnSk/krKWpkkaGmvi83z9NEFfR+jjUOyxbAbcvmo5FVyXQXrGjJYE0RaUeUu5fwOS
2TKfTwgK6YtzK2Spdr3DaKFU/Q32PcZq7F59zmP0PN9rmio3lafLKgrydsjRhZLsNsC/HPkpWu1F
96E6n2s3BVHC4S/MXh2midyWnIg+Gfk8NGdWCYrQsY9WUoEGmNd+PIB3TnOx0PbQcjl5wHyKOZ90
JsA1ZHuuCUB9u6SENOH7mDJUrdAbmA23UjHHccyJHg49D8SSi4ZY7aXByVKxkB6xwqTkVgaX24D6
rLmAJG5Z7pwIxHkM822vH8GYSyRXQNUT9/OPLDCbPtupgcPZVS9JespecOm1pyfYL2sNLINJMj+8
cYKRbPSU6TQXYcUusB7WqgIC2FfGw5XxDNcxgVEuYgibQD0fB50ui/1V0b6AEDETWXi2w5339fuU
Ndvn4Feo9kkmatnLZ6982nfEs9zCF9UlRcvtoVSQUQ52c83bbWP038JhHV/D9CJZ6zUdFmuyPHTp
ul5/fmgHNAoPzOLoDCP4SoLij4ACZBzJvj47YkE7e/AmLqqNHWEHklZcMydFryCTH7iOaRWm1aUl
FkBV0RL9TdqKF93okAIfbbhP6O+F2fW4gqOT+bgMvk8gvD/8+9il5+3pQ7/sKclQTTQ9a0Je/BzL
4GwOVRN21Gc53r05sYV0I0LjKcbWT0AayCistVlM5p4NPdRV0PR1YDAS7a+ctjyiOSLGrvul2kna
8APAeYvSA1E4RJzdTaumuhR9rOW4/6TjasRtjQ2aQamzLou4I2ycy1as7ioos/m6pwIM4jjSz1aT
9XF9bgPzFHFbrVwR0PVDSIBdXip9AUe6m7F3OMMotOJDz2i6cQnTNWtkrm8vzWyPO6CpRcUFtJr9
GwgTDPRkDkgn95Iuwd3Xu5j+qZW4Udiv4ElPp46yC+jfGmjTtTb5XyTsHUoo/YKKFz+7kMax0F9N
MAoyi5hrZ2fhxq2ciIbvDzzhIbbDV2110l59pm9qm5GQ00lJNmKFVKEgVy48j5BtQMqCV+yuOfPa
CbTbH+wBrzTxZOBUB9+ZG8z4rnN7EAt+W39rDSkp/sBYx0l6gvNGpH7g4H7mDjwBLrhEjrBYK+Wn
bDeYDzDG8ro2S/144gy6x9xrGtRCFOWartRkjdN91ZNeJGWPUadj426QYAv/i71+4u5t3IT2WQ8x
ZooG2oUOJyH4kUK440c3QdIIA8CjC61+ZYKMWAW75m+FJW6BtuPbgrVO2hbz9ipHxMHCpy9QTWmo
+JFgU/GTGDjX/Ye1PgiG5WfN5INLt3up8Q1SgW6uj866lAeYjihTbrksAomQC+qQADPq82gI/Bgi
v+DgDz2gsEYl5MJqOJd9q/vi06aWRaehmjXYJ/qGEXiH013gSwWbaYFQ4Iyfc2AdwTClQbbdiKO6
2FMFxE4xjt1qeiV9iBdaDtdoJWiFj8/1ZeHGXz6K/LkRAy+V6gpQmwvjR0+AK4AzXrN5Zj5yUadL
+mWzJqmprw3ZcTi3PiB+jC/bUjlZ2+p3C5uraedxN/3v6byOCok4gGFnUUgnHw0FwO7YH+qRnRcF
hYiQqjiNtUJMY8AXE7Qqzv5qBlHVyBXXjZ6W/bCKmjwqFWVP1T8EgCi5E/wnrTVV/DEsdrotzCP+
k9fxY6FHAZ4q/QptJtfnljd2VpzWXCoh6Z+SGkmYfkfi1VOEuwCTfOCk6qTKFejlu/pRiUTvIHuv
dkAFo7EoPvk4fyui3hlUL3uMrsVcOQz7ognq87pdmtc4cMki2f9C0IlNtWyBVFrGs2h53G1H4qBm
C5S6CHn0TVQ49OyXC/GGp645jj3Wa3QMo384g69CDJ1rERY+2TKHZfBgL2Euusa6fK/6tPgb++hI
8cNB7Dm85UPOxEjFhpI6+KF8xpGNl2bi7Ov8x00AYgfSGRlkT30FWgy0F/2pKIkSpKvHa1FAjB/2
MX9Vy0OPNjKRmvyaRPnnShCncBNU4JacIOIO0EhRFwDyBU1MbdSCQSvTxf+GGogwtrCZYvfrmr22
5sfxq4X5XXMNv7pOSCz3fChVwuDRk+RlsSIEd77t537R5Yf2zxe1Krzo7GeiroUertyUWdgs3tEs
sh+lyMY8lssR+enr+lzkv+PQ808HZOS00tPgzMhIY7mim90R9FRWUtDD9oaWEr8w9JK915VTz2ky
hEaNkcieJOCCEE9VF1xpkcxLzf4OsJ1CYG3dX5p2/zwbJWv8KHkZwNIJz+KqkucW2n8G7zIs0sHq
YyaUrXNw6CtREMhv5DjT4q1Zfz8iEIaYMVt5oYONfUbYtFwxNrvDXgwSKuRSqE/AVirJnTTRijHa
2tB77qLRxx6rtUNrvbEcGjQXRINeEdDMbD1YvaADd8Hbj2mlHIdutU5/tZwkDQCDEWyrGjw5wSgB
Am6M9UcSXjjo8G0dK+rrZTz5quUXroNNHLB+EQAfW7iIvFYW4IKkrD48qt4lVHAEvMUwzf7GTtLu
SjGkhLDYkP3QG2xDk8AdjZNJ//0bPhXcBaCxobelenJyzqszV9BOhIKJnFl/a7hHb9KxLCZaElfO
bJnf1+FF1WzV+oOPY6PAa8FLoQWrdeplK/ZBGQo5toPDL059z1GTiMCmruQ5+G2fD06Nye9Wz+La
6JunpAvdw/lwFeuYLHz26WFKY7fU3kyScmU6ZY8X3tT7WHnThQ8EP6a37NBKMP8r/hC5z/Dob5ov
S0/PrKlIszAEdxM/+3aGicmxNe/K2Hbt5IdxhTiiYPXAWbGnqKdQcBJfFQO3YEiGQKCyjBhquvSQ
ew1FpmNx43v4yh2YXu5mG64frCXg7tK+Ucbi7fKciI75vP8h0hAdUjhdaYQc0hRBLxrkHKumVqE+
PiBRgEwrm0NYeuvRrFxf8NzaAe0EWMQT+8byYHvWbsn7r4PQYIpDRF+CPdGD+Qg/SAKnjaH+jA7k
hBOLdxDd7W7HqEaPdH0YHYsT63bUyVXjlHD+CRb+7bghmpyhxgE/K52TCERiXqMAY0YPPO20eivJ
3m49YbNtUo0TM7gVk6RIn8UAZjTbeaWX7i5PN73wNhus8VnXfK30xD+XBP4BtmQ4ryhaggQmizvU
aAUxeFnvpoALsHUaGYTKzU7n2rg7w/BYmAFddXnVk+Zaia3/ArS+/FERsZRHkvSFfr6HITsr8GR/
Pf/27aFhVleVaD1H9zR4o2Yx+IOHHHbjBHUaWjWyLVoNS8L4lhSGk76/6Lf+bC/wV3z2JffLiyn2
nF6i25CfY6eTdMbmwg4h6aN542blCSEIkbh+Kg2LaFvV9oZx14t7OvS6g6m4YOlxHatU93petSR7
YWZCYH5zBSj6s1fTv7P9FKkeKI6kl6wg2y4CCpiHIrZBuqndafYmuoFLAjI8A3RZWrPKbT8vGOpy
LFvVb1ggaKrSyoD24Mi3tzH52Ma4V3YD3pKNsOuFmeayiP9DAxDft3xLboNtK1cqIvLfkFHAwWyw
kyyiSxWB/ETtApxGA32NcPmhiAnLIlqoa//VNsP2ahio9SkP2YQO/AU7MX92O14ZK8ZE+C0iqKVJ
ame4t9CkAJMSj7YASoMq1krlF7aUt+oOiCSc255OOSLpCJKpLuOxmYn8y2TEbyVKHBXJbi2P1vZa
E2OUJ3PB/lQgx46Bi8UBWA7hpXryyyOs4mQVVcU/P8aemKI3K3UcQT+RU35dwENI6hYjNxjOaHbc
E6jlUxeLx0P8grcm1uQWz7X8nEdBK88DZjzyO+s3dxSurHk+6GKIK1z0I17kVj30ezA/L2scdRgW
GH1I4dt3cUNoJs9/a3M9JGQRWLp02EDqvmBP+AVGmRk09BAgUqNGPQaN4hdKEiB3xaNdE2qFLKf3
aRxO3t/R9+TnGD8FUkKuZv+4h2cW8un8htUECXz+47R5J6TCL9kDDXDHS4tDHHcS1QT8kBeRyxZE
+XgvFwUXV4E/fwGMlcR+lVgkfAhIvafZgVJ/BBUpsDss8SpMTPt2GBE5LMioW68UK4pzAGAaDWBd
rL995VeGdIMtr68gvZ63tIY36+15hHNLFXIz1xdeQ/DQxFaO1fehq5QeohFb73rasSpsgvXH5Jzc
863SCSCGhkZmpcoc7qCE7M4b1DLq1RO4whTcEG+NHbR80JSYjiiJL8qawLQw5YhWEHE3tEu/26As
KB4xBWrXBHFvvwKAu4kkr1h6CKiAkQ1EHz6d/nV4sg0/jzU9H6AcMyzmYPI8B/wWHRBHOP/ASim2
82EakuxHpPch70STLTGdCH05pr+EyqyiAfn3nd9bqEwJh0sCPMNQZrDTnq5p7Mfly0zG5AqFgZ/6
pguySachH86XiOXLLJ7xlHYUob4y8W5rRJ9F1injCjGJZfuAZfRYFDaZMj8COnrb8T8a2cYbvFe1
uZZuwomWIWpxgSpYwO+gZ5I9gTXUU1jbQjBqs66J0p1K53Tj/Iu8QYi2JDUlOKUh04L84ttgTzqd
M7IrGVz6H14Lpux7PYiB3U9jhdBzUlSYp3R31/R9hX6lKr5r3/AAt/Vzvl7m3r8HM+LAMCWkzbDv
abXkffQnG8YqSKBWWiG2xQHfB2QPcEoJYfdb/KCR6tiSno28FpVYmSyDQ/AxFDKDDqIgNwga2ru9
fdJDG7inwda9rtvUznhXeZkv+T3jS6i1hNhmGFANdkOZVDNWMEzakdyQoMYnJbLXQPukOnwb3LwI
bGnTCUUiaqrlN+W9keDdR2LJdt38y62Qg64rcULplGTHfkNkenLvEG8+8ahIzpWuwLJcwAWpFVV2
2ixtFlhFBAwKE0p5oeoRV+O68PvXNbi1lKTU2xDv6a1kN113GyTNiFhlqpy6r6NIGxMesD8fu7MQ
BgyIr6UluEWa/X6avn/NQJvsXpFKSGABNITJ9qCwVOuMJoktb6l7vugxqyrx/mkhBzaCtIuVdq/H
VlEn5Wjd46izWoT4D2f/2+Akp8cVdCzZhlB5mqbPx7yvyjD56NWbzOZbzoewZZq5fEuXegcCJfmn
G6sFlg6WHamVSzV+7MXFqHH6tGQ/gjL6OTDUXunTxoqP0xOrIZxmPZpyFk2EBxEarAqwEpSawTNQ
z60OHwJlcaPJMNTz7ldRPqqSiHXc/ojeIteW/LdcSIJvxZ4yzaGWfG2xoul7U7bOYBTPWAdbA6Gk
gavBJ3TLGoql4cGVYFmtFFR8SV23lnrA9JTO19eHbKSQfPED9LdT936p8BJnRTWQyCRFxc+7Ra1n
+DNH804hBmMolREkAM0/i5CShlgFOdJ/WQvgOKR9rf8HXQF88DRoaY1TUA8IXBVekqLYH62cQmtQ
AOM7Znwc00Ri6/FYfONV1956lbe9MmJk+3Xf18SvFAM7TXkTD6ygqeyMrUaj4rixqFnOmsVWat/x
5M2CHjpK+C8Zs8V7+nCM2to5zm5YAZf/h8qi9kKRy9rdnXJ8z7WoOMJogFzg7LMvIFEonOeV5trr
3g0NQKHHhOJ0AZVjMEJy6+3951q9vPsfQ7Akgw9j9SA6DeWvhOzXYqxrtdEvPf2d6hIZuzxUzjGE
+h+cs8oS0JV8DERQ8K+DfqZwbhiPhMu74URFsjbWYS6xXUeT8yVPEwE/r0XM2AFVUnJGL/mRfZJ0
lyMn3/Nidr+/cJc9PT+8oq8bvlWeZlijQEKj+3MGQqUpl3TWaU9EnBiEqh/2Lu9Pa4wPUugNK5UK
qoBdkJekxRumua1Pf+VXzROx89WwKncMZe4s/K/f3cwDcA/CmhGErtL6NFdnW/83VrkP2HfwA5jM
HG+L03H91NxcUWPcdP3iXkFbHh5EZWtjvNr2sDQz2kPyV3YwWqCowfjhDdOYEqAjqQoRwas1t9WX
n8AzRoPy18c3r8+vMDrMyEkrYbqG+wMxGFAKHf1XYI9ISHB3qHAj5E17MBPMDn1J3zyTpo5sYr5C
yQ7FKZk2A5YdvkIjH8OlP9k3gQMrgQP8r2SttYZS8HZFS8N6tWyIjEfnOKIg5oua532qhG5m3SA1
T1io1IUHB+23O+K0JGkNF6PJvxh4ne/MhAvFJdJhSfvwInipqWIwI2sCEFZAbbPqLgq8e/0Y9OMx
Y4CRwc603r590pRU7wlfwK3wAfcGphFeWgsJS6Q1YnlerBCcpcAirfdc0w8HfuFUzbXciOxKmqqK
jYmFNctUzIF7erSqMX3VQC3W23SBJZZWRohAosDLk9FPqHnHQoj+VAUcWJtUooZYFBHFzjP+rEBX
C+Z5+f+65+3Q2ebFGe2mQMjogAyuDNvdtWYyN6ttDSyJsbqU7OC6R1nO3ATuPGbqAVj5VqFqMMKq
Km8uaGUXG2jbiMzzSMSmz+P1hSMibrG5Sw4ODH+zpsev3CC/tm0763Dsc1QcAbtPifhjufYwE8Cn
9TCcYry9+TosMbaooYSkydK3tNlnHILkOjWIMk36+JtOoZh45UNIMYbivGo2E05ly4vFqFy+iz1Y
KcxfESDkmPgiOdH81b5sZ+EhHBTYNrjGZ/PFMkhNOhxLLLlZFnY0j3yVTdouAILT/eQi+KXTA+0K
XDLHsJW24VZcI00dFpl8v4kRqbSy+K428MCDgVXhEO9Ur5aoR/6CJE00L/y8WrPHTP5X4+O7aUYt
Y/FgUaypprsI4jHpyPyMfAgfyeRzKZuW2Q5gOBRP82iVvzzFCEeJHCuCbuscuc9IM6A5R9eko+CM
+7uiGRHRxxp6TeZTJELzxBI+fUj3aLMdsCsZ6r182JkZDTKZR0IRmUU9cf0E9/06VWP1yikDcMKX
SVXRR82cyBZ3iYX/mRb3ljooeDoe0lw+S1ZS2Y+je+84C4nW+Upq4m0lLhxEAf8UZ/QmiKM5OH3G
jIRSiylO/ka3qPR2vGskozwcN6vrmAGy1xNfipUr9Zm7ERcA/0MjexAMn/oXsBH/FtjbzbcIJRw9
4J2gWT9yds7wEThb5aRZ0slxLfpSbjV3xRhHQ8t1gg4Ql1OYsE79bX9cVXFyJhDMuVhFfwBQ1H7q
RVpvTCCdYOTXicUrdeopvQ5g7KZRqiQjbUuyagowUth9VFa1kmEn86qNn1uZjmQQqUXWUQm/HG9L
4jR/rmKjF5o7wG9g+VHYiLHdqf0TehjGlkvsoAU67aLX7AYIo1FLg3bxhMgPBrXtIuNUkhmMNitV
GBbHaKjm7HdznSW4aJvAfIsQ7XkngmVl4heSdYjG+LFGfD9GtuIAp8dP1KxH2dGtgiE7k3nAYGzU
7AOUV7P7UfewMog2cKPYQKv8FcM2Qar7GHQcZ/CC4svwWDnQ/N26kqw7SP17OH8WEtHGmRjLDFL2
rnTKe1V0r25rC3i6zOJ7cyB4rFVKP1YOMyISGiLhacfND2BhUKWNoIQ6pSXTkAivUjgeAD4z4DtN
xePTlXmkD0ytpFWZyFlLQ2e5fQc1PvxxB5Efbx/RZhpx7B6ROSc/If3ENG2+cv7cvzIKymAzlV6L
0tlsf+r5dlyoiwci7u9QxOT0jpDkaQJ7OlVXP17JXtLYcsCDIqf7zOLvLsDZO3WWu8YKGhmWXlsB
m04x/DICajFXN0aiQnB5enJ/Ti0SPlBNzCiyiQNCTW0AiPdwPEBgzWcJzideOd85NCohwdF/bLUR
Nx8oxeErhtqn9H1VRFLoBj0hf/eO9556nl72mQq1wIC+55BmZ+6N1O9Tx1wxB52VI9wZjr7H+Wdd
mlEVl04Iz4wG9If6Y/zggzxRNZyfUVo+hZW9A7rikQnzUt8VmyIg6rbmGZQ3j1rCvy7nulJlLabt
czv07gdMWfq1HfLfitWON7rxgFjX41VCOPdEMaKAEGTnGufIP8/6yg+PvGNhXjT9Zbtq/4IM4m4z
pG6Z+VL327B0poI2FxybE8eCzkAeW656sdZo4uHQnhwRd9EfZnUNGWBkj9LF+0sNb9HO5u9NbNLX
HZr28BHrcRgykgjMdaKVllAW31dpu3JyQmOtBmxYR8F3G/e23DwYixSs9vwRRjAJTv/v71FAyb6j
80vGKhp+zl2MFNMIcAav9ZgwAUNq7Fa5Gm1LC6gk6o7t3oAhZtig2DbqxxaP30p3D0VvSI7+tagb
unOWEKNr2p3LWBkurfukNOjjUuYh2PPtyuPrd+viD/a9gxuGM1xwHn9bIEv8RCUCRHvGhyXBJwG2
qJTf8dD5sLqLiDFd0Iwo4aYQxObJIYltIQVNP3WAfaBFnqQFD8iINdSNbk4UxXBpfIfcaULI7Q7j
7B81XR8DJECtjoxMtZ72s5N1ABXJpIAynvQf9fViRyKd2BRKZg3yA64ud+KMksTjbc355/jMj04u
/56xYwIHcm6Htpm3kAt2JhO7xta+ZziSFMLxe7+hww3ojwdxXy37Bq3U9zjbx1v1AjXu1mVtW5QI
8IIH1aYpTIfFtR8AhjWVnFW5pV4LFzO1TOvEpFW3ntxzIwh8eh1riGFuRAlvn4U66KmOFEEJN4ia
WJJHKIzhFvSMDt4xisjf8OHkMVzvM3QW3SybXK5fDq6ov1x1FOltS7EJh9Ne8iIEIZRQmc7F4kjb
qKud8s1459WtWIbxluPBBGyJAicRPfZ1HMePvny4wyUZ+5eFMx/tMKjJdPUAtjmK+/9fZB/AMspd
MZL1LhLoGlTBM8TZLb4Fcsz1GDuqQ6iGERC7cPSaYap+htqXjzj7Imuxf9IZvljoGwbUvEcTc4Js
Ms+2YfGCHLnsPw0ikZ48gQ+Dv7ThxV5XK4f7O87EAhz0hMaGqQwvjclqVM9AJdaOQqn2vCv/vZax
01w+QT/aqLAuiAw6L/nM5j0cbep1Z6UuGAwvyuLYl0RBO59YXh+RcFoWoUYqXTstMkprCYyjj873
AykwNv44t4aFhA+VioSl1Rl2bPvF0omaX+awlY1rZpM7edm4l4/Q+hzoVD0WiQJpEEAhagvWgKfO
Ap5BqHGOMHI6HH7n8Agf2GYCNNmD1CEhP6todLDnAlB7r8bBqmCmdRD/NYQV39djRxEIoxHbKj+V
mkyJoI1wkfTlnqMugWNPsUdjRNo5xXgai6YFrSNQS07LHV6JV0tfrWZj7L47oEz282rDBKVS+XW+
78gL+5GV9dUgi29uRI+cDmdwLpGlwE2220wk8MgIyai74qJJbEGTbvcBuQsxvRSHsJU0mJ4o8xIG
8DMC0h5phLFFNwOI7CQPdNh671aKL8fKckBoGlOVnLZAHFOvI+z4+nsdi/fkzLRitb2+954sT0l0
DsBtkmfvo/om6U47Pywt6PnIBLBw4RKuSvyWBpBHMnHkow4m62rYr8PfYgsmQUWilFfrQ+BS++zd
Dn/XXBJXBlinNoDquQ4LO7jnYCfPl6Thc11GxNfcyYxquxTkeVSY5WXp+d6dVNmINTuTaE2uxgOK
5KPIivb3pbPBiymz7gN0QzjfbtOofu/TUFKQVpz/7XQD1BUfX8GxAXZtGeM7Eyn2Fb3jX/02zKai
sCkBAQMxW9UyGXCwk3wtF7PvX51r7B7cNsPUEHuBRmKj5njdrDivIHJuo9jZ6oJSZhxfpzO/3lRh
09i9qtSqKFUhkDdJZXPRDBhKHm22OUgHnSl4BuzSLY/hB8x/YIIHCyANpsVUC+xP4ehU/aYOSAth
XwxFflrl20jZJW69t2qA0JjcoHHJWdqJBQqODnygzrEXsOi0zr/KR3ZtuM5EasHF00Of59TE1hNa
W3a26rd7a0bvlaItNYa02qw/2eb8qvF0mMgjVnLCwOQrtOtTxUrlnqgx3OGuroT5N5pacdUHeLlz
tfySLrS3TKf6IyPuhG+905hf4jHqpWp+aB+oRsSiE5gUwL2omYt7qfgmQgqqXN+pVD/YcYBEVi0Y
IYxbSZWXMR8Rga0XAYtT3RkPab8pFzOFFTyuB7kghBJQ5XlilQl9rpMJiodHsyZP1NjHEaje75dH
43u+lLwVzLOyjBdfRPc50QVE4eqCsuPYREduS1LSk4XfoQNJpJdMQO/dPBLRaS3fRihxRHVKQk+4
kwtdZESr4RyZhlhie1/TNFoVh3B24ZY5jLN+Zr5AoM1eof2LgmTJjE+kG4sVP+1WOoh/w9hVKYkk
60oxHjoSbvu9SDYQXSzR3LR6Jb5WbfP3H7gpTP0QzP5LiYvrOQCjxnLXVLcKUbGYMampAnk16OND
45R6pAAB0ukWlBn1T/82QhOGApaODV9AEeIoXUQidhtabs6N3xngpqobNzve0ukc2Bab9ZBg5iiG
H0cIaYfLI57DhldXK/6+co4ScjqU7T0ov4RSP7GrkMijyQdf6y4Rr9f21MEiR5weJY7bBqprTtZz
pHI2JWEeYCM1kni2pgDpqY6OtRxyIN+ZSTu/ZDKetNVLP4X2lqL085qrArkxyIgkaCLDYBMbHiDD
VGmTb4ThUTXzFB7UvDEy+nFZgYAzmgbnnegELhkuZ5vH+6VJTJ3zZVQnZ3Fdx9r0+hIJNcwmEJ9+
0XernXjYHuxRArXLk/9vJUCoRlKQq5vNtmQzrHSbo6dAhGULs0ii2qyyyyQNY74lRYDN0ZkvIvuB
cBRGXhEG+tu8TQMGU+ZxkI7736R/wNTuadEhEsfdKRP3UBiMqNT9x7JEk7skhKgbbOyhASqfeAUQ
pazN1R/Mgn2EKp1gkzhpwGzjbABt8urHypdU6Tl+xQGHIScFOM3ev+oF+WHqphh18NmaUxG1sKeH
PGsw7wE8FvkLuUYJiHsKJpHiXcPmPkaKmYI6iWEiYXd7CWoTBAU91zj980F3jVrYp+6e+pvKZGVS
/67rUbh8vbJen9iHLCPxcHDW3dI4D5O5RUKK8OxWCJPZUZVB9jL8ChjRYUTi2sm0MWdllg2XV99Z
ErPh8oyDJ28R7ZBoOUcowLALogyvDZXkx1wGgsNTCG4vF+N9NxJgIPN7zz9yjviaclY/uXzGI8QN
/YopE4hXSl7jO2GiPhlt9jf9Sm7CN58U7deczLlzTnSLIkA7oW7RWoLD75v2QBzwZqkAlHzKuKQW
i+kkPqNhPoJdUJ3UVQ1EvzeUPoSd0f/KTF8OXnA1V6zZLE1xBFCwW03VE+9shJXCUv7pT0wVkkrG
gi45vNzgv6od7Px5JMNXwqCMeBFWkYUYcmpK8HeIvZyv4UNmE2+POA9CGQGiUVwV2kXFpkOwqQ7y
iDh2qpje8zOkideHm9mcC2SPlD5Ub+KUsyhFhCneBjKl0LdX3GtUb9zkUriIHEQ1DR8uSfak6fMk
kR0vHmClnSYE3piLscjia5d4GyjdOfExnBzG+P4oG2igPf7tsqrCa1KsSFJ+Y75gYemTVBZkb8/4
U8IBBQJsmK51kZD0R+W6Btk+wQSHv9gRWJkbOa4dkwc+9On002MiJMgGqvognc+wtze2SzCtWgi9
SoMKAFUNyzXsc6Ipi6cU5csZdkPXv9K+yUgjy53jwhG4M+20ef5E9YEZBbfh4zIs6V4iiWRpdFpu
0eWjkrA807JhzFGUPtOl+FkKzT94EesxMThmoLRChqdz1o9+enMCW3htwCQK7aq8lW3FyI9F6u4O
kbmezrWP2SBe1H5ZXaL0EIW0jNz+acN8wKNfDwvA/nGtU2uVRAKW3Ep4MwBXU1dThr+hXWPSKx18
cwGMpOHyVePyaYLPOcomVNaw8ojz8AQahuu4FORfsxvuiPMDNq9RX+JamNaFIO+M/22gWAQRfl5s
KYuTg1Dv4NY69aB3o/6ZyI739+Cdd/2EXrd55zX9wxadgrR8nsWtvADJ7y5sOK7UtJjNnZbVYtG+
+VfuJoh1yhuhwK4iqSUl6EnO2l4Bw/TrWlzhH6AXFF+AU5N+5ZOurXpAUnynJE2pRKCflr1sOHB6
1fSQWuv5hW71+n/w9u5O9vVG1psAn/N48JZ5MnENnfHzjXfQ7HoKIb2iJvkpbdwqize/n6PWNt7H
HWrds6bjSORmXrLODZeRjSSUprMcReQeDVUlVVRCKmL+JFN2qEWrEVl4fhDnAipgqvjHRgfCidBV
u2NlaSrQWDv2KdhxQInust49f5sW3eJtzdtKLe5LlzGi+S5A1AnXldPXczlTZL+6N7FlJhuIWsTO
i0Um7FDD0gYfqrAA/KNRAWaetlhGkIFZTY9n2V8Co/jU3H7LLP4EacjA5fLrP3QYBqKXW1KyTCwG
/wwkg9Uuz3DI0wS82NTi7s7YIKL9efO1fMvPCKolBa3ln3llvrFOatoMupBaZZV5tTJt6yx0vHV7
CYUL5RLsI/MTcYivLUiHX690JiDg+PYVkjLDTSLxQYsf7kwBX58LXE6t/ToW3ECj6ajWkdXzYYKR
Xlqx8yzEPJYXf3vHKB/YT7DB50Qd/eBxwPDmSk5IAa8pq9B4PoqAAi/t7ZTIP/6RePlrAMa76hNG
wQOGD9mvn80jzfw178/NoxwojxPMydHp5MNsNnYfgrqoBKyh1l+DP+Dj8BYCTNKimmHkvRDWZ6p3
SKSCKJKnD6jzW8Lu0aWHWN5Pc6B8N4nBBUzNAhdNH7m8lEmjl4MsgX6xjjeMAAA1GnlwuajhRnn1
9IeEEJJPePU8LGCstUQ5AvVAm9ZGWKOHMTE2X2k0YWaYskTZbNAjqGJD+fy66yekTqhi5stsYC3r
HnmoWNL76jeTF+Bd4n6+5olJhh7pACzn5B041HfXuRo2HoUrGmrzw+w3q+frKCvNWa3U4wI6Weww
Go3py9U/QPehwFloxu0bi4zI/NdeyJItt59aLWNfIqoKgcuMrV26nyHknvMVRXMT/w6YEklDPnJy
G1k9sb2NggEFCxGv7g3UvZK3Ffs5rPiwC9cRdzIDr75P6WB6m6swC/fr0m5TrkT1sgbKpPtDGQy+
Q1RjJJ2ePT6FyiUwmRSL5+O0vvGpiwRN7qs2irRzt5NQka6Jgy2g7o3BbCmu4KrZYA==
`pragma protect end_protected
