`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13488)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCWkq9Q7sGKUfekyOUZQK4PRcosgQmmcCzsxuTnFB3d7s6toQeIIuciug
Q0f+emK30TdB91wsQZSjuTAIoNWYKRzulmWs/bNsWh72Usw34oZuM18r/NXqk/zyOpOYqDbkKl+d
JK7fcaF2pPPBhs4212VhL/lYQPvWX4HAzOgKKEY4qsegKi48TTT5/R1zKGo1TeJoACqoF0skc4P+
9K20Gb/OVuwgIO6sTywV+kWNqNvEc9InNKTpa507rhJGL5ziqhsTxM/bfvx45KcW87r9OpW1DA4s
XQiG8evw0YSTiqM9ZzJD6VWIIwiB8POps7EnV4lstYyR4ZA+LOcZtCv0YGSfzdWRxDsS071Hd++X
n5mudaz90pfkyJBx76aNoo4m/CUhl51o2TdMxn841uuHdxcOol+OaYAK6E21V5U631CedkRr4vkL
gzVeYehMsVxTb+656aTi2EhRZlGlWCkwzLx7mxbVveATjenBPc39++93L1IybQYB7qNmKAtNyV48
xZ0mda9NkLKw1lQIsrHk9iYJCSIu5SWvQy2R4gsqMCvQfLMBnrfwfOK4FyZk/9I1/G5e43ToycQ9
BtzEnpE3yk08pKV/pUZsFreGUOS26jJHOg0yAxkV1zQ5PBUgisaiyd01EfrZdt8IkQCGkrac1RvH
4LJbkEgIC2DMWmK8P9mJNyFStDqDNIXAL9jcBdb1ONur0ZHvamq1Lecm+x5XWO9H7vSovtg3tGB/
w4ohjQw5fePzboR9AndgXrzakuyGDIrUmP3EEIgNWC4JT3eJfHy2OkFJs5oEoMqAZRMg5yxKQjEd
40XZiH6bXojjwG/5Qx+hIJjA60BJE8ry5NtBjP9wzoedAf47tAOrhT44df0L03TTdzPECJtRGNnD
sm48RZgKRRy+t3nyMiIXvy/ySKSip8g1kQSZSlVvOb8pfTd4N44fnxClUpLXqoZZPVnMPY0HeBp8
U9LLEIMXvdl8C1/ZDl5+jzGY6ptUC/XMJygeHEWu9xOflKqdx0UD3uSWXsSiIDQLydIhe2Kn7KBw
cX3mizVssgXK8qkTWxVe12CH18A96BwKV8QLiJSgVU/usDoQ2YOKPdqrqaU574dYqBJr2wJUze9L
CRvZ4oQxbfJ56lH2JPAUEsbzJ57MTNno1vlAOjJwsRzBUHFTIE6zTcfsNEBA26ypbARj1yRbjXZn
+YLcHd55ysUuibQHY+lXHjvg+rzbF8kH5bB1ubEmze78/Q6yt+kIWFBwu4Pxa6JDSFPLWLCDuyiw
4BejgpwUIIRbfaVmFcd+5PwRmTIXchFUo/T2e+KCqnKBNAHIxzgX00oZK0Ujg2R0iTkKrU0Awk9U
t4Prnu9WqX0qJ3WPFzYT8soSyzDVU/SZrq3t8T4/dsEGUb8uq35KBfbC2SZMk/g/3jUB4GONPmdx
ZXk5Riaq3F/nnuQY91Hwo+NMtNWRJbBZto8zcf3e7HC9Hzzk7JqIH7FkwIXczp1ra2PL7h1YHSIC
kxQh1+cYHAKP5F4gASz1KfNuBAnd83Qii8swkxFUh2qUOM6rMQ5qjswWXKHS0+MuPCaXnqiwgpV/
IS2bMC+Ztv1rfwljbU5zICWc7NsPTg6xD7OtJ0WYeZN8IK8jC804vXXJP9YaOuFfueZT/033bKYs
YUmcsPszu5c53ZCkT0cDssPJdfxNgV2j0GD3mb5PChiv5oMkpDRlMPDbPGbPIinpl4QODAREjeeD
GlnWuaGzmz+5HwhV+0imwrh3EF7PsHO43gFFWiiE0ho3Nzd//SKUfmkoLKsuqPhhxR9+I/vvIhTG
GuhyfLShTL4Bu5rQwqpPiS8LvQOyIXFlqA7/TJFqBmRaOISSxNBSHnQDdPw+VUEzCOGBWxP9HVNE
2XLL2X95rKFs0oWanRXR/ucZpBGulwtbufjr4SWQX/qy2NMLBp2PLTxw7bOyRLOgwAK0mA6bxlYs
xoNYXgDa+VaMf9qq0uSmDC4gGl42jr9Z+hq1zZHFV4Yi0vdnGpkoNQ56h2vDr9JhpJnWpYfyORQx
YNZIIN1/mTw3zw7NWyfFdUBUIoMifop9QEwFdwrzu9gsMPQM9I89ARq6JuUlbMsHJXrmaxQ0EsfA
7OOtQmyXVn/+/wMfU9NdWIIsY5SJmhaeZXSUvh9/OnbL8hUr/kuXgkAdp9eTPglyPqT6EyuN6Qqa
nZfVuOqr6C1E5pVf1+bipLSFevCg0EI4XKBxLWqZ4SkczSQ1dm+t4EgcV6a3Zjn4xbTNzaSUJ+zW
nMQE+nuvLe1F6ER5LWHglJroGOO/2uckQkve+mH7bcknpnMDPusCU9rKd+icQjsZKpnjYGqtARZc
5pqphExYvmLmHN3TYWiMyGZ0ISsZ9dhKXp88Bunl6fsJog+qNDSmPejzAxVRbkLUs4JtPQTnoSHn
k5UpuNvr790W6aLO1jZZBQ84VlXjUZLk+VQ6gXgbRA0NemRaXDlLk5+is5Y5dr0RzioH9RTs88OK
s5hL3VPId1/vfWOx7/iHtegSGMt6VGKlRas7g/OYUP8u8eGdfz4M9ie8nCQRMB+Z0cXz/vZlhMwO
cVU+9Tf1cke4IhSvUCzImzgOfihk4gpgrMjb8fHpR9x+0cRg5wvA82J6+WcjiezwLK6AG11Y80t7
x6LLpBw0o0TrVr88G3B0XrOXD3HbrNxzjDnYGy6/UncvaRAwjc5A2k/ln3Rjz0qcAAoYoAgP/dd3
fJSUWhz1ttesCfaAvYsH77qZzeGWQYrQI+eAlvtR0OrR6q1IoDM7L7WqaPDNWKT+FnAXZB0SPsct
FqmRWBoHyF+yWjXih0Diz2MLYhvcOU9fQsftIJvMzlZ+Y0vO1LBblmUQQGCRVj4An6RouP4Iq03H
cTry8EXr/qer3SRDS1vht3/paNEyt9dW/yecCpeCOSGlp7kJVgQFZl/4biEsy6imyoF6WcX+XTTW
4wUMBYjUtvg3eAz0Ov+zU8y1UDQX7YoMr/wRZEMPja9edo9QmNoaj2zshW+n6eqdEBEWSLM2tP4S
a3lQ1Rtxi9Iw6LH5XMMMFPKYuqEiRUVoR3Tq3ITR33MdSMiosaMdF2u/uwVtWAN8WgcLQfhw9qKG
7jPnJAP5D24ve2Ygv6vDDQ5enxlGM5BFtwbtPOR/hYXF/9DGoKyujaRN9EUgCH2neBDoD3USsKF1
bZuieX39K4foEyATLUhNFTe3dMoDrW7fdTqINqp5a6aXgzzh9vp6weidAr4XG/NNSnqfyqSDhAE1
vAsVZPHDJzDCgxNOlSBlb/69zc+ntutmymOH5FBUys0zMyM0xxvaGUl+V6PHicaiQIMKXpFD3VVr
Q2EJNqejFXdjJAwkIhsSuJXGlzeaGS86i0TM46UZLa3qjeF+EjXTHV0g7M1rhZoWFY/saxH0yile
r9F5uxHbagmFMqLDj2hK7KiOXkvKsxqC63nbjhw/mEWizhvs4saPh/9TuQr4OSluwAycQsydIvxa
t9voDj1RYCGIAIbH5rCfyFUb5zw4rcJIU3/zmMk1PIp1XllwmQhQ1DXLLEyw+qna1F18CntApp26
FMjaEQtDBOaBsdEY7eXUCtgLEpSPdzlRhql7tdhpqDSsB5gF2mWb53h/fMQ4iHYxHCWgv6HC32Yn
1SMN4WmdRoFfpE/bfgKhUulIJdojwKQozoYnqQpFKyS2a60goM8PBk7Yip1FyOgGT0jCFyENX0z3
huF8zXx3CJMkG8KnaMJdI/ZESv9x0hrmkCf9K9ylN2D2X8oULuPUhShZRDWYZ8gTprhgd8CjI0Ir
M2fT3ubzw2m408aODtI7DeaLjBu79shXVu6GZnFEzOmKMR484ndyUOmlhav822YFiE/Sa6UYrom1
3wuuvyI/FTUDmJj/aWjxCZ8uHWeD+fDYYpz25VlZn+EIA2wPHGbeO9IleIr4Dcc+8KRrCQuk9wLu
aOUsWmVYykUEXLBrUftwqrRAIuLqd0cTWJhwhNf+dD9lOp1+jVprbVWvUcV8m3So8t1A9bbI7wy6
i0TCUYFS06+gnXRkcr1NG0TuJ81F+pdvF+qIRwJn9E69V7b4rwlqJBVQ6JZSZidom7j+JlCqidHA
wQJ0ZmfZREWIc/MLQKHHHS5io8wN6Ct8GI7keufOwEr8qpY9Zh0gh/V+J47x6PVquxJ6tuYwiwtL
e99JqrirAW8YmD9zGfOiSioGvht9BiA/BMddVnlJ5ptVXeVTLVcE7RH9f0FuCO7rVmE9VGuzvalb
lkMIuUR5e6aifosBvaXkuAo7xxpPZ20cDbAz358DY/6+rxoW09cQ52yMvMpz4J3jiwH13tQbb+rh
fGj0upte3k6tq32zEGwHO8wTgrSqrwUm7BPY0r5n4zJ1itSvVHNJqHukXP4ytQbsWA+cDvOlNv0g
5IQGZjnBhGbSmvpgYrfoX61bFQzlqNyPJxx/7v47+uEdPfnN3R/LTXgnnOgjfRZqONY1gR2dqgPm
mwwB39Trvb8W7C7R0ByBUS/YkghXexevm4j0oFWa+Ot9TpxK5APYSvLsXSDoMoOtOy+3E5mhYyL9
E6tCgTL8H/qaBugDhMJKyd3ZHAITnrbWhI7/GvBJe214tDlBIogXWckTWEHNRyFIIGpe9JHsZZwA
ZzgmeTGDH7sxdqnFLSxC8V56vFcuZvLu1pGq3Wlet3lJsdc0vR+HCPD8KMZxFoOoIVQlJU3CUxJi
PswXqSVnTBPfxnGpTlISQWefjdXpc4QSy88DQuIPiHiutQz98Ep6RHcfUENuneI+HHv0i7bgSx6Y
GcFsJyY18xN3a2lBQrmkT+RRv2KrsD1TiP2yuQs75XR0uAt5VkjraIthw/QKGF1qragY/Wsn6yc8
mfze8oJidci+iNdHC0oOtlP+X9f7MhGA69sDVON4svJyUIy9GlL9jcSrR71b6amff+TWY6ipIVE/
GcWZqDGcFojNPo5Z5ZVARiP5q5D2P8n029OqnAW6SXBVdEGE+KxIw/vy+p1SvR72EWmtwUO2pud1
JNxRNb6UxWAdm6vfsvs/McqmJR0CCa/lVh5MFW2gPHCfvIadU5gzz+M1K5+5ogqIiPwecuYAa0Pf
IwTv7Z5lYVB3GhShNK07EuGDgVX8/OhXF4f6q9ZAj4dGPIl83vcFWbpwXae+DCikKFIFegp+fm6I
rZayYM1lSAX2My8rg9vmCHoQqbBMVt76ur15SMSLjp1gTx//2ZAD1mlDHxyOjODS8N9TF8MhcwY5
XWFSsHf6Rn1yBFcqZ84c2znHBT5C1MXHtvq5FA/MZzmjWzDMIo4MruRLA0qpy2bQLnmbU9qknwIu
D1FUh39ZERRsTfS5kyPCxer1K9ho1cAilHUi5b7BnX+bammUcY/LvXuwu3vyzvbICds+3loRnD5F
pwH0+CBdzhzbvmDFxYtN2RIUo3uOjfWXZfpcTLwb7BKivpo1hiJ3CWUtO/1iTZLEqWgGkwG5nRFG
8S0RzMRm4zCWtrZKFMjnwV7J92h8uDUwwCuLm7P2Rhzil6e87NjzCi7tM2KaoPoWGzWip4zKrMNA
PsXAOZYLr/DYDtL45MmkNkIjWaZdBbOoQdw+/ZIfwgiKYWUEUMlrhmpmbKk1ao1lgLuKcyE1/FC9
KiNzOZUxMN3T1raY7nrngPa3X66wTB0Bbrbpb7SrFjgcPKA4uK3+3YHWkEufBVz1KtGXn3ZdejYt
RSRG0HDa1oyteNvtgTk/3+biokFtd1VDhzd87EA/RMCuc/tD5pVbQgmLxfAl+dNItE/7ah4l+x59
1OLY9aOzEnPt5MUOxdU/Mt+bFiDpBdzAJnZp5wKsOJVZKT5YO25iUpOAzQXgV2On9a57HcSPvL5L
5Bd7SGGozS5n2M5RW9USWsuNP0GUvYw/FcKme4zf4XzfndLDJBzeM4uJchz7+2e7/j5fXG3rCRDG
KCZIvaWZntnSek8RhXHAJbCjoMgxzn8QYhyhfrLMjaQAFGEwZbDNz2afoIPHcHi/b53emdMNRc2c
eKOPs5CmyammyaOkaOuAyrmA6SZoI+WXmPJgYXWwTY+z0GVuHkp/BQDFQTFaJcMWI7zjRUK7xOzW
Z+S5yZVYGS59b3Z2L3H5u8sHy+GqmPL+jIGqnwiYWPuYkEUKdLLxcXZwKRQynBN6aRLlzEfbEvkk
x3/lwGcVOWuxoNTc1uXAMF9IJQJSV+WtVq159f8W3fmBbAD64T1jK0Zx89E35DdWldKWxvdPaxi+
R0w12cWOXT/j5gGjXG/xJGjDtRjYVuG+pzzma2ow6DXCknbhSNMgbUnkNC8vxEZB+6DcDLLDc46m
1mer872l0ujMjD/ajQDAsnpHN0bK1OiLpw4MLQyEXSq4lbbL0jNNwb7MjY5r8Rrztj66b16o6Mhc
x0THONpUzCV9oeSYOGFE5P+LRl0vMD50yQAeeOEmd3gs3uHO00TO54i0B80di5RtS77t4lOkBe80
+2Z1JaIFclXVZhl/iKpDnkWqZ8DOuqicaqpTA8ypMLA7uwqmI8fqKFkGxCEa3G9aqI+dSMCRANqR
HWK17xmWgndpYh83qQvDHT2i3BMvL5wC2YNQ3L0NX4ol2rI3QHks7LMMWog5df4Syb+b3/lwmYCL
95OOrsHWsv+VhI0SI7hGye3wesLK9j4tvwntlQinguopd7Z3sy4NlTZTubl+j0muZfyhIAzup6A7
luv2etSzzdKYXgpTXdqaIhrN3t+2LPxw1t09lta7jsr2V2MW9Rod1gOOUWdWXPi/KdzyBxOx+HYJ
EN/uyC1VERQ/cq9FNI+Jcqr5efjTADB9St4qS7Lh5AiDOEYZp1zTTydvdFOfSZ+/nzbW6c3CBejA
TO5y+lHWTXAYQ2k1eDWVnnw1f0OcjLTu45tnrvu0Y+W9G0PwT9bfnL8t01ZDeoiLpVQMpPPZZoOi
8LfxAA6O/GBtYY9nshY9DtTYh8xIVvW/98vyWOxrr6owDc9TJgp6XwIqgGdUj9yecCJIlVmHkCE3
BSzq930/vz4h1nekbQEKK2ofWtl4Q1rom3cnXjQZ84zLVq8Ir5+15X80V5AN4MpmyumpNWRCaQL+
a1LRd4AUhg3YkbpPbSN4iapNGeGW5+tCw/tpqLW+OKZmpDWmcvHiOtSGedNHl4zgX8MZJu3DkaYV
GVRazDgzcoXZV6TcqaVthGozgmRNs1abJ+ELb3Vn08ATTLQqMbZsn6z7Un1RgQilGPvCV3BgWSTy
8Ct/AKJtZxOC+aB6wZ2AHyVw8Xrf68VNoHAq0RYKeDiInpABwRon0aCHP8fsOzhEy+Efbu1uY8Ld
9ykqRL9u9UNyn/q45yKji+F1zcOEKca3VZAlXa8dAPKWVAaagHT5VMwlYOW+TyFJ+s4rwjwhcjE+
rGKm34pbAA8XwEDGrEYxUgLN3Krx72rLGXRLuIseKKDVzs18bohGMz5JXrK21raeABAVoWuUTCE4
MeNtd5Kc0Ki7bCe1qVCr6QSanHH24OlxC1s9KKYH+KHu5AhG09lbt35n4K3cjwds7apna5penKIm
fm78mpIv3qjdAr5k8E/L29iW494q3iq/uQYfI+6mLG1jmRabPuYog/tS5ULGWpQsRvM6nsk+i3jy
0qh4pZch3PcauDSSMRQxjM1rBKkQXgw37MnoF/3cyp3zH+DQ/ZHmeAK+BXaG0IFjf1TwWhwdKypl
QqwQaDYhSdukBNRX+MFGpLXOs4C5WLkU9LGsDb0rwZcoP9ohG468rDjuk3kSHdzd7QWRG6s6LNnf
hlF1DiV/U/GWjzojBYAoQTkP3HgdtI/59WHUAT/eHjaJrANi/KLXegNWUBIVs705T/SAl9L8W5eu
+F/15NIQw0lPIiO86U7U5pAEXxck/hqLiZdRZlHM0AV2GVVFc/OyZrivgCAAWc6pVydBuHHpIHBn
krFxS/ZUb6j/pliHFtwXKi4vYE8p8LVIlz/v9BFTwSb2dWO0hIvOk5wqlQr7YMu7kj3DfQWW/GIL
iq4VqSd/i3EZZbdKqn+WROeyVVBGz5b8Y9JScl9jWnF/SvZZ6mAQ6X/Eu6vIVQuYsWF71KhMqvPc
Em99PA+N81z8Sq3o6M/KE9esya1aDM3zMpqR2DRQa971RVsjsebFbKTzuDjwiXReAkvwRW4Wl9Ku
9BRNMY51BQMcNwqxB42FVy5sRjHUyvMW0DUEhHl8DFPVZqswnLWF/lLXIIWx++6VmQsoyDQC0CG9
du3GFAZBC7jTEA2Duv/JnPLqqOscDQ6yQN9gSzMdlTvozqx45LwwR3F26hatN8il/HHj+gaTyTYF
g9d+cbzNp3zaYvSpFjruBmEPH9csHDaUL/4dzxzmDYSoTdzBezyAuGzLF2SYYL70i9amqIwmj9P5
RbGxY/a4+0eQgrYzdNum9ks0rzp7jw6d7PCZhyQuGZfx4QPc3xob78kDcTl7RMZftEC11joN1n7C
5/4BY6ROi/kY6GFzLnxTNBSoI4yc22CppwrcwV2c+m86zd5jVH3uHN8mGp1t3uvSEOv/oQYgA2Ck
epKlST+vo02hNSLbAoZK9Il4mtUGpZBwKToaRjsAKQ9L3aZ2xvRqxsAyay9cwiBkbFhMRftKHSXt
mWOCQ34dVWuqRu4GQsxo653g2RLtY1ExNPE/SVPpaIN2cGgedxnsBTIn0nRZ9UpZXRndXTXxUOwU
Xu+N29/s+MIrYmLYUNeJFK6STjcOmQYTtqWOTiESLnSofWcSDUSc78mg5UCdp98w6Tcsag1jGmTT
U6QApjpiSQyl6RicNrf8Of+B/jk4a3CQWelWsWKLJrTbjfpaMrDbTJw/ndqS9aZrz3fyOvVboERM
AcHHs4mz0GZK8J1/Mdc2KBQlVyj8bjvku+xWNMVkDtJF+Pfhr9WL8C6fKq/2YTOuAcfX6tfuUlgF
gOLNOraT7srfirxQmPZhQaAiJrQL2T2+L9EcaEqPsvmag3DbU6OJcg8hUxEcZ6w/xWRvOWWn732o
c5d1mhJSycwJadvMNgcEVNmHGYUVOsBiC4UvvKhnkA99F9Fy8Y4bTT5oyN72kS+UjwDDup5vvEAC
HfhMO6RfcyNwphjIpbVxBwfZYD+5qHlzdqm1jICrC2xPMz2meIg5hHZr67ra/LHHNcijeM2uBu9P
HL4MXgfOv3MZn6SD4SSByCUVN220hD4283p0qhPaJwu3A19FrjC3ikUFYwCUgSKMuZYHy4cAyIrM
XRSvH2kUhiKdmNvYZuKdkt8RnYN/nrElIaAu5l4Wz8mjdrmdbrQGlG6yAyEy+Hpv3vMImMcstuKj
Qcix8ORTOKgU1erJBNRjpV3aPGQT7pOASjjB4HyO4BySBeJFR6ADWJR1ai3Of0PKy/JZrm5/Cd0H
m4uE4cd4IF8l/ZIYr1+aZTCUAbaQC86tfFPaIeQ2fzDwYQGJiq9SzNQn3/AhEF+0Np11375QQI+b
yP3SoxmGJt/+xj6fT56sJk+j48svQ+a45/s2MQ7a1Rhy7MJP6KOJpXHHVSnSEbkGEHyCmF3cVjA1
k1oAsqvYmTGNGoOIC6Q0sQEqbScec+Ct2J87+T4Ewal82jnXZkfrHUdDsMTRi2+4lPjUrrJyRZRP
zLYzbgVBQbvbYMViQTPWN8xCDdcQ7H9n/Gu1aah7iSe2kt0wo1Vu5WKWhlb6i6vkOs2EmZWtHxY5
NZB/PCxhwDdoihdP+lRufhFGUryULN89JSasjwkaOfoXHndDGZ4jWPRsTtmINQhMLvO3WIB6npjV
phqcJ/FVRuEn32JgktQ9Ifa4hX4jTbovLaYrsjReIUu+3nzk4XJC5M5P4vz3WywVB9ADrsYmNaZ3
3p3Gfc6/VqRYaTdFsAm1oUP7pQl7ltLjpI68UbbOUDhmvJjSFk584D/N1s+s3gcvAS8xr/3rjlrG
B47eCHTY8y50X4abRfUr0/jhjDpZZXTQBvSmOzi+uJe5eNjwxGtJRnBxSNkusAf5u9PBePgc92bs
u57/plurszJRo/Go2ucmGfbJLgHqhSo9JbczR05ZGJaUCOr4KDvvykpDIDjY1GOBL7R+a0E9StMB
Q7u12J/39LiyvpRUySuNWuYdUohRV2ETenomGrf5mPJQAMbJylOLYLnjSkeOiXOb/JzIWeVVvVxb
HoH7qJI22UA/UT64qUi7yVd5nrCmQko832OxjEjibhR8oZDa6d+X+aM88Pp8s+drIQPdWDdOA/x5
f0XgT/b50DuwQG12ANS21kxh5oDJF41RCSc/3g/3EaGSlsXVMSrN6jP5mRB9LTOKXpUMV4jwtGcN
jlxX/Bn8DW8tUD9vSEBI+AGo4ZuSvjnBlu6LPRTBqPYOGKFH8ew4KoQEVdMuMl2u+4BmnatnSYUk
BsXsQljw8hdzWwCXX4UVCRJZQKglHP5ojDTh5at/X5xFZDMOlXDHPdKx+lUT4nQehNaLcswgW2qR
74JB+0KHWSm1vEv2RJHOKoIXdkjt7j8taJOZtmpgqLFqyzzw0yaVbQMQsRcXuESxHCyB458gDl8b
S3v6FaVIQriHuYYodm7DSKlUYLHidip7NZ64mIs2O8MHQc5iSOIus+OS9UIfc5GQK5b6OzfYX5uO
AGoKN7CNMeSDz/DBsuShDFJ888CVR7JJV2a9Itbpokmh/HB9mfGHBr9ki6KNO+UVv7lM8iENR1+1
m92gEk+r8xphWJW2NSe8T+y1owLDtXOOXELvq5nc6LRWkeZIOIO4d1osDTpMWsr4O7RyG0OqQOq2
4gybKskehtfcU4raZ7m+m5AxgaG9Y7uDtabG6djM0WnRGPvfARRJkotCHGpW4woTdqrX4vuAusvE
qTLp4vise/uo7OvA0+eYJxp0IA5wt+v/nuZrzN0dPCJ1gf5Hd0Oq1b4y9E4l62W42o3lTdp97bHs
KoBjTwQRdc/iPXDdlhRXoFIqzcw/koypwk3TVnzL3mrbTn/SfXoIJUgSWnBbAYqUdy9Afr8vSpxM
Xgi8wrPDZ7XG7ipWG7ZvZEmHdEyUP9URw2lQ6qmjc2SFg7lJoFtM3//gA1D/wjNJevSTzD00db3t
a3x7WVchELwPmNjqJrzi4UH18t3lChRQWqjPwhKN3L14UJ0H2tthQkfzabZpF+Yo5oNbhKyV9oc0
WyJs5YnuF31PcoXBFjLeqRUmNMKHqfN52PMX745CRosfx/74j/0h6VvzdJ/nR2GKANAf0JBXTqaJ
DXX1Y2J9iNYN61ZawWWs+rKub8NAF/FMwogQqFJJt9H0Cjb7mITVdZELH5DetE/Q71AmNkJzg37e
paJTTILFK5Lw1dqf1QR8Qv+MZImAqSoWIVvMlH59KGe3T1KTdObXSDCoKUExB5tkNP6QAMG1ilZ7
FDc3q0dpOh8J3AXcRKweCiHcLprTEH1pWu5QTE/cr3nat/H/kZfN9kSSg90U6XlMh1wOaPOF9Ctj
kMmAu8nRXDvL4JrvayrZeCSpOBFCa0boi+XFH+eL/+vKjxhGu1ymZIboYVOqhgINT8FlIAAmBQlZ
87euJBUi91ck9P/A8+m90OLG39Vfgk2ymgdFAf7Ep1TWq+KoO/SfD4v10HiuICQv+pDMYegJ5FjF
FKOyUrP9J8mTE0jVRuyZ9eEanBAabgWtRudCZQAnjngpQdN33iaU6xV8gqxSWRD/2Q7xl0XIAxi5
sL/eyQkqns7364laKF7jESR0KmN/PT0fRPo58VSJ3ptQybyqrELjt9MtPzfQ4H9IvcfHAXCT1jkh
YN2CKJB8uDaON2znocPvfjaRZ15c7+rzTEqaE8PdekQFKjAH8ezyq7UO3Ft6VL5nBKQs5ucGC/gL
5CtW6n8wNXIi4TdfXsDMLknxhZjYQkgEQWgK8fHlHiMCvMBjCayEmxPyb7pVeRJZU8XFSEqWJny7
+wEyD4N+5YQc0KQ1Tcfb5PL3J3yjj47Po7Drl5al1KP8Nua1D6C5PMo8c2EXPJSw5CljcLepASvT
3liAnVEkwrPLA4ZXxeNNbkXacBoCvXqIErfr/+/wOn45umxrTyL8tHUzmAuTf0/IETb4Dk3sYKIS
PiLAgam38j/sdzPhrRD7vb54p9UNKvy0QzhlUwJGY3SM2cL7OhUkN9foSOjWLxab8Pm9uIXdECPA
7L1gBwaL7eoVF6ygF7u9iAXXfVcDrfyGlTiRE4cp2mIrFnGVfne2Sp/kg2zs11B2FvOhQ9dnl7Ip
aN6hslqMp8cZw39eb5+UjW1Z/L0MrFYVN7UsZAEYghzMYf0AcwQF6mgj+9peFp7cHjznyQ+M5r+7
f6CRH1Yk/++9x3jinAREht5Vd9sz/ZeHGwK7ubyJAA1cyaRPNrcyTTgbUZBAJi+sUDDWGLJhcPhd
wRJFUU7bLNL3ktwtBJlJOCukvjYdDk7UQdLWXrJN/LEEhKBFQrRXsyMlr5CatHtbUxTgM07LxLkT
iVYrYcibAgn752NEZB07l7ym3WTLCSBG5VmTVMb2pUQKipREtq7xOkVv2UbdSUd+4eJLt6pM6+Md
AjF80eK2RgQfVG38TCFamGHPFkkkT/v2k+MIQifSz0GP4nixi8KnTuGXYfxgUiM3VokirIqNkTkD
2z7CwXN9+/IE5smOKnlx7SLcCahjmH1/QphKvTyZ95jrhligucbwVSpANJvpDictVePn0SutOVVF
HRuUXsRgqirCyqOA342qg5wDUicjbMb1KCk4+1n0WwEQfOIpZhYg0yL9Y1nplGB0+6ul/T8fIKGW
ikTaAN0YI7lPDwyu0xOqsX8YP02NgPZfFyhsvNM+tni0uhVTSB/hpb/7d5dQwjT7UuvQAgGvEjnn
wIIU0bOJ47+WKgq02bd3NYUvlR1UyFRsVo/sOF8TrFMxRx3WdjZo2hGhjg61vzwRGLNAe7PVM/m7
GXZAOoXC/YwygTjsebb3mBujVnP/vQFqUa1T+2QtkcB//rgHe5YcxGuGsoO6SCVit499HNHfvnJX
dxRraZdEKe3Gkrg7VZB5q9/tp/AwyAK0hWxu0unQQWrgYoi+QTAOilglC0xH3uoDDd4LYhSjJx//
E8jDF5gGbCa+qhjBZsR02XaBFQBBcgAkzPxyWh5j2XE8/YsdUmBBvfl8mymqmknI1rEVPdJfklMR
E9HRG9DPhrIvXYa7s5xRmPizm2IAtic5cnmHDJddf2zstv3bCLgZcXUCmvy9baGMdzGvk0/8yam5
26qkCyoAyf78rRiASYGyB6RP+9+o+x2fbgTXviqoPqtQTla9UR/JNIklFn/9LqNDkaqs3TKOPy4c
5WcfcGedrnmI5vsGD4D6VSclc+TiY7Vzu/Umrk26bPAFkBFn9VILbkQVjcSztFOSNsrwj34Y3D6S
wCwnCoahI7KqLj5U6M6HJlAJrLDXWZ0eASkGQY0Uir4hjygfQj6sN6wr9IIYT4ZhJPs5XnrTqjSw
LldwuNmOTKqxSKYfKYgo8+0oOAoclO/3BWsIGZk2EM11WCG8ZOrLR57750k+yDdYt2F8XxOa+r2n
AY9iVoPayxXawLsPPIZMq0zxU8K/XAHiSS5kR8GPuWRLFqxlHNkcMYb4SMPjk0TN/tUrMU0zsD/i
w5h9iUhioZqlN+oumX0IMt3MUXLyOSGOWkfY7Mkyn9HId0eC/wfguwLT4Jb09CmynfGFtbs+//zq
ymfE0URWooGlXKCr6V3G1aBHe5hpUk7nLz//CCEZaKuUyd8rR8iLnkTDwbrt398iMxpanhukcEu8
m/r+yySKmDux6rR3IfyDDhnjmpIm573oe2QYn3nTXuop52ImjUEFcS3QtS6qpbiNZmQ4Dsx4pSHC
RizNe479VKxXgd61VyOgOgKPukGCOwmFMOmJ+KuAx4CldYhK4Ojpp9VdZ4viTq0/fcoDWoCg89B+
yTNwn5emSBqn3hlRWwZJY++evUrgH7NPvmim67MhYkHeXy6YJnyN91dOIyDCtEF4Yg87jI1som3v
6yi6OLc4n+v7/Mh74bAKMlKc/990ODqv5Eh2Sx+FiY7ciEPZvK2nOQ1pR5/nVSgAdckrajch5TN0
1tj6TfnpATVvX7Dv0Nqb+aLL08JPer2vFF8rhAmqkgPmCP75jHodpiiC+FMys00tXkdjxQ7OopQy
xoktDtLXzYWhnFeUQwBy9hXpZRRFnao5brFg/e9o7kKbtyAArRL7TvUNfP6eDsvo5zkYnJ5WlVWE
AKwN+vWd41ZIuzf7oY9l5uhjcW+k7D0qKtBpgcbG90HTzjOlemJX/84CBBUQMVe+Sw5XkpLqSV86
3yuMyoMJ4I04tggRkaqECldpHw6j5tyTsrRTSH1TXMtWdOJev8X8b0d9JjFc+HMYjJp1SAfCMHv9
+BhfCjTQ5wQ+WHoZLU96ucw7wReL5EWNqPNVctuzORlG8RCB3GMGUsNQevjnFxw3p2Ga43eTjqii
QoOz6ynLZNi18MdxqKozAogPMYge9HM0WicGTupoEgn6UhpJCYEdijCV+gWkk31zLM43iAHIlLZY
J3CS0u+xwzBXM+9hxurnrOCuu0KaPfqMh5qTVVDo7L1JLbxuervFcWXNcUExapKnD253pVppQiVv
Q2ovaoktshwFWffhuXsQXfVfZ7qjAdYulFFi8IVGHUL86UAP+KkRBNQEs5iMS1Ea1M6uYWUEirYr
ZKtE6AqPfIxY26TFK66/L5soPbTPmCywsEgQf/5YLvzdQPMfit0M/Bdqxq+kRfGLuBjgbhWguxfA
gJUsggBth41XG0o0FgL7bKKh1BzgRjKww53Xm4cXGeutiLzYBh+RFlz3Iihjv5nSlf/RPkes6g2J
+Nqus7VDp6S+hP3Z3oanc9rwLO4ZJ2ZaI0O1lg29o8fbz4Ns1EhA7bp4/dwpjCDS6vzw2XeCf/a5
nTSUZyKF1pubchpBE+OJo6fFFallLN9MuouQjByQoZxZ1ZVNApYxZpa237KLAMTv2vPLgX/WKe/Y
pvXo2nw7AGZW76W6y/wGtZ5OtlRvt83Z7CQw1EqvMjmihrp5AaJ6eAqz92IJsbJb82xLAbw/Wfbk
d2f0GpnIfhG7AMa81KP+rxgPPCvn9qgTFrYqqM9j0JUvNPomUilqC8Tmlxo8ToNkgX3sJxEy1gbL
Xp4ovg0jHIqZBHIHRlvRJmr/AECRn1Dh2rlk4CD5MSEuKCMYnVdlW+pZNhf29QMZwPNmQX3pdL0q
EvzjGPFYI3g4sn/PUOSz8zmBnKBiuaY4TIyjtqlVyso3qVaNpV38UodlQzmBXZvmJTHq09Z5G7iT
JZP0QQqFeOIUDdxTkvNzUfuQJ1IsszDpjDv0B5cL0Va5cjsymcjjb635chBOhbI1MTqs+x9eX/xj
iG/+sB50VYkTwgngrS1OSGxx1ONvI7EwJBCnjK/Y0xUK47qIgCQDgRxJ9HKnOSdoCBja5thp00pZ
dN6f8Fe/v3aPguG8XyMZGI5wvmTW22g4nUPAWEyfVoxCryFK1mGPNNKAmOmxwsV4jHR8I4peqeQk
y1kXCPUCLxxFfNhEEEOBUqLODfUTXH5pntQVJvoWs39RNfSkH9XQzizmFI5m9dVprNHGeR6n6uqF
VAEl9nORx1rtqnCdlGfc21uaR8L9GSmIhP67+QKFggLdxPCFIfIXn8SvVlwSJo3wa5IKEahMY5Yb
lFks7gkrm1bzEweLqB7AZ38ZLBl1VJOzFs42+FBURp4aeHZGnj0Sxt5U26DSmr9KCoupfByDp/Jl
DHRrgJPv+BzIUqF1uKTkc2YX+KjuI/lIm/YkP2CMLNaX4y15Glx0BIOqAHugzUgyAjeT8jegaAP4
0CFLf0YZZ58jnXpCukRdBmGYSVIptpUbeomUMXYxU44pNOLypeV3ndol97bNuDTt6O7KPUr7H7CD
/3NJU3n2RZJp4wGJ57MgaeOznU735CuRtT84u+x2Q4tcbBitkZ6+J17Vuqzv0oFnzRxUZU7Dk4Sf
qi2XLZd8xXNkF8hMOydm+wRxsVIqFxZM6h99pW6y5plmxmtlrA1gUw1lWuyRQP9HGl5GIZ6CfpWh
wrklQkqQFsRQ0q5hTyqupPJsNBSpub+myA8wEAtFVBzza636e0V7TFRIIIKX7qHguIIVrzxu003a
sJSA+U2BsvClfjWSk18bWxeIjvKk8TzVYuFyqnjcnptnKbh05hQ+tP8f1/bCUqYqg8ilgvoNW2EA
Y+wyPP/8pFMl/resG2o7xT2Ff9Utwfql54hup3A9wu3oftoNOL/5lZROTnMh3VxjTOJBbhm81Cfr
o+PTLSbmGmn2sO7/h4fYGIotJM9gty/f88MWD+lbktz8U2HVK0Cj5jrAowoncXrwmaMmWPVh3ni+
KD4fqninPM5WswM6ITkG70c3SZ9d5qVdIoodLob5kBSl3qZoTSGHDvFXDo1FoAAvc8YgWfCG9jKc
LbzoJfPxSZLuCviRL2Hv+/g+OamCvdsWoe5E8EkXyg5Asmer6bL2uib5lR/b03M4ik/wvg2VD3uu
LIO8gYcoZ8WWjOKCNW+exLpMZmbLLtZG+1cz7SxYl+LIl4fgsHoRMkOAxXBo+kZAtUhldcajTwCS
3JHWtTiuuYkbLCaiY9EJv7vLrzxyfAUr1SDMIA/tE6ZvC/OMchF1UqVOKUrNKLcA3hs8z4WFk7dF
kckIeOovfOUWcYapOK583y3KPZxvMXczkOqJW9CC2pQlg6Q9Of7FwkDQNAL/7z/nY46TTbroboxp
rEPyZFkjuxo3QhC9KwX3vQEEwEPcPNsgAjDexo9q65zr5+1PPbmScV2FnI2P5pqmzZkZKVO+0mSw
lR71z+3taxkd29wToDsAhB+7Ohgbn5hPFD646DV6xxzKXDZTh+D0ohQa3A4k9hUJ9yYFBUXPSggm
K47rit57hi+A6yRYT9FjIf4B2V4xn3SekWx1acwxy7Jb9W4JMdI6ePCm/PuDrJjP+uvuCefY5YQ7
38HGlJBW5lHFMN4hqznPo/EN2xHwTyGNh6qDbrGEIFt/fKOmOQcaghgJ8tyAna01Zl3SBxdHPV3Z
AdndKDrdOvcT/wSFmUiVaKGJsavIZJOlEeCtsctzNQy7MPxNHMP8RQgK71vbl8dK+w3smo6l0z+k
6QUnjazZ52hVY/lTVh/7tRM/wdl3zMM85jMiwC+4woh798y4KTKetTFQXMWPcqUNAgLG2hAkLGej
TM5RNCZr9TtFDH1izRuFDT19jq7m/8kzLj3N7PArJ6R1r2DEj9bf/wdsaKapfWOi+Rfp5cjfoMMF
PwCpxfFP2F7aV4DuTkgGXGpefXcg2rw1VHqi/xaCteAGvINeQNHlEbKKIFNkrNWdaEvK8Tg4Nzas
rOjDCfgo8KZOCbdrxgNRFL4Yk868Sl81ZpLHOW+kvH1TOjsF6MZMBQjfUgRwTE0MxRLkk4uTfIkb
XDY9lk9Ao7EqI85VTeeDvvRmLnF476jg3In+aqeOvIp3YbE368C8HF/Gw3HDEgIPWu3rBW0914T1
VxI4m1xb4GzSbd4Pd0RWdTO3vtHQ9V4VPCr8fi7krlEZX5liK9PenMEgkkcrIcBHsTYaWOrYbKkh
v/UJIQDLI+u08gy4WwSYDgzZAPnCLVE/JgFn3bEZjqQgH5fMMaB5TQHZmyxVnDH23Z/LcufIOIca
OIDAie7PwuNcfXKymXQ8hu7jF8fX3R6vt8WFEsYnWA00O0Yg9pVk8Qmmvmhv0hi89ju5qp2+4/cN
ksqHa+LywPn6s/23WTbdEBBwqxnZQ3aKcAs2GTjePnB++H9jQM4pz5WvxFcJuE4D+CwXlq2c2pmb
ntF/+2VS4h9QvYZoF27SbZaNny2v/117epmnLKhgUEwphAjsnXv9jDfWUA10adEqzxs0akmjJ/p2
Ym2ngAuJ7HotpcQMWVEZX0seJOzhZxJrQP4krY3GBahzQQVbLn/zYCt/RM60+t6r/M7s8THU7EtP
Xd3lOULksVfPpz2/4x/eXNdolJVuorM0DiNTuRucSjQZ7hItKK1VB1bx2pJz1B7+9VxKhEyj6Zt6
lxxRRSdGEcM9qYUl6OcnuuoYOzqk5cveQVNlpf7lH8CdD0tE
`pragma protect end_protected
