`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19472)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCTcg9EscIq6lRv0lzTzbJat7rHahSqjIbU3zFXiUiLyB4p19hmBlf2kO
ErXmO+zyUrpHtH+vFEB+9S+DMlDFTzSLVQ3QtCqoAblsgowCZSzhkjhXV5hMnIYrDnTVcjlWtnvB
xB/lQaYGwuoCH0QRY7IkHh+lSpKLQWe4v8644boHQib27VFxhW/IMk+xSTaT6UBY8hDxuzhEVDw9
+9NhTWehM4TUujW75MoWQioY6XqYPslz8EldiNGMRgx+jASP19Cr+5MVPH3ZNbr9WwNZi19t2CqH
227v6DhfcSd35hCD0NXI6uxbe+oZ7i895Ag81p2TeMcCwZ9FOAKlMV77aLRwtiBZMR2/q0BBQAwT
bil/sSqzZA7nG8nW4fdyTnLpknTbW2CiuUVmjRrBvvBp4i2XEKQb5B/aA9mlk5xpacP6yAtjGCnu
5kMJLcMAjZ2MSthtVNaooqVlqpTOt97Fo+oY4iSFjdvXaI0s80C5JiWLK1fXIwGhu1sb0IZSBfBe
q9kcdJRcS/x5fPpXCZOZbr56lU1C8a3ObdFTuO540LKjzfLgfrSZRxTGkIPkWm+Oj5VszJeQwACH
i/TQfrHJiMTctgM1yaAZxieTzrnQm7vCkbgGG749Ae8+l8oWcZoQ0acbGWKU+YjiU0rv/XMqypmD
4aopSM047MxIUuAsdDL77wETVUECdiVBOHvwBGesSosBJYLW92z3g8uV9pKT2OO0s06mxg+sS9UB
yEISa1HFw1nlGdQu8AkMSZOhh0JsvMl7pbKMsv2CiLzBaUiCFM18CxalWJjSBSE/SPz883N3Guyx
biP7f61eUjqL762a31tRKzOEwDqFVjTcJSjOVwB/gY0+L45hdDCmwR0/rF953csD7F+uVMDQSq09
BSA9bXJSSDBWv9RlRbqLJGW+BcqsTwOKMRWZiwqMGru71dFC0JT4AW1d6Y5lFJnVCxLkdAQjQabg
4rO1fMb6ULOa+BzQMOaEkIUNhqBSoUeA6fWnDdYul9HAlbUgaRWx9gfjPV7yyzIb2WhVk9rx1EWI
7pNPAWQ0tpP157LpQZAFbsqZbZ2wE0Twiso7OCRVM/EmAxPwvOz5qvsvYORQGscxld9Y2a8SYeDO
rYv9d7Kim6xnaopowuDOiW+GgbsIhzoGWxXMxxkX3aqzaqiJ60ev6Wn5n/teTvWJfcb0zzWbnlDE
JTN/bW2lAH7xdSWsoskGM9e4hSGX/58LgZWSf7+NQv+/ZA7eRAVUePtxq0wWXihCTd/PHjeu1OAz
Z69WzFsnchFv9B7LLfktBcyWjKsEQo4dBgw7PRNV/rzuMkT/3ca3kClTnGCkqcSri6xNk7SKskl1
Cnm5AFOaH9hE5Cp52fiMFW48SzIE3oKXLVNR4Hlg8nwS8Phyq1JWR04ABrXxh+Nt7HlSEh0Qlrwl
uzkA27+2OswEVgRCcbnte+MPYq8Zo8svQadGiYngJ3RFnCl2tXnXZ6BCWFqLuKQUheSRVXjafgKN
fFvMFG7VVQULdkAOn4AKCuyYQgSUXZ4948c5jf+5GedTjT9jpqe5njRujCT9JYXFg7KCXbwENAIJ
Gb9X9w5m17BBNqNuCZ0ltCtB0VZlXrpv+spEiJhH2+yvD1ODsfIYT8t9fmx7I32BfJBg1fsIgTwy
g35UBBZ3xOhUcijB0DHDG2dd7c0Sm0lWfJDWapZPmeXKopS8KJ2p/s5PcxuF5TOFzRv6bEaGIDea
g1cojefoo/rQWTMfBM1cP0kUSKNhGvpXJg8YZX6nE3gDnXMGstcO05iRlGk+jetTeo4GuAZn2hbw
oIg8XytvnPZhp7IyY/iHyP0ITQqGHm9atDF+OynhcnI2ewGFDc6zCOd7Dfodo9OHmcUbeSCJ4BBw
DRTJQRGhFSv1BBYVwG2sdyGL0oFrQJjKGCTwc/WVG64fZGcL1CyXO4XLd2y5vO1KbBo/DDxLuT6m
Ic/3YU4795S7vqy2aS9IOB5lyKhyW/98n92tU6eTSJKXaCpjSHJY0JEbdzKppbLWzG9X/eFnxj6l
yqmnmhWIRZWNf4aGrZ1fo/7wIjrYbMb6eibaCt+Xj+YAGQksIcDAVhPCu95e0u5CObY25jvoxLlR
3UCnn3izl12As+9gRc5LuhB4t4xczNbgTs308MVb5eRR8OP/tpiS4HygV690g18X70sklxCTFAk0
y4T15TNPuUE3iO9gg0QYjoMMtxiZhyb2NtHRWQpPoMahLu8JFccnDViJGIkCDsxvnMjyTONzJDPA
TZNbiwsgyknlJvKQ+XN7NhhjfSrfOfE2XDdUBWMN5XnIFhqB7ZXKItOwxSE8wfZY2OH+LTl/HD/3
QVL/PxeJO4UsEzcqd4tiVghA2qLlJS0L0+QUo07IMpn6Tnw+i+V6O996xP3lLjQH9xYk1hAGyLuM
uvCBbYuIEKi05j5JrU75xzwljxFDSg2v4EZmDnFERkIY60blLDdZAHvBgQryCIdyWZSnrw6hHv3g
ePuIuLCX2Irx/zPoBVhMxs+f6d5M4nIdQPimjeZWHM5lZo5Zmpbrs2kbXgSbrCeZFOS+110ZCJRe
3zOJ4/zMDIFWtbRauJ03sKIrfuO3F2tI3wukclIcE1zrrIcKQO6mSOS48BExySMJ9jmFwzM/yQMk
WOrPGIBadgAt8jYearAHbQqW6U/A5XTJcFW9i0aC0GGdiTTeP/wsrVWePpVKs8iAw6TRp9c4DjZM
7pNiwoojDAxmlZgHS5J/TWQnVq0zOWWYIMok8TttWJ8MFvdSWdHpncX5LCfzXmI0wbqTSaiQqZbl
70CL5wa8bGZf/vbTuvf2RsueWP/CWNTueRHUvT8AHARNcBi8denarv2YiVKQDGuv07lKwmpTjkQ/
nRrOv/L0Cet4cGFGT36VHv3A7BE9uMf+hbXpRASDiVCt//cVO4PdJ5db8RBmVWz95dZ+bAIigkUh
vcUfZQ370qBsDmjsvqDhXgrfssr7VRpSwE0tmITZlYd/VdAZe1ZgJ0DoLd5hE3tqpXX/jvudTOn+
qz1WIZ3SZRcqgtUrBKBFcSYiECA27GSgzT8wthFQtTPHFdIHv5SZEji3+zE1IE7hLTjLC2k6YXTn
8wYPylFeBj/sbJFaWRP2gpPjBiy6xQsCcitNbp+VYvtJ32KL3lM5qrw0OgM5xwNFGduES7pQ2f/r
xRzaRJd40kgmTQUjI2ZCw5fm2mSKAZ8GWseVToNg76QXPZT/tf2hBgYleRCVSKUpF7rjBrHYY6xj
uajS+P5X+T5Xkv0VJflIs2h3SQmaH+uFQUVpZZ01Nw+UtbF7PKPntS2y8lUACW01lwp2+73vXqy4
Boh3GKQ1LyMvWKtaHS3Hp9/zxVdKmlGyz2pqfTuVwFzNUEIjeC/4GgNT8G14eJqnDBcuVtzGBcOr
QDXER+XeXdHjV570vXHLrDphIJPksYHyzRP3TZglpjToPo3ZPvVsiuZKAM2YuILBdvEYdv7zBgEY
VBkHwjj3ANW+mi22LArLtmwzkRAJp9Ij7foCN6e7dgzgyi7Qo0VJdGFRT8CsR47IMDPaIOX0qDpw
TsUVZ05yOZHVh2Uy03nHVVtaymkXpDy4mQn5AbkpkExo8lOJYTl2xNEPem0T1AoebNrQ5kUSfGcd
N2lLEkd/TZgc5PPqqhq/tneWI48c3bwM5gNEaHrB9Z0JOmlt6m46hBEh6B3JNlE6b7uWOfCs/eMk
wNm8ubqqZRgxmpaLhe8LVLXdUGKTyheN+C/B/TC+LzYgoPWOBNFY8mfpu/+cixv+qX8s38QhJfzr
sS9Z5V9TfXaIlIcWpOLYFofIp69qRi/DLmYP5UsPKM9s2USKshXwACXc/cLWWSJP7YupLN7bU4dK
9aiVc+nZDtWT+SA2PASj3hSfhOZ9jGWNfEhEsPy0tkCDB2WIhN9eQNk7sKms4cMBKfo4slkbvTPz
qRm56oVHvh8pbW5Dufndik2ZqhYsGAi9knujfFad7tJXA2+fsXsq/NtB366XlkhhR0wGy0NojmuH
P1QyraSQ8Tmez+2rAxKVnMTsZeULi6QQx5+lfn1sKL/egkXgmc5sPAK+FSD/wBuS4xSiPUO7WwRA
+KmSQcoJmeqZF0jvc3vWxW/W2OUj+rjY+ovSCH1Y7rnrEIqSQbGa4yeM8CHNJcje0AKCCjJYy8uN
wRdHy9C8mzMugnpbfMVoThTZxONXd8x5+9erIxazwKAzTqZycf9tzddTbNj7ePCkhIA9EbCIMvFn
XGiO9bfmrxlyKMBj9pXb4aBdjkoVz4vdt9rH/0G8jaFooXN0lGG64gDXHtYGzLwKhxVR7kQ11gCk
MV4FDRhkB5MjK0AzX26Na2oiGXrJYkBiBYbjCX56/4aVlPVUaXAmGZBgVdKcNDt5XR0SYae0RqsO
wLGs/wgZcwAuSOIeAYVNW1COw92ahBcD6WYcjuripLGvz9RQDN94VMEld1FWYN/TPzVqjG8FbK8I
FktKVAQNFTxaMrM2j07Kjee1bbW3ddSUQnIQWTYunGCK3cWgnpZQthxUxKekMBgqku6CqvfGKZZz
yVzcelSbtDP0LzBAMDLho5HSLY86XAzGx0CQ5yOh009tffem96Vtipt/csmNnvxK4BrIwyD2ayAg
GWf1qUTnBiK8hbISQLOwhU4GMWAKuZ06i2zpFwLPkXOdXr42M+cZFWCwRo4r6yRsOoETrfgabnzV
JUe49l7xRMiVPz7O4+jdAtCH2AoL0AOI6I6mFkk3p8sRJiYO6ctIJA3lLxnAsron2BzXkeNZd0lF
nx2Q6wFAKgQw8uzCXNOSQnaHlnWEtbcpDGU8z/Tx91aBqoBtDJa6Rj4Jw9G/bBTNz8cYfWk+91Rb
AuFCw3Xmw+O82uIIercD2xeiAeVlEXH3FV9nsCeB5+gEbjr05Ty8tGx5/RnGbfw1lhflmq5s/h+G
zJ2V7OiwXXq6PyR8zmgQp44m47jGfUz3+ngLIBS+yWDWbJG+VE6MP3JNBl7mxJBX+C4shduRNbgF
ckwiGZ06u3wo0LRomUb8m/6uHuA/hdSqZvIbekbz6hqiHPS3URB9swOPz3TAn9eUVQN2qQ/tyQzl
I8ZbQP5GuIrMH123fGN4WdJnJygc/SL9x+XJwy/ttXlzOSgnbKrb+iP5Ov0gCi9OL+dYqnpTkXbB
wdRoiVN5AVXBakOVgoFjC9HdJGhzvkodrOKh7uB5e2gTF4s7ghnBNoOvPZ4pUxnzNG+ff15SXJNw
vMKCg518pDYMb2gGn2owel0AGt+KxI3DyRGT9oC0m05G+Kt3a4rekaGVa1KER9t6EJjhZWMGSOS1
rQqyJmOnSWLRRmv1e7kCl9TQgV1FPV+QgOJra0P2+WHRRlxCM/3rufnXNuks8siApXSaRwk9f+jJ
BByBZ47AdHfmueXPAAMcEBUvKabLqc+vcyT2HEhCYnvE/F1bb5K4lNk/y84N86Bxw9tpiDW3O4cg
gI0Lo7AY8AqQDipHxVLPYMPUH+uTJi+fB0KlWIbdT9sgesc9VsBCvlMOiuuHsYpyfRF1St9nwpTH
cwhuSI1wzHszfcgImfhZa9K/Q+tlZkuLHX7IgizwEeseY3oZClKtlaRN8Be57kwRlWJDuXJ4VIZ2
RGF8b57JToJ74ISFPmRg8BJTYfsn0ebqaIgkSBYgReob6jZKQ181ohvkABiuRDsO92XiUHp4IWK7
pKdTdmp+scwagWzmEr/eBU2SBQfW55uxx7HJcNM3nDpyYGhtoHIluQrTbXAl0qjbmIiGJBBQJfKV
Cd4aD3FHSw+wZHng6K3P30SQVrXzt5OrvLNJEqtcOlyyeTJzN/MGNN6v1jHGSYe7KC7XcIEzo4Et
dp3ajFblO6diV5TNO8izYI/heCxzyoKg3UnGuc4mjs30KattASbWs47rsMFbzKvBcSM9ukaJ5zhO
8TbfY7uft9WU32L/807SWXx0szM44RjOJlAfePYlcCfxzrBoMfbXE0DMVDohGABSzudydrkibVH6
6lehS7GKImaUlwZoDpSdwydC4v/PTPqx8VMg7DV0a0N2eB92/h5Jm64tvZjo/kpSMaEsbkCVtH+l
+2GMmMjIoqlJJ1R6yFrGDmP9hh14RqB7UtbAVPH4LBv/IaWJW88M4E6JrA/zLjxxhoTvXuyAKgRJ
xNxxsw6Up0y/qhFCBpi6cwjWnEod0d9D8+ZNili4i2ozU4MbdKpL7ghotF2irOmLGEUxH/Gg1RgP
h6KlPmAnCNEdCV+DqS58qjZ24WraGKRqwRO+isuPrEfZ5pt021pP5ib0CkLex+9dv8ox2YmjvCIM
uu8lxlm+LGegIgCNJRaxYgF6SEbI7tkY8aDvF1bRCL+CTPYVLTDT6IY2IWL2CMoB09jWqi0HvJNP
R5+l3kKRFomRk3cbb7Plvwj66G1f4B6ZZyjmL7mjb8tNBaSpEmytK6QW19pioUuucHhAssaQsAt2
Vsj9eqP4bL0I13/lnW9zqT48RbCB1MEI+yFyJ+PInIHyCrlRHHJDF5LjrBsu7uz1L1rjA6uD6yPu
/WnQYYOetFAVuVcrbtIcPF0e7fm10U4LP0sdQ4ltPQmSq5ly1IYXZ4glFCI24yNbEUn5wMT8XgBx
pCG2PDrCrYKnRQWDKn+pFF63d3ud4luCg/FyysUN9Hy8d0GBJgpg80/8i40YMT1qSEFekJElDq1C
sOs3IxjfK0E446NRwto1aGo6Wv35XyY66+ZwOG7ltjcdM32jFilktxTqvd//9sYknEjAsvvM6BDC
rK9CQ+3THF9UMHBbyVW1+xIe9FwtOyiM2b+VH2E8B76G8FyDERmZg9O1ImCPLP5BF8wA2CI41t/f
Vxr2gXNxfZMKllyNeWP0sc4jN4O6HCaFkav7UNYXaclGH4+fVtxooO1XvqS/zntzbehfR0AUJr+H
woeZ+P7rWteksIaX/u7WkwhV1fielY+ybyYUD0uuRy6HeMokefRGVn2G2pcNxc6S94v28mzjrmSS
S0RstTX0chgxCxGxefD+vfoMgRNny6DIx9zkzBg/r6QTqs9fchJFKA2QZ9auiUBUTDszOpXGICET
9rrLdSjp/HYFoSKNIwY+QRKZtgqYbttpokd52q/rWIoFg4zxR8IjGVbsQLdlrUCZWC4b9lGhBUBT
9VILKgI2qeGKGlwXQkxFIpzjVV4tY9gqPUgiS8MYXgXP9PMWoAV7OgsnK2G5GqANQilaiIMYSQ31
1c4K0IDXK6Xtsu+KYubk/l2tow6rFXVSraO8Ssy51QFIFJqhpSLGDnWhvdAsqYNaL47+rT0mqGe3
LoxAHljV1r5nPVZZNjJzTTixBHOh4IF32dLrG3x9a0mOTRZ0BxmzGPaBdJu2XvsxY3MtIjrr/+PP
l6wjtGgFPG90Z69jZMS6YA9RcJ9HK+QPbckZn+UMnS6QmscGND3QIp5jgzBz/XUwhNJR4ZFyAh6l
e8xlZSVkqLQut54kPj7J8A/bG5QGykp0iBLY7Q/z1uC1uyx7P+ISvEDJKk3dlMPbvn26DXSowjlg
RHVj4MCsgRyvFgMFOkWWq6mtn5U27PHG+PE0s0PQ12YX2NWqS2ZSgUBRpjVi+rgXBcXyaEFHEBrL
jS0SwDe66QL56T2MibMlMvG1xOsso/oVVhzMdmbORmTdMEEEpob8n5j1d8QFLvNriBLnnCKnd1Uf
wr+vds/li6yfZxhLoYe/sFLdKwzP5dW0ba7e4GRdgzx7HCn4KuWToXp980/Y95iQVwAYVvC1lx+7
DSTUHKHfxP1q77W4/ebDXqSX0nW1aXsEzUufPUOmvSpOZ4HT4o8gIFy8yldAHs6gnU6Fp785ee6P
sy8VJz5XHaWmD49CGDrSjl3BBUjIrT2GYG18/6jRX49hcXb9WwwKKLoHSRkGXEcvPinB9r929xyQ
Q2Zw+EIc+tBUXeWHQ4E6Kaqil1W+5lJaG82TfDUZXiEnj1DxpYcoN78czZqU++1MKh3CCRNcsAyT
uEV3MTMtM2S43dqN6MkaCAeUtsEH1Ltglst5nLFI/fTrEcP/8FWCOG6Ir/yquUjtb0BII8BVNSTV
WH4ZiEO60W6YkQxFATPBjO3OdX+Nxne2GVm7iCLQwWAu319ATyBhtH0pPzfVSIRV5+/uvwcqOqJS
3o+eBhpxogZL0ffChpQYpAJUHRIAdT6oKA2yYgtW0lWAcfU/N7axpmuBqOE6yihc6YL7U//hcZXN
U6S5nnAZ7qV+5Rc1S3Xclm80SaT6FXsa2fTs2vmkUWEznvIdatOVQEpEwEU6bC8e6gvEDnb85ogK
+au5fdWEbPi1qtdml6FTQ1rOGA694buuNaAuJ8MQYLT+51zDz7au5uiW4FfQIJUEccTrdKiRjiTl
WGkCSE0OR/Pl9C/XmZJIoaoS7Cx7GhbtuBY1kyjUWE+MbEbjZx2F81poMRRCZ5sZbnEsY8AkS9e8
CC3BbWGVr1cwqSRXvnCc9ni0Os5DvdTCkxLBsUp/3I1bSCOl0gYRiW/USB1OpV9ScYbFMLJ2lcLL
4mqhCVzjG7J1LC5Hy0gRV/KlQqrAAKaAT5aEeqYhH9SoxyCov53b7WUbmDxFSQxskFjD8JReyH8s
ZoD20JaVX2n5mH++hZnMNgNCTlxMMFV0kYLX7XwBf7EdU018GNTTuS5FJhr/Xxj3q5eoVD2YvWYP
IPVShXT2e9xiI9YeaUra3/wHfwHd+FDdDVB3u3LeILrR3M1t1FuHfvBjQp2+wlsz/v6Dyqgr+//X
QtafVJtUKYbY/TvrllPO1g0Nyvg6WWTnpm4/wzKzCrPXZ5cQiSO0Hq5/bAFbmAKnIS+/NWZTrG+O
lDJzBkfHUDbSSJCGcuScaUwEVLiVoTcRSWX0KwrEt8czUuJJG7iq0H3Q/Yvfsz9wfoT7k5GpiGo/
36rGrZsZ+w0SwMD3GVwsUraGLIPF+5Ls8QpQoBEXRRX2OicsRwpn+4ngpmuZHq/GjyZVm2QBDgi2
p+RtVtEUFeNbK86elSap/tAggtdMWsDWLugNLbDeo+PzHnSfEh0oisjDsZelmSR5XAY7TUduv7mF
x12JljRK8UPrULY7c4QlmeFlvAws8m5pYHXQxkiI9Vh9C4/zF7jLtXL/qiZKyywP03Syg76KKQ0+
1eW8e8Q2uXVOa3K5d3MN1O2yS+fwjFEOUwNPhP/er6lz4a9R79MuCr+A0chrNWfm44Vaa8XeQCkT
H5xBH7BpQjNyvtR4qrwUZqXHxIW3tb1WspXCXwDZtnm87G+eOzADg51fkI5188H/FcVoZc2tAsx6
SEzWxToiF3+Pinq93c4PK/UoMFdtfqy5PrsO9Teo5gMou9vBH/JRNE0hAhCuvFDngZI//B5ZFA/r
m+20n7qpJ+EtOAqiR8qDSy10VsqGbSUp7/CqUN8n+vBE6MRyMo/22UEzRbY0i4j4btfEr5BayryT
7kJUiSlU1lY8fjpqzsmVMixeGBRH+mF+V+mgFMStCS7YVsMHO0pkdgAtjcH5CS1d85KB5iJ6Qdym
piT0FzlClR+0b85dXPYLykaQ/0C44aTKKnkZJaZVW1Vb7d5rudO45Ku9bkGqwOF/1s5DPzqYnjhK
hoDeqzHZKfGukT4PDrhoNckcspyV818vU5NVQe/Zo0MR2a20tw0U7aMNdAXO08pWdrbCi36Lkp2R
nL28a3TG7k7dP8YhlT6ygKX7yy9CnLrXAj38xv9j1ual5Qjwer8R3Pcnx/Zu31WYPN+Zi/8RxPFZ
ovaR+FqHFN0fT4okgkN12iVjVgHyH2FR7QtNpZThpZYgkOe0LcWwtRhWGlcgjTxtASnQlDTjlCSS
1w9PTou6EOwkM998nU8XugZmpCNRus1mtmQTO3A2puYljdqcEahHSK8tCS3ym6Aabocq3m9Z+t+a
7jbMb6VsOBlZO5TL2OG59vNKeu8Eiq3qQwojhjU3sypYXF05uiZDJsPH2HhDN2OKmm1oFilTAgsZ
AHjbbfQQPheqA2uS5R4SrBLMzWLw8H61yWbKLuP8g17PRLOe/hqydE2go1RNfc/K9gUiHhzkz+O1
McaXq5tUxRssJiCnhl0fncAMh7RkIB0Qkc8Cl0vTRBC10sr7KFdd95BseumSKShTMs+roIFdDJGj
u0nSpH00YDXGoyUchdXzw2k2QGydUUo0/p5dFlPh0N4wNpDwMrK1l8dyeHpJp/8AnbgHI1XODaci
/4fzWcEaV2q4+AcVJXgMZrLhrSLwxgrKFj42wtgwBHaDEJTYv/NXQCaSpyAQAuE9P9Jw4H2mij7W
n4ept4t6TKd0GTrEalSWFnLvtvyxCeM0/10Ja0D/HW/XTkl9+JYfV1VtZ6WApjcOxtSmRnNBBxu2
BlDz+awlTC9OtEJMPc7Nxa3JobR4YlZupwvQnvqLlUMHT0yyypQn1rvxJu6dPTBb2dUeY7M3D2ux
ULLQazhSb2/WdyoiraU3fgdHnqcGqfVr+2u0KyMBXy2JM0CNdnXRNoknt/QIICJsBfFEvZgdM3FG
6xdd5xNUwACHy1fsVoMcpT68KcOTOQ/a7zK16TKFrXoCpu0UHAlfWEMDy+RcyRhxBZBT7NTKH6pX
zWH+32xxe20PJ6NwgZVmIW6cot5laY1l35ODwJTJZHXc1lX8cjZFBwIYZb5IKqB0a3WTlFBOWHum
KITMuMiQ+WjzlgTD/3jr9nu4Oh3G6+pkTPSly1JdF7sbw7wTcmqY9k8JcXtrXSi0QaDCclrVHfMj
KgDfiHBdrVngPKWxk/j8chf4HTTHvgRbQ/vAJNC+TYIGsvRjXFY+OuHS5Pz93KtermrUOj5vJMTG
xygvbs3RkV++v05h4wfSUeGbTz+fFEPE79li0ZYV1T+sANWtAm61/6pnYKIMTqtba7YACbiRYCWD
i/DBodKQPpvFpWC7TgL/7omO3ok2aISMmPCe0404NNKzEYSX2QQkS5yESfOS4mkHMqYwFxFNAZL1
QqIJOzoByBJT9rPnIginvzJ/ZvZmjNWVpN1AyWCP21iTswmdrLjl/cGrtm3a96LOaEUtK9T6lSHT
vS8iqqiXf4Yh3zwKYGjmKCOSYWc2LpTcKYQmRcEAPH0i3Ttjvk0kNx7KvS2MF1rDTuTaPOQMN6c+
hg0FSsC6Pb/IgHhct+N3ybpJQZuK6la6DMkq75dVOepsT7CL6zprv/7D8/DCd+lyvIts5gQYeBg6
Jf6U+jUcDqGdZ6ifbEnq4UnR6lbk4kvS2v5JQxpdjOZ15TOCfVrxI29HuDd7m2tdCo5FdekNyVxK
x9S3/oR887IBhrKNNyt0OUZaQYFbES/H9toMorjR2QpOnqjit/s7BH31xDPFoynshdOUZaiRlxX5
MVUelxWUjWsJzpgHdkGXkFcExHuSFYprwMJLRaMkWsfUjvcgM4MWvfnj87nq7L/qI+zrk84O4/0J
4jYXa741Ycz69lJVXB3emrL0miUcToHjehjL6K+5Nwpc4FF+MWCXOb1gvJMjyWdzXy5WgRrb/aBA
wUM6jG4NZK8vM61gYZgRa4pzu/sI5eXdy8eeToezAob7CGixm4z5EI1mdZJU4obeK1uBZoxKz+XE
XMEsZwx2tMNSyEffomeTmhfZ+7/v1hpMd5oiceLNmfZFJHLOMN4oF8q/0zhUnmM0AQB4/X8WtShG
sPfJYgC560nwt/qcXZK1oNLtNN/yUHmv+7e7aaFRVEb1qlJqPzNcnWgwXRTK+IEhYOoGRZEbhqwF
iw0kViX3s8E+v1tpG7xJqqpxIC/cbJs0rfqeqm6xQPg0nMMEB253D1nEvB49BMuZT++5klJxNpM5
leZb/88VirWEtxHOo8ccqHuKL6ge2Ds6Qt1uLJycOUjgQZs3A/HcZewaR1/3jg22ufm3wMfZWE1O
WeXtyMY+6F2mZD5GLhZdoouW2QMoWj49qDf6gyzbrE2jj4UFfITvzG5siOI3neI/Uw1wJHLX6WYj
HCRsorNoJmd/NgVqGMlvVGQ7ydZg9Km9DJwBmsXzHi9jZaZY7vEldHDZ7Rd1sxZZLo//bdR8VNZf
o1nPO2Td4yKFzftJqHN9AZ2rVwfsaKKIqdMSWUPJl0WwspuiKKgo7eknH6fUncScgJxrX8BnN7VO
s4S1wMSGECM6Z4wuc0Xw8LNskhn3WXffsC2hpPvQCqKVBvVW3SNuayXhwfe1UBB8dnpShHq4kakG
rWEGafocaXOfnkuew5SgK4SuTUxH0BCW0BUC2Om4jhlTOxr/vfIbIyK8pZgcxQN+47Rkyh5OmQ2t
FUviwaG1moLAhsrylgc0gF3y0zkswfV4B5L+7mk4xz7UY1i3vGIrj5XYcPbJmBBeb5EB793EAdF6
F021P0KGt0nI/FmU+K7mPfDv5uBoMWnNGOXQDrIYVt6IGb7izGi0/gHSn69BALb/0v9FA8J68u+p
SyPHsApd3YgeUqH2o5ummktzD5iisrVbPwbAgi1obNNKOtSJFbQOxO0aX/k4wdtykTHo+RhcSP6i
s4vTC9dElTu/wJjQAQGFuOxraoMkZBASy+Om/hNgLYG70k69bMuiX0TVwhRMuUMuxoCkD68Faa3q
wYpiGigL6w7Pd+ms6nMrMRRnTqFWOcKS7qCLn1hjARKn+kEuiTBrNfiA4EjkApKdPiDdtl06cNwO
dJsdfndDHzSMbphEJMfnDJ1+a7myFtOFN9DNAxkVlxhMPPm9+zZ9SKEJNftXuZGn/mM7td8aajPk
LHkEa7zu8UDJKg1Lag8YXC0PVNWcVVLUTnMdQkFIXynAqCgokCGRqy4QkUourP80XC4TAerQ6l9m
LoPBsscTBNW/InJk5nvNAOpTGZICW+duYP6pgNk1/LgF1kNkn8RCxK6rrmbdRHxmKigEO989ehRC
lXtKbMQwNBg1FjejOTIjNRdNpuUFysQYS4wgNrGQtvXvudYsAi+yFDnxeoeJZbzaP6YNfgZA0LhN
nTBA+OpxTkRbKJOp+H8IjoeSqm64Fo63HLy0z8231oEr74ovLuWyTfnJa3mMMREj2FAlY4h3wckW
8xBixdr3JC/F4Y8YD12iPImDoUeqdgZ3AxGC6/y7cpyYjXo8liQtsF6erdGeGXM/QSUAnNWMG5i3
/IJdGy3UDkKGWiVGI2pCTsssbsWUMnuaLPYjflyvnDa1IkmhE6KjIcIN3uhYveIdXhJDUgaB3OHe
L4osV9vJ9loj0aansWlcuUFrvGOeGulLqlmV6JwMpS4sbXpgxwRLrkKodjluBuhk9ml9ebZjgvvk
nCYfVg+5X8QBEMmVHKJ6m9Udf2m3wGrqWcw76c8bGKXr4x87tgAkz+LAo9F4bdbvXyQMk8PixCoW
+Z5alOew3djNdSfXknyyCY0idAxo9h22jFZdKXQt9Q3++Ind84FP9pE9khwTZrThblW2Oet6TZ2r
qIr/B26XrUryQQHRQnXSO6qDAVRowJyT2LjBTs5jIhpOuyutiaB0iXmMmp0Ozryk1Q1qhsvhgwtu
M9HB/IY7XqhcfpT5SORF2mFsi435yCUI2x3UxerTmD9CPhDhyxOnhyhGm6im/BzwK85uRdaELtN9
/0a61VIf+/3K9Hfvnr1c8lZg7Zez0cwTYk5qrKNveItphSziOTNC5dsfcLUE0eTmxGKK6+HHaWo8
4nmWjHRny/gdLWDA5pA+DM6c6OjTnoMq6JTDEa4OVQM3jY9T6fehyT4MgD1osLkKXLO84pVWZav1
eNzvLwCydGKQf3VJRXzWWBezpDzn5EsTrAlp3RrNgN+HaoppJ6g9JSZd2JMKJVfJ5AX94jlJ4PPF
sFwrHxADgWxZFoh4nUXLhFqRiOfjhfMoYVLMKpKpqyQiV3zngqabGd4kjfPcioPsgV73VIkFWZdl
vlmzM/K72d64qD0R4Rm0P3ZD4HXMGZ7anvhvN0gyp09PkZwEykzVQN15IgeP5QZ9q0PXvNnjuy7d
rTfEMTAgR+rgyRTwsu7KJUqtwH/nWG+3y0d9a0F3QVuKyCjnendUA1n8Ds/m5ynAjNhl7y/V2hDe
YEX2VeJ63hjvCRzxRtY3x/9aK0JEDt6NszB++oTNDfo7wBmzYhKd5ms+CgOHKTJJCNU4i59dyk0z
JFY72/hbf+haeItriXmMImnXJB9UtC/G4pIjl7eX7CRTCVY4OnJLkebwsA1MUE2oSjty466v/and
Y0DfnzyeZ3FhXdPSWuEQMc7qL5HhFxGwXiVGN1HLDi4WTh6ij+imUeRBIO67TSYwWL7Ax3VszfnN
5TWOnl0ZAh8BC9ixbMfwLHPe6tWcBWDeeSBmWT1exUFO9bGEaPqti/jVZ0ViqvVivk0D+wI1LCzz
6QgyD9cQ7m2jCSWGrkvY6X71RN80lAVrdxMXMxaghS9O2Szothqow1fgT6p5Mj9+AGs9aQhoTEUi
RCL1i3x4eSqXYKjZhP6Sr2kH1kkU2icPlBFnRomay1H8R1Hxnx0EQiW2D9E7Ra+voOPZNXc8Jy2w
TLnb2co2dKIJeLFppsYHi4cyF0I/3R2TX7HvEIffYkZluVBqQuEBkvHS/9KJbaDmeDw9oF73z3K7
kPOgwbrLIxoz5D0Fg0Lo+7ERJtWGW7BfId3gU4J15gETKvoj1LspQYR94srFcHFwmZqGiOZkzFg3
3svy9rrGNS7Ub0fZ6LxeWaw9kfdIRjFrrVu98Q3AfSPNFcxCRXZI+A/FD6reIo7F/Na0yQiOW0yl
+cflTjH1mUvmdd0XIKK5xMI3zve+ZDQYIEP5KSnEll0CJTJUIaYay//tiTRS3yZAo32g2akaYcYM
aRAFn7n/yiA2DOR7rT9oELMjc135dgZadiI5Ihz8EsUDRY5datI9kkUsmBHxBmACrgbcuLHxqR3y
/zynzNXvlvAWtI0ZUkrLUn7mmQxmPn5gUA/HeiZ6Tka2kTBNNjcnsxlE6MksZtqMaErPUgwPtnQE
76AqBW8VDz36cnG4yo9CBbhF7L2n9HETX5tn+1NwcOj0FUofeRNrrgT9i+BEDx3VrUPZGTGefuHC
lrdLTxIcXJEAesuGts6obE41ZPR4zIKFIF96baRL3lTtdghXKCVh+RV3Jwdr/7y8rkyYqPSRRBIs
jpfEqGEW3rLaZcf5CIrmG8ShwVBsNB953ROwwkmwZzE4NmjMIFa6awQhJdaCvpMuq1tmc8rOpDRY
dWLhLO5aBBY0gvTXPuHl4sN7wcTSASR0TwJW/MTygrdOMZ98pRdGU7SPhcLMV13O5EsaUF0aJAP8
gXWNxBIQGUW4Iaut4xhoHjlfkr49Z2sMeW5TrGUyI4CXEQ5zTOMDPecNMtCj++nir/syEUgPJi3M
CnvyUB0InJq0ny1wlKT1sreHxTk//YtL99nbegIdaUHcG243gnenCJQZEFrF9MuvRPY7OxHOcRux
Nv+Ntktq8wUIg5QSfT/3PG10SWxuTk5O7npDIVrx6wLmwOpmEzNRjmaNeFbQvIeT0Rx7t7MrZ7gc
xoNgBpRkYndxTU7GPGEONRMtJjtyGssVFgNm4qVhXoHGhGeMPjw28AUIPpSV6iCf7ryQuxgiiImJ
y0ABEEjuPSlysQVL44JSUokVeqOKfBbhg0kcHf/izqFz3JpzUGWwPoHmz1pOBY4q3tY1HbIwPA3t
WdzBZHahmjDDktoVNdhwlZCFFT5lobAypcZ70EwQ1lztwM/0BYyty++X6riEGb4MpJkNO2r1pjfp
WjOvQZgRIOZ/yQVEHxvdUR/yaTxg2dkpBeL2OGwB0Tfk6xC6mGoydEy2JFELS3azUvsRU83F3qWt
mZffM8S71W4INvLbnovfD2I8KGPiIQ19iEg3NlYimjNDOY2ifKVfBfsTu7a4sW9WRAkY0GPQIM/7
cp7ehLPErUzSVnwx2Htqeh/kJaX7WgcNpmjcJvH0O5jlSh1CZT7ZL+XlMm6SAddmvoIAow7eXzpZ
u0bFNHW3Xlr074yntHEW7vMYkNL0/M1U8Kb9hshqtxeInuEHUKNFRHZZnyJTg7sEARak7ghpqaTP
tJrKxjmSDfWfC6dpVpod+WGfFYhdKtOhpj8sdEoP/gEO3UJahKT/9Q0a2qTEVm+2hB4gqGlxNeWy
ixxR2WyvsSopnxbzU8HtddEpYLVr7q4RFbvFLkyRz1/GVhW10HAnyoZeH/UxDCXgTzjbTH7CyKYK
07u6DNQzufegZ5mm9YpJB1ZNoK65FddXMIWkv3BMM0SbIVeCMj7JiMDQ5SceLrBWivU7jawjoyEk
jGrYJ1UlQYy4eF2dUWBQZa9avK+YdCPUHdqgcWmLAyp5UXG4Kc+cNl9PQsxUA1055ddNZN/UBm0f
tgxoXD4CDofck2/G5fAgyBpUMBows2G9AT2mRUp7yoqrcgLcI3I0EtZjqli5s3UlZFDmcoag9n9y
vbPLDfIMUuFOzZVQErT6OUYa0H5rBHH7lyefwGcJROfKl97wfYk5JG9llqf/qfRMSXl6tT6vLtFi
qX47T7kNJTaTZzeZUtmQsRAmPl91J2P76HJF5aZng6PGAmSI/T7bwsLGcXYVY8+SRWyzrM9ecq86
n/RheIYB69m+553C0j8azFPQLQN6CyQlk7geSVhvSHa2vYsd22ftAbM0yD3EIqvTdNkCcPipK9+k
I+yWBe5/4wPFRdpMXZwbGHO0i80XPTcMmIXPs8RDovTT5LWfCpLTykm4oxEHYiGxntatQkbIhWuy
MtlOgzuUzk5DKuI3SW+Id50Rak4wS1buyZ1bI7/KBdYx4CoYZWm7BysD7wSW3RUf5yJ1mec9hbLm
q+s9ft/gsbjyApZUswoeSz9xfmodnh3oP1Ng73YIc574ybZdqMNi4rhx2UF1aXioqGKTW2l8jdyd
JAXnheoGcrcD482OmTs+cnv/mz8pKTOEl+04AIPTblTFrv8xGaAwYMG1t7IPpjlPEIMfdI2XEFrk
JthjD5HwV8LQEx/d/n0uOuU5FmDGpOlTjtVpg+JeBeL6S2dlF4On2HOcFENPQ62/mpHE67Tvh+74
85e6jKAGwYdeMmdTNlKHkk9RDZn7uyZOZ2gzeyHBNZZDwQMsFTqKGBJjtJGGF+ie0Ld2UplCXDOu
jW1La0tUAkO5MuQzFVFunWE4rL1vvZPYo9owhl6QPwvKGsLQTYTvjcR0AkdhOf6ebmaeGLBhd12i
G1F/0fitOG4JJp+EI1tS8G5PQtJbpe8gbVJJGYZRabH1bYzrHN64yDBxqZNGMhKQ8qUne3FZuybj
XztimYs95C2ZZe2MbZGaOK7PEYUqCUokE3g3R1aeBIMhw9B5Ofo7gmBjmMZmanqOtyt1xSZGfoKw
nBtFM33jVNQNov1tqabdE+GEMLpKxOniD8tNhg1zJhDqDuRm99/MUjpvWs6hX/vskHtNc8KyEnpu
sEs1zfZwCRIn7XUWKiEtf0nEH3S+jXweW9rrLVsDyGWtHI6DG73coIOmtuVWrWwLFq6PPGuCku3n
uG9BbI06aRENm+RizO4IEBVxDrnnS6Dre/e3FujVgbcwCr7M/uP9WIOArXMFFhMu1rZkYpm1g7SN
l7j8y2+qdDD4zuJB9OvbeGzRKmgWjkV9z6qkSKGOypKR5EtB15FmhxpoAO6LUCEwa0Pg/4k+XcSj
bY0wjrpHqKvjJrODQbsFHtFDNIsMxk6Od+y/LFMoW3x1MEG7dy9e9YYI23dvdKXkwK+lgBryNbQX
bt6zNbafg5u6VEVv+DI3hkGIgAfhPfecGpIUk0fIBMJwXAJSJX1Yc0qGy5FUfSZyxJhjtO6QKQXL
fKf0ypZREFmQhE00sp5AwaOceM+kIh/TgcNnr2rlRAoNxkZcKkMGLb0lZPKKw6CdfrWZSfCsZCUl
HkMnopXNtp6TRzpY1A+OpWOcZtsdIu5OhRfBroaRa8PNgWoJV2W5TRGvXSgbSYowckrQIDeaOd6K
3syGNKjtExrJvL1NhQrP8GFGlYp6tg8kOjF234akcla+oK/GmzaSBOqzfLatbhC5VHijOYj30ivg
SF4lK3rd89LTSUVKuI112FAbJWScvVtkQm8CGnKgRy+7mayP33Jcb6C1svAYF1OjjL8F/oJIPd/W
3BzayJCb9/ycXP6CX2BxJ1GNQetJaE9Y9fIwa717CpdjC2lL3+cSTadSyhf4sTU7T0LwIxHCrc+G
vE7p2wF5HRIiQ3D6KCBODlhTfvF8Ra/NyMgTgnnPda285HN398sGWJlV55b2oadrPmpuo9Lfk3+b
r5w4d9bj1gNFPVw0fdnClwO4RXY3nXPQ7mW7Pnqxg5qNQiHeeBBdt2S5Tb9jdtWxyEZm32CvQZdl
yCs2JKpqW4XU+GryrYj8oZM0Fc5iCo/SSYLY4sy+FasSO5fWwp+ClD3UeXXLzuSC4biY05LacHXf
OYDYj+ZteqVRkVGcRu1WzbrTgTz/Hs1m6KU02+/4NkfaSCSepv/cez+VR8fcnV6ogXuS2rBeXegf
WUeGKWJEvO0VAftcZ4ESERZZ7SN+mjdr/nojo8BIMLLz5PSiamJBo/DsFU8FQI73C/M7ZH+CRVqx
6HxpIpVMqRk2/+JOmMOIaeqwISyqGvj184xkoVSdiWLBThpuF6Oa2EPRMTYbmAQtGgChbDcRiYh1
racMIPTG7Eo5GMBViQZ9EMVS2mv1utJJVkuesO4E9Tc74sLF6fpyhKd3NAyXebfD3pB9bH0ZNXb3
m1CD8X6EfPN1WysMoTzoBidan9wHJPQffV+1clIC1F3e2oXVWBem/uZI+o+n8Tt+q2g2GRqtn96Z
Awk956A0MbJub23ZzFnXEfJ7lkv5LniEvgQWQFVQmNUGnUz2ZqJ7+jxH2BJ1WXdSDOBfT+ahqP0c
oVnh2fIfQFXBaf3N/v8ZfzMDnSzzzU9yHGt7bjeIiycz6Djt0yx+cU42t21c2lyWQeQA2c7XLnbJ
9KgBczD/f9r+1DDYKuuDVJJix1VFo/CVm2ZxLG7z+yXRZe7IywAjR44j7Uvo+jrXQW4QgALJo8UQ
ClaTeAQRVeSWWYvx+tgS7vGl8BOdNArMwz91nB/Pq3gWu/4L306hGSpcxw5tvjIaR3caGZ15PFNr
BYoBnGepq3wQtyKO36chN27BzdcSw9bmNLGuWKPllpwvu0TBVyG681lLErxLigoM7wZwrXl/0rbC
76hS/mOYv5oVnjEFcLZtL/Aq7NQD6qdj8O/BhJjg7zqQ86W4imSW09wXMCFFZ4wfoU3I5qs27wsg
4v6YtLag8MHSN3HOEYLnrx+fVieZYrjWiIdQ+MzRPsXO8YyzVxOTCobPIEgiMR2QuhPdNqqG5NTp
njdXM/ml/f5DhMrKG34/7XsBFC6ra98cdS/9Rsu70mXMA5Fzd+UcE7HdlfbvuH/obtcy5vZhN9tH
4fWHpPi9yN5/e8tNCoOY6/L1UyvKhOMWl4UnukiDiD4q4Ycjh3bxOjxU2ybaWAfvWITgN3vFUz3E
0cmThrKvUitjFJDnULU2V5Zw/J/MAE9yuAoH2H8dhZTp54+WMRRIubRjf7Wwk6GIhmCvR/qIZ8YG
rA8j/uXBCcNV1RVCGuWOdtmSHuaiTi/OzmQcgimYAT8ehDTRzCRJCNc9MdW+rUJefCmTHtrqJTir
kRVxIoFBVJZzS4FV+Oc/IxhOATggPW+gIZWNnZbYzdPznAwXy2Dw0dvDH+84+yRlLz59ONP2RmKR
CUK0ksVGqEc6+4dcNffdVaNZGHN+JnBADK+rgaJ4yAp+XCwtOKrD0rZjBXvK8FUxi3L4rPXjoMHp
/tBkgLqasEymnCCstCOIaWjPpxe0vFd9pVQTPtIj9MKiSERTjlsr3dK6MRf0L+GbDfl3bTsF7S5z
TaBHa03KANa93PC/iwmssLwPEEAfWxUKPbd6S8bfS0FBCyJWcFFmaPkx40Obfyg8ETgfXO/kSS0v
REvO99jz2MxqDOY+K6xNNBVqh6k89tIz52FLmIuIUV+4ivx7fVs3dSSfVmUQbaSVg3mKGgaadqO6
JVy+0VXBO+OcgT0UG/K/Wg5Zog8Wa1Xfy8t9aDnO9rItk4abL/Izjxd9DEX/pSIsmnS5ib2QinYi
PE75EBBgIy2BPzKFnxc11vVbD8b88m4jvRXWoPQj/peAqjjxicGG2gA26miUK1pDMtjDlejnl7Ep
Q4SM/t+9kd6sW9awi+jwDNLestIGBbFpq2ai5ggVc+BcR8++xVzPXP/pFFYwYGydx/CxDO2x/uoE
GY5sEp++kD9+A9Cmv4NP+k8fM30RFmentmkPSfy9bfROAoJlD6iAN232TPsBE28yQhUITMkBH5aX
33oiSiJSuHJKe13Z9OkdY4b38TwHgC3DAsgt5FcwEeMGx7V/fpSG4QlXUgEDS41mB6H9JpsepMur
cDhTsInzBKjIn6UoeMQ+Vp7l6NSsYJ0Hdb3f87YtHYIHBlTO01NMvNPcdLxr7ENuLU7lUU6eI334
w2c1ZM8Z5qwX4m9Lm9LBChB/ETlw5Sq0XYmYcRI6zFn09RuKrqp3hSVEV6MnzlPb7/JUfWWYIoOs
RP/t+sO9DRhkx+FkvoN9n9+SLykF9TOb+pLJbuQIYLiItvhuaCOFr53+SPHt8k5zWJqW4pfNWzAk
Ao8jL+SV5Zz/6Bb0jzXO3M7su73bxlmoGmDGSChSorSCWjiqG6/xXpJ6rB5MgcX4NtK0TpU7jWLZ
MSNR8YER+6yYvHsQ/jD85jze9Vo6YxS+Gl5svqKJb7MbUp0WnZu79v3Jn3Avhpv7OBWYvDC7AGTu
S1C80keQ8do9/jxXXx/Kh7mzhGbdikc0KM7PqDEWaUBYNh5xyjhzvcgR2aFE9pfeTidCRUdA4hbl
ZGXiTFriGPvvc8sSpQWCq3mQ7lIvgZk1PC2ZL74SkKiOVqzrGfK4Y3CtUnHkJ0ps+9IJVbpKJ9GM
ItuQBmZx8BK/va1dFoyBYFGsYK6IYgpIwtP3meENBdWF3ysA4jiTPYhsOhEnjkzyUhEZSFtpEd8q
v2mvPpafHCqj5PrFXfbBBymPG9NuCM961UpLMdoJ/My2VU60kOkQUfiQYw0EwqfLQxhGcvIahY3y
NiqSVObO3npqAiKYnClSqRNK1GFgAsoMx4ncS/LP+umfscg6O8Mt3NqOXTGwgOGGSkq/fWtLkSJs
r8jVc9CUZXTGRqBrkmPX3DUsxjQaFhaa2Bu0LgwOL5zHMn56vMgrN//gUeoP4b9haWParia5nEs9
S+j+/92GWdRQAsLSWq46+DU/u5WbHtU2ZMBWAcNyC5JMHhKzRm8uVWtZXLtmJDOonGQ4PyJe9idn
WNZHCTcdiljm7uLyZk6ZSHmarrpfKwXmhNf05qE8Tzeox3/ts4DYB8sIhzNH6nH6fTcekv+p9wx7
UphOqL6db3tISFva9IMQFr3fpOItvZj+4IoiI+4ZZfR4my8xd+HHJ0TNaLhR7rMbWM64k2DlSJzw
Kv6MbLnANqI1ffWjS7cX5lFUg69i2h2WuD1/b8Hmk+7NgqsaGkYP4woV+f9jXeigyyEs8rmM9hjn
6mImPnCUQ+6fO33Re3+i5cvv/JyMmOccdoMVUdpyxayP4JsiNgueXfKX33JaHSCM7cIuQmXv614x
gA+LwMgHIoz0rKkN9HNRCM+zNWwvtaD5tbYtkYkZeG3Tnrlp7RQ+jz93dufLqiRwWnk30Mw4oUKe
Z4ozu0oQ6DFMDjaBLIeApFya/Co7xCF9jg9LkOhrLOlytuT/rczQlGJnCI0K/aw0FQsFY+TMDJPw
LcgvJkwyWnL9Fuwt4KCBuMHe16cr117xZsNKyyH38jBOByPDhzjQV4E70yUcY1t53qDng41pqo9c
sU2mnh6UJnZrUgrlev1hCIqMJx2UgzSvOvaN53JgmTn1G/x2IEj1Y76/I/FQ5r9KjIQ5HSoiGTbN
VJutsqukltDzLoWH4kzHUqIvNvLbZMASje7TdXFxHs4bfVGLEjiiw64mTL9+RRLKkaO4yLKUSpOv
kNmIySM4HNL/kh1PO2XJNSleDQERoLxwKm0XTkfN0yHtTBtFWehVgPnJfWukZoCeTwkRTDSoRSOF
KtsEFDrmy22TikX6qRtL2Iga2TmEM2twgrZo5nTRL22N/yowgo0o+QJt5AQwfxH5hsIuu9Hmt2ek
zv8sR9RqHgaTUjTJflj3kHrUUuO1NQny3qeQVRMdsA+egd4GNv62ho260vCfRQzQXkhprihHUKEt
7HW0qYPhXNdylc6t2XakDOGtAz0QCez+14YW0tB1MwnHmCAWWi3YISWnsxdxZ8i24U5GcULmuCe7
w18o0ko4X9jK/+d4LgSeaJk6maszXWMnduk6rbjJJC7wXjpjmhBmg6sou/82UcSHoj05q6MN59FU
UjC5KvBtCCA/e2QIs0BHxBgTHEu2issCA8ce2Ch+sx0/TIL1YkAZRdylPY3EfNPbSJgFgkejDrZF
wzYKn/tdsQ0hZ7WphsruAh1mRNKeQSjOCtx629ahKUtuzhPW+CNG6HnGN8DvVxsvFJDMu8skLDV1
GIPSOCgppoYtnpRPFCIYDIt6vKhUbaSt9RM7KiwJfYzQ+F9XDLAGpzlq4e3codC+Gu1tx6pdHiwf
zvp7Oh+3wJOSzmh3/6SyhSQyWV8qSqqnY8yvyVEt/kP0F4BkFaRO5rGLE/XgTUm6m2zGzRsctRxW
JJ9592IgfBkvXF7m7Mas+f4JFrA+BkizMB9As8ymFsDHxloE+TQAB5F1ulRSIKnBCiKdNihCOSnY
gjvPX10FUbfvhQ3yIrjqNOkWm7IGhB9DycdQ1v9OzIfzEZ60IZcrbYvxlEiGNbBnzvTkeqt8L8Mp
ICAPoiH26PFi/b4Dc+I6+cFVa7wBxNFLLiz0ePulKXV/7x91umODYvY/CEDjMBBmj6T2ePSZ7b4R
TEMcpd5UCsi6RLy0bUtu/PiJdE3e0a7H7Ebr6FpW7hsw9W9jiFruWmws/cC5VwnvfTaYk1sz8NxI
ZL4J4QhSe48pReGQUBuIeRvXBmyOnZOvrmH8psOmfe+6vhWT/AZTu4TLlQq2jStMy3xvuVsIHq6h
r5+yBUFZp1KxN72Lwcl68GvvELHt8pbVv+gZp+Y1nV0HodC854B/jJL7wnHhJk5aZfo6jH/gK+q0
vjjlALrXuw/k/ViZnithPYVtwfN8lddgA4YxId9Tf7mkiu6o78YZwKXdD1srpFr4FkBzp7/+NR7N
teMxTwQsdUWfowBKHfSpWIBbfcXYVXeX5Pw4ExCqmYe9w3ustT41AmR/30nI8p0m14IWCXFwxuzY
RSWGM2v9IxiCgXKYi/R98WsXaKISDxr1qoESYrQ554oYiB8j8sGH2yXGHiS+mRBK3NQiQ9HEmhIi
WmYKoTlkcyIL3B0yQvESBNYBUgm0/TkHqFtoTtOCYtXVpJheLqgDOYQ9uU62qR3kZkWIL1A7+7BL
HYULKHok7auMBpqZKzvsAEZk1ElHLNa8YboZJNtyNAn51IoDRvrrwG/4GhCYR3mJtq/WGu/YiN1B
/Kvh7BeVARfKMfIU1uWqlEnndQnwOL+cf+luIae9MHbei91Ftuy5UMZe2vPKyUTPQvvyKHiVtiYd
OkKurr0g3OV+pHl+C9RhT40WGI6qrTefabWI0fk/vcpIZPRwJaymBULe9FuTmYpJGy77F91G8Ucs
uO1IaZyXTcVFRPcvUAc8nMn3EbObMQOSYopyW6fAA9ARZ2OTkVKPcS0NikySO+vyPMU0yvTBx8Wa
/iIDNmahFRtHHYz1ocl/oZPmeubqh3cwgkIdpPnv2+CiUZXGEVoHx6bTHZOxQHX2oZQimWBEOyWS
KF2J2jM04BQVa8N4SdxTKBFhR9W+V9VMQ+Pd5Klp7a4pAXf50Dyor3FEHHOdVTMnCnhfXRTbcy43
qRFWFFtSppb9Pn67GXfzuqELvFpbemYKdLEpV+Lc+NqIfRQZNwqG2m1s7DPOfdnW672k+2vRj3Uj
vw2ZTy0JDb8RLT1ujqR2vIoD5ugdkJKXMPp7GFZWQPCNx5aXc3b6G9nuQbZ1iLymZCLQbkozKmkS
r6U9dzEeb3z4XZVNRqsuX+NwHUD4ea/LA+/aSwJhIpflaX5NgHppdfxGGc9vpQFTH8dQ47vMAAey
ebF5lGcSOpEVmjTUCI7mKMEqNy3uo6w46QET/3UUWLz0cKhQ2YyxFOJVyhZ6/7MQIYnz25POG6PJ
HkofDIXejeNC/TVZ5xg0wZnuUbZ7i/EAOjXEEdaRQ1dTPu8+eb+9EW0DBOBsXq75JYROpy6QzJVT
tHX1Y2mXgVvqvZIfGtPbmL2hA2gtq/4VnAJmNj21ITZ8Q26/5KNRdRPNlHfyL5y1tXamwTs5DhXb
ILHC09pRsXcQO3BQP0h4bqFx1xiCIW/AhXXLETV8F14me/fBYxndrS8yGqWGS7IomNznoBUj0fX/
3GD5942rkQ6yN9TLFdtfd63Hmts9Zyq+g7dTM/SUY9btQUIjdjbhq6Fp1sVzD2H6a+1VPFxoGO4A
8fQS3GPcBTZNqsc1OB+a4ccn9EWnw/2odUm2ZxORx/E+3zXiS02ArMhMfIL5y7KNglqdDHwUbK7/
0Ogesj3xjLHZURd4+Ox952jRA5XyvcCYfhaW3uXHA0aQUTZhxFhirX9J9xUfzNNxaGjdPW+p8r3A
VEl7b6/FrClyiLnE6EStRUHdZ5KZzrAm3EYC3fzN6NoDmzZ2tI8OBbJr4mMM6ZrygUvM9Pa4m33o
/YhZn2B3l023UxKG2nRVu6fGRQWNeQaGwdG9XdrD6hqKyAHTMlBQ1YSh4P5yhF/pNlxIxq+d5Zhx
Q2J/4vRCOFkbGUQP5X7aKtTbyXqgKp743P31T+u4WAs97sRcdmfGBPsV7Ml7Yw5drrnvHHOTFrzH
x02TQ6tnIKVK4oyaAGm7HMTcMBwSPrsWfGIXHOWI333ce0Oc5C9OzfKp/+2nXUQafqf5s95pqY/4
sO1SGyuEMED78FTgAzroL4QDhlre3L5lbf5DJQYIQrZFNEnFZ7UhfmatfcnXsq5KFnVceLQOE0fT
tKljcQQ+qAGHW6fCO7NB3Vsx6lmvKQrQOCSI+pp9vuv/WszgTH3dmiJ+sZRxyRMew6qSRT3FsFwL
KKOsqTM8qQbpds09SFiLs5O04WvdTmFnkWoe5149TOlKsc3SKRHiRe2fUN3EpE4xon+m8Fj6rDML
DJaqVuusoIK4BtghhMC5SoWXYKbgLwSFEk9ysYJDCZIgtOO2DfGKeagPhYw+s18EKdxyfaRF6/lW
tqVlQSufSfnx86jypdav5KOddeSomhak11JQ8iBiWUAE06xxIEZPCsfVe4o98KAxmdXBft1m0m5/
ez/tm/N4gUWxHOxAPWAlFAdKqp+cGUADydNF24TUBxm91zei4QwCjjMmocD/zA+ThOOpeCqgpydA
KrPB5SyMmXHs8mZ7Cbv14U6+b71/RLe4kWYMcPx83xbNIumbWA8ZZPbHpPrHoSSts9+DKbN8WaRA
qkCLXathbgtlPMV4PtfI02mBskZX9RpBYUSH2RStgt4UcwOsvkZbMNIjvIjEcOCeF1xA+EXOx+sW
IBOeCkZZ70r3pOqXLjONGsbqOx3R1l92go3f5pWidUHhW4EVgeSbeND0PrWkSjnSjFjIGjkYnCgR
jghTa41GBiUmmyHD16bYCvQlY+h0/0OLrV/JgbE4Nc8Z4DpttbNUH6xKI1ac5dPdJ23HnFSdBoub
3vtP2evCpjs1q+KhGXd9VYSdRUmaSYBMgKA4fCqjLOV6SAIQemqtuMes2Bd6Lgli8vNdU8GIX+eu
/JmzVjTKwF+/LFAEDRsDIo+EIZ4WHyy4ipJCsgoFEQranSOG5VrbnAgjqvn0TD/+NPqMFP3WjIDR
20rn13XfOXd/j68rLD+LLJAww+0CSLSMeEmWXpN48yjB5Of5HMBERsA2ILSz2VscgJCmIrU/DcpP
2Fi7Da+ZQQt5sKzlus7MpeM17s6om096nvwoEbTqZNfk50QS7V4XzcsMfqwWSJj0+WLuXBcfi6+B
cKAYflqauqB+FTtSCC1NH8fxsFzbwijqj86Wx8RFLJ8OLCM=
`pragma protect end_protected
