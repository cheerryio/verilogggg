    .INIT_00(256'h022bfc204e01d003022bfc09c070b002022bfc204532029d022bfc09d0732206),
    .INIT_01(256'h022bfc204e001000022bfc00ce020780022bfc204e0202a6022bfc00cd032206),
    .INIT_02(256'h022bfc2052a20780022bfc205062200a022bfc204e0205a8022bfc00cf02057a),
    .INIT_03(256'h022bfc01c002b04f022bfc205122b80f022bfc205082b40f022bfc2053c2b20f),
    .INIT_04(256'h022bfc204e02d010022bfc11c01010e0022bfc14c002b10f022bfc0d5042b08f),
    .INIT_05(256'h022bfc2054a2f032022bfc2054c01001022bfc250002d010022bfc205060101c),
    .INIT_06(256'h022bfc09c0c20508022bfc2b03c2050c022bfc2b80c2052c022bfc2050820596),
    .INIT_07(256'h022bfc204e020506022bfc09c0c2053a022bfc2b02c20542022bfc204e02200a),
    .INIT_08(256'h022bfc2b00c20526022bfc204e02052a022bfc09c0c20536022bfc2b01c25000),
    .INIT_09(256'h022bfc2500020536022bfc2050625000022bfc204e020508022bfc09c0c20544),
    .INIT_0A(256'h022bfc2055420508022bfc205542054c022bfc2055420536022bfc2055420540),
    .INIT_0B(256'h022bfc2055420528022bfc205542052c022bfc2055420548022bfc2055425000),
    .INIT_0C(256'h022bfc3663820530022bfc1d00025000022bfc0b03220508022bfc250002053a),
    .INIT_0D(256'h022bfc205060300f022bfc2054809001022bfc2054220508022bfc2052a2054a),
    .INIT_0E(256'h022bfc2052620526022bfc2053c25000022bfc2052a20506022bfc25000204df),
    .INIT_0F(256'h022bfc1d00003008022bfc0b03209002022bfc2500020508022bfc2050620530),
    .INIT_10(256'h022bfc2052c204df022bfc205401400e022bfc2052e1400e022bfc366451400e),
    .INIT_11(256'h022bfc2052a01100022bfc2052e010c0022bfc2500025000022bfc2050620506),
    .INIT_12(256'h022bfc2054401d00022bfc2061601e02022bfc2050601f00022bfc2052a207d8),
    .INIT_13(256'h022bfc1410601000022bfc0b11325000022bfc2050820806022bfc2052601c00),
    .INIT_14(256'h022bfc0b00f01e00022bfc1410601f00022bfc14106207d8022bfc1410601103),
    .INIT_15(256'h022bfc204df25000022bfc0b00e20806022bfc204df01c00022bfc0401001d00),
    .INIT_16(256'h022bfc204df01f00022bfc0b00c207d8022bfc204df01100022bfc0b00d010c0),
    .INIT_17(256'h022bfc2050820806022bfc2052601c00022bfc2053c01d01022bfc2050601e00),
    .INIT_18(256'h022bfc14106207d8022bfc0b11301100022bfc204df010a0022bfc0100025000),
    .INIT_19(256'h022bfc204df01c00022bfc0401001d00022bfc0b01201e00022bfc1410601f00),
    .INIT_1A(256'h022bfc204df03f81022bfc0b010207f6022bfc204df25000022bfc0b01120806),
    .INIT_1B(256'h022bfc1dcff05f00022bfc0bc1703c3f022bfc2500003d7c022bfc2050603e3c),
    .INIT_1C(256'h022bfc346b220806022bfc1dcff05c00022bfc0bc1605d02022bfc346ac05e40),
    .INIT_1D(256'h022bfc0bc1803e7f022bfc346ac03fff022bfc1dcff207f6022bfc0bc1925000),
    .INIT_1E(256'h022bfc1dcff05e80022bfc0bc1b05f00022bfc346b203cff022bfc1dcff03dfd),
    .INIT_1F(256'h022bfc346b225000022bfc1dcff20806022bfc0bc1a05c00022bfc346ac05d00),
    .INIT_20(256'h022bfc0bc1c25000022bfc346ac207d8022bfc1dcff01101022bfc0bc1d010c0),
    .INIT_21(256'h022bfc0bd2003dfe022bfc2500003eff022bfc346b203fff022bfc1dcff207f6),
    .INIT_22(256'h022bfc206ac206c4022bfc0bc1725000022bfc3269020806022bfc1dd0003cff),
    .INIT_23(256'h022bfc206be20284022bfc0bc2001100022bfc206b801010022bfc0bc1620280),
    .INIT_24(256'h022bfc0bc1925000022bfc32699207ef022bfc1dd0001010022bfc0bd2101100),
    .INIT_25(256'h022bfc0bc2101100022bfc206b801014022bfc0bc1820280022bfc206ac207ba),
    .INIT_26(256'h022bfc326a2207ef022bfc1dd0001014022bfc0bd2201100022bfc206be20284),
    .INIT_27(256'h022bfc206b801018022bfc0bc1a20280022bfc206ac207c0022bfc0bc1b25000),
    .INIT_28(256'h022bfc1dd0001018022bfc0bd2301100022bfc206be20284022bfc0bc2201100),
    .INIT_29(256'h022bfc0bc1c20280022bfc206ac207ca022bfc0bc1d25000022bfc326ab207ef),
    .INIT_2A(256'h022bfc250000101c022bfc206be20284022bfc0bc2301100022bfc206b80101c),
    .INIT_2B(256'h022bfc204e0207f6022bfc2050825000022bfc2052c207ef022bfc2055201100),
    .INIT_2C(256'h022bfc2054c03cff022bfc2052803dfe022bfc2500003eff022bfc2050803fff),
    .INIT_2D(256'h022bfc2500005c00022bfc2050605d01022bfc204e005e00022bfc2050805f00),
    .INIT_2E(256'h022bfc204e020280022bfc20508206c4022bfc2054c25000022bfc2052820806),
    .INIT_2F(256'h022bfc2055001100022bfc2053c202af022bfc2500001100022bfc2050801010),
    .INIT_30(256'h022bfc25000207ba022bfc2050625000022bfc204e0207ef022bfc2050801010),
    .INIT_31(256'h022bfc2b08e202af022bfc2b1bb01100022bfc2b21a01014022bfc2bec920280),
    .INIT_32(256'h022bfc01c0025000022bfc25000207ef022bfc2007301014022bfc2084901100),
    .INIT_33(256'h022bfc206dd01100022bfc01c1001018022bfc2500020280022bfc206dd207c0),
    .INIT_34(256'h022bfc25000207ef022bfc206dd01018022bfc01c0701100022bfc25000202af),
    .INIT_35(256'h022bfc01c010101c022bfc2500020280022bfc206dd207ca022bfc01c0d25000),
    .INIT_36(256'h022bfc206dd01100022bfc01c040101c022bfc25000202af022bfc206dd01100),
    .INIT_37(256'h022bfc01f001d001022bfc01e000b01e022bfc01d0025000022bfc25000207ef),
    .INIT_38(256'h022bfc207d80b517022bfc011000b416022bfc0108001200022bfc207e136347),
    .INIT_39(256'h022bfc2b00a04210022bfc2b3892f917022bfc250002f816022bfc206ec2085d),
    .INIT_3A(256'h022bfc250002f818022bfc208492085d022bfc2b08e0b519022bfc2b63b0b418),
    .INIT_3B(256'h022bfc2b08e0b51b022bfc2b37b0b41a022bfc2b00a04210022bfc2b2092f919),
    .INIT_3C(256'h022bfc2b64904210022bfc206da2f91b022bfc250002f81a022bfc208492085d),
    .INIT_3D(256'h022bfc208492f81c022bfc2b08e2085d022bfc2b5bb0b51d022bfc2b62a0b41c),
    .INIT_3E(256'h022bfc206c432309022bfc2077a0d202022bfc206c404210022bfc250002f91d),
    .INIT_3F(256'h022bfc2b5bb20631022bfc2b62a20646022bfc2b6492f21e022bfc206da01202),
    .INIT_40(256'h022bfc206c43238c022bfc250001d001022bfc208490b032022bfc2b08e2063e),
    .INIT_41(256'h022bfc206c405020022bfc2077a20565022bfc206c4323b2022bfc2077a1d002),
    .INIT_42(256'h022bfc2b5bb208bf022bfc2b62a2f21e022bfc2b64901204022bfc206da22388),
    .INIT_43(256'h022bfc206c42f115022bfc250002f014022bfc208490b117022bfc2b08e0b016),
    .INIT_44(256'h022bfc206c40b018022bfc2077a344aa022bfc206c41f1ff022bfc2077a1d0ff),
    .INIT_45(256'h022bfc2b6491d0ff022bfc206da2f115022bfc206c42f014022bfc2077a0b119),
    .INIT_46(256'h022bfc208490b11b022bfc2b08e0b01a022bfc2b5bb344aa022bfc2b62a1f1ff),
    .INIT_47(256'h022bfc2b10a1f1ff022bfc2b6491d0ff022bfc206d72f115022bfc250002f014),
    .INIT_48(256'h022bfc2b6c92f014022bfc208490b11d022bfc2b08e0b01c022bfc2bdfb344aa),
    .INIT_49(256'h022bfc20849344aa022bfc2b08e1f1ff022bfc2bebb1d0ff022bfc2b10a2f115),
    .INIT_4A(256'h022bfc207fd0b013022bfc01ccc3633b022bfc206c41d000022bfc250000b032),
    .INIT_4B(256'h022bfc2b64932336022bfc206d71d001022bfc206c432334022bfc2076e1d000),
    .INIT_4C(256'h022bfc208493233a022bfc2b08e1d003022bfc2bdfb32338022bfc2b10a1d002),
    .INIT_4D(256'h022bfc2b08e2233b022bfc2bebb20828022bfc2b10a2233b022bfc2b6c92081e),
    .INIT_4E(256'h022bfc01cd820646022bfc206c42083e022bfc250002233b022bfc2084920833),
    .INIT_4F(256'h022bfc01ccc0b032022bfc206c42063e022bfc2076e2066e022bfc207fd20631),
    .INIT_50(256'h022bfc206d7323b2022bfc206c41d002022bfc2076e3238c022bfc207fd1d001),
    .INIT_51(256'h022bfc2b08e1d008022bfc2bdfb22388022bfc2b10a030df022bfc2b64920565),
    .INIT_52(256'h022bfc2bebb2052a022bfc2b10a20548022bfc2b6c92052a022bfc2084936354),
    .INIT_53(256'h022bfc206c41d001022bfc250000b032022bfc2084920616022bfc2b08e20506),
    .INIT_54(256'h022bfc206c422388022bfc2076e05020022bfc207fd20565022bfc01ce43238c),
    .INIT_55(256'h022bfc206c42054e022bfc2076e20526022bfc207fd36361022bfc01cd81d010),
    .INIT_56(256'h022bfc206c40b032022bfc2076e20616022bfc207fd20506022bfc01ccc20554),
    .INIT_57(256'h022bfc2bdfb05020022bfc2b10a20565022bfc2b6493238c022bfc206d71d001),
    .INIT_58(256'h022bfc2b10a20526022bfc2b6c93636e022bfc208491d020022bfc2b08e22388),
    .INIT_59(256'h022bfc2500020616022bfc2084920506022bfc2b08e20554022bfc2bebb2054e),
    .INIT_5A(256'h022bfc2b08e20565022bfc2b47b3238c022bfc2b22a1d001022bfc2b1c90b032),
    .INIT_5B(256'h022bfc2b22a3637b022bfc2b4891d040022bfc2500022388022bfc20849030df),
    .INIT_5C(256'h022bfc2500020506022bfc2084920554022bfc2b08e2054e022bfc2b57b20526),
    .INIT_5D(256'h022bfc2b08e3238c022bfc2b6bb1d001022bfc2b66a0b032022bfc2b5c920616),
    .INIT_5E(256'h022bfc2b66a1d080022bfc2b6c922388022bfc25000030df022bfc2084920565),
    .INIT_5F(256'h022bfc250002053e022bfc2084920542022bfc2b08e20548022bfc2b7bb3602a),
    .INIT_60(256'h022bfc010801d001022bfc206c40b032022bfc2077a20616022bfc206c420506),
    .INIT_61(256'h022bfc2500022388022bfc206e6030df022bfc207d820565022bfc011013238c),
    .INIT_62(256'h022bfc2076e2200a022bfc207fd2057a022bfc01c0e01008022bfc206c42056e),
    .INIT_63(256'h022bfc206c41d002022bfc250000b002022bfc206cb20294022bfc206c42028b),
    .INIT_64(256'h022bfc206c41d003022bfc2076e0b002022bfc207fd2029d022bfc01c1e32396),
    .INIT_65(256'h022bfc2076e01060022bfc207fd20780022bfc01c0e202a6022bfc206cb32396),
    .INIT_66(256'h022bfc206c42d003022bfc250002f032022bfc206cb01000022bfc206c42056e),
    .INIT_67(256'h022bfc206c42b04f022bfc2076e2b08f022bfc207fd2b20f022bfc01c2e2b40f),
    .INIT_68(256'h022bfc2076e2d010022bfc207fd01020022bfc01c1e2d010022bfc206cb01040),
    .INIT_69(256'h022bfc207fd2d010022bfc01c0e01004022bfc206cb2d010022bfc206c401008),
    .INIT_6A(256'h022bfc250002d010022bfc206cb01080022bfc206c42b10f022bfc2076e2b80f),
    .INIT_6B(256'h022bfc1d0032057a022bfc327b301000022bfc1d0022d010022bfc0b00201010),
    .INIT_6C(256'h022bfc207882d003022bfc327b701002022bfc1d0042200a022bfc327b5205a8),
    .INIT_6D(256'h022bfc2079b36426022bfc227b81d004022bfc2078f0b01e022bfc227b82200a),
    .INIT_6E(256'h022bfc01c0e20473022bfc206c43240a022bfc250000d004022bfc0b00209002),
    .INIT_6F(256'h022bfc25000011b3022bfc206c401e40022bfc2076e01f0a022bfc207fd20499),
    .INIT_70(256'h022bfc2076e2df0a022bfc207fd09d07022bfc01c1a20453022bfc206c40120b),
    .INIT_71(256'h022bfc2076e363cb022bfc207fd1ce10022bfc01c0e2dd08022bfc206c42de09),
    .INIT_72(256'h022bfc01c2611e01022bfc206c4223ce022bfc25000363cb022bfc206c41cf20),
    .INIT_73(256'h022bfc01c1a0b117022bfc206c40b016022bfc2076e223c1022bfc207fd13f00),
    .INIT_74(256'h022bfc01c0e1f1ff022bfc206c41d0ff022bfc2076e2f115022bfc207fd2f014),
    .INIT_75(256'h022bfc250000d0ff022bfc206c401200022bfc2076e2045b022bfc207fd323da),
    .INIT_76(256'h022bfc2d1080b119022bfc2d0080b018022bfc2b4192f220022bfc2b00a14200),
    .INIT_77(256'h022bfc2d1081f1ff022bfc2d0081d0ff022bfc2b2592f115022bfc2b00a2f014),
    .INIT_78(256'h022bfc2dc080d0ff022bfc2b28901200022bfc2b00a2045b022bfc25000323e6),
    .INIT_79(256'h022bfc250000b11b022bfc2df080b01a022bfc2de082f221022bfc2dd0814200),
    .INIT_7A(256'h022bfc09d081f1ff022bfc09c081d0ff022bfc2b2892f115022bfc2b00a2f014),
    .INIT_7B(256'h022bfc2d10a0d0ff022bfc2500001200022bfc09f082045b022bfc09e08323f2),
    .INIT_7C(256'h022bfc2de080b11d022bfc2dd080b01c022bfc2dc082f222022bfc2d00914200),
    .INIT_7D(256'h022bfc2d0091d0ff022bfc2d10a2f115022bfc250002f014022bfc2df0801200),
    .INIT_7E(256'h022bfc09f0801200022bfc09e082045b022bfc09d08323ff022bfc09c081f1ff),
    .INIT_7F(256'h022bfc2d10a2063902d003011022f2230010ff010501420002bff0250000d0ff),
    .INITP_00(256'h4cd4435c52d2ffebd354e07857c547f96475f3efebe44e51c8c7c64e594d66e0),
    .INITP_01(256'hc672fff461f46a7ce45d4de0c2d16279de585fd754d95358f87348d85b4755c8),
    .INITP_02(256'hfd71676054f944e44a755779e8e67bf0fbc7fd7159fc6d6ee3757cf46a42e6e9),
    .INITP_03(256'h49c4e9495bf044d574c35de1ddd9e041da71f6f148684aeb5779ede67bc94f79),
    .INITP_04(256'h40e4427a56fd5148f3c17fc8e1cb7bd048e94765c9fbd8fc477f475de74edd79),
    .INITP_05(256'hc57d72e34fefd4e2f5744ce3d9f57f67c6696a5e774868c663c0fdd17c4b4872),
    .INITP_06(256'hea56597c7b6df57b6bf8fae17cf8e9f57b69f8787a7c5ffce6c5e770fb73cbe3),
    .INITP_07(256'he9c0f560e87fee6d6d78e2cdf2fae0e560ed536365e5e5cf53e661f9de5ad649),
    .INITP_08(256'h7be7f475726161c6e76f6573e7f9e5e1eb75f3e071cafb7571766667616b71ef),
    .INITP_09(256'h7becf64ef5fc68607b55e6c873fd6de37064e960c36ef8ff7de6d875db7162e6),
    .INITP_0A(256'h74f27d64eff9ce78e7f9df67f1e949777bffffe8c37a5e62fcf46b70797df95e),
    .INITP_0B(256'hfff8e7d5f64fe5f2627e6d58fb72e4e0f748e16b6fc37df37175efc4ffc3ecf2),
    .INITP_0C(256'h726d52e57ffc6f6d764f6d6afe7446f87dfce7e96347646de171504dccef7beb),
    .INITP_0D(256'hfb746841e76278f3e1547ad17c6b5af35ef2d6eae0e37470d5e5f06868c06264),
    .INITP_0E(256'h615c4cd8ed4069ccfd61fec5e9fb7340e3e3e65264f96efde6d661ed7eccef60),
    .INITP_0F(256'h736c37424763ed4446f47542efe6cfccf2714068675ad1d8fc416df6495bdb72),
