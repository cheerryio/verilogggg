`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2432)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCe5EyyhyRO4fMdI7LRralJ5ETVaHYmgqXXa3gUhMGeR0p7jOU6FgfuUX
y46TbaKqFF1YdGBw9IpNtATopu5ankKVeOD6S278u6/l9lN0Lt4pe5oIOXR65ug2kwIvXvnoGc6U
fREqGDChJUrd5arlN1QXtSRTeDR6fg9eTcEHE18kC5IZ/PRnLnp0m3Ib1cqzRUaF7OPIxfPAhUWx
w1fUfkswH68t9mJFrRnzi91vD+Xv32RcbEDCzgO+GGw0fZuH+bmL4KAQSSxhnozCzpAb9CQp8Nph
BDWukr+r04NjO8pFDU823Ea+dc8yaJ7UsK7JDxdbi/gp2TyLF7DTQRRcWe/XfaHMG61d33ST7KBG
1oHiCL6n8GLF04J274UswGhRLoZsJuZtMMiDBcTAeL8i5UXZaBevhxHZqfgJnZXDXqAcH6dxnbqM
lO/HtqRe3oyG5aTwCEHnRWMKAgM6JopnNJ9P39Mhp7qhqltjv9g98ARnRdDnFuiF9DsOj0oROm3n
LGFgi4rrFVNN6UGiUBDOEZSayKDKe9kBHzlskBbTcGwNubHFV7PQO/np/G5mdDVzVewuqezuLRzz
PmbG0C130UcO5ZmF2xHyAHjlyhkiswc8N+VBxiTB6KyFT1R7YkPJPC/jAyxa2S/+EkzYMbviBkgz
2HgLklZnjNOpLc6u+LEj7W1fe0N/HnZD8K5BrwGT/3GIUUvBz3BWDM0U84VohrHIqkGvTJTfIW2G
R/XogULhjBmXQcKLCRU8bCEZ0PAHiJFF7gSPPRdozJm+a5Y3/8V4w/bozdGi+U2b4oSlmLvqRJCu
osIbeV0d2asT9GTvRuAZ52DQcoitWzsb/L1N9zgmAiJGf12uByy6BJrYeoMltuGTfHj3hVLkiRR+
jIvRaCj44PKeP/l9i9fhMjSMIJFvP9Ns7fOYR5xk2gv6FiB5z3bndUgjeBFLPYoi3SQ+O0itmWZu
ZR81XgJs9SW8TpaCo1uKiHUitTF5pLIAOZaUlCtSSG5jrjz9rQ/FswuDN6nDiJBUEhmXeh37VJT+
U04y+fBLiCpKhq4eVKMLMnra62asYmrn0MZSPOgi+9pks0hIWaBLBYo6r/vyf3S5UgeJc/7g84NM
VYjWWQSvl5EExz2eqdPy+ea8qSeyWbk0H4trpOWg5QA7K7iNas8Pn9pkJ1iDzAobX1kUPV73ZOJL
05disjfXKivhdgxxu2PZN9i5NHm/bqHHV8tVN5FGQ10VqSt/ol/OmAZ71gVm0xFtUk2ZUOzTCxPt
3/2bCJjsF9eDQ5BNhNPwasKGpZM0DsF9IYP+p+9vYAX/caqTrysFzkuWBAkpydX3BcqQQc6BS4vw
/aFHwMl5A2xqo8fqWsbIW/8CIdjognZZJlbH8tW+Zn2ZZtQEM1Qxkyti+UOPIFyfa2WqbEmTlCl2
b+iqdQCMr0abGLIJ2pUIaMtaXmdfevH9QgR9KtQTbS3gXj0HqC1ycH05c3TZk7AzYCO1YfvKD4QH
Qwer25N9LE6G+4PVghINSAJV3dHYPfbAOJP12r1i7wiux0RhfmtcLHo4ZO/jQiSQwye3wdkzzePN
JvXVRNZ1HDx+rd48wdA1scPSU4B54GFsXyWzbOLDi2MBCq3R4SXRzJTauNtEFPS6wrGgjJTf/ThJ
pxBgUzAk+5CExzvjQUm7twtEjgPxQKvN3fIO3yHYNhj2iNdkiYSUlT6Ao7Onhb9H9MC6JUZub7Wd
sEXNRU8lL/zuVIynQg9/8+5Ogd574+SOGHrCrnndA3lB/El8e2w2F2v2YLvdifFPAYnYOLDFMw/e
qzHRikX9805eO7fs3ERyscij9YSlw0Vhpujzu2FIa4UNPRDssSxDVgDWbV/WhdEwhZ66q3T8xO73
6SzPz5/dARmaZbADi7VFmXmjWzbJNi1YbnVsozF6th0VremUlDw9q0Bxb0U2WLGpMH9DFAGiDHdH
VRxNSTYLcNrl5hqsp8iq3LqGpY4QAO9s7JiGM/TdX2sdFTMsedePgJU5f9OCgGdD3GYPtWQwSC7W
29IOvkTDBVprkobEzf/mCjq21qg37XSJYoPCDKw9Fe1UWLwn5VRsQuIc8URT1wn7EEFAGxZVsFQS
nwNwB45X2a5K9kbVeCtmJ53vN4Q/vteFAVaU3MAnvNlSZryCUlcwelqhS7LJiHoVVPH9/MsbM5vr
fD/nhM4DTMU3sG2EuOvm5nNqt8czRe7E8Fa6IrZ81kYK1i6VVng6ovoDtlBw9hS8p+BWrU+dXmVY
k811yToQcd0uyHSELZgwih9yoAXW/p7R0TONxTAVtGF3NP1lW0eNs5VQBFOT2uZaLozH0AkLeRNF
tVOIUrvPfwpXuzveqLBZ5WIOZnidTcif4etbjpxhgMUgEPgrdOBYwd3KDmiUmClN7n4mgGxHID3f
0lnkqcaqP+RihvKXLymfQh4N//ltIfQbPhy24vrBTpXnfIAB4Rlj2PIFWYAqhXlEkumN0u5k1yZB
QTIRtKDOzzoiwRJuqFN6KdG1eGCQhEYo915t9KSa6TyEFC/H2WnClqN/j9fD2pV4/7HSZmnk8D8v
C5a/cXL6GPfVN7LvCJwLJu/yee0016QKBsg8GQvYqanHvoriT1WrgpE/bItQSQGzYR/6TVZMJ2KZ
4vP4+33X66mk7IV7pZAJLO8Z+MYRpMkonadoC/pCibu055XKCpmF/rGBW4eV3SH/SwLLy232C7Hf
4v/DozRaSJfFyDarrDxF9ed6AoZfL8CE1QRH6u4qYA+TqkmHYW1B9VXoRZWlosNiP2fx2CUnBCDV
MD9EIjnHonBWow4Qip17dEmZqVAMxf2I//b5McfL45LrnjA9Ohbc6iHFxGg6aAxWhsy4o0UPK+vK
/sS417CRCW473LCs/NtGQCTDZStiCau3r3E6eSMoepUSzA3rGAUwrlIBW9bKBEkE2dk0Wb5Fm7bM
0worVHdG9Ri4qTpRvybsHwJ2YWmGVbBQKTVWMBntddZnXGwk4DJfvTPseaLtks0bqX//0q/4+Buf
88gKeTA0+O4St5Sw9rTYDx5R88+u1uIxzT3nC+JXeUlD9sqpqMXHfwvdvU26OnACeK5B0uec5ui+
9ORexcy1sFiIb/JHBKnif/n8Pws/ySZ+yG/fY5QcAo0nq1JMJkpnUJg1IPOXtVAn4OMuKsKK+JTj
Fs3cquLDOhVEtstCtgOZLWKXA0WBLUl/3omx1HHVTZtFvSH8jSo=
`pragma protect end_protected
