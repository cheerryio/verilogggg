`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10144)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpITdQgHaMfHKXyzEKgR2sCFu9F4lrKSPEpXn2SjDJTqo3VhqOlz9+WKRz
Kb+5a0Xtqm8DpLqhRwTFDBiuSKhVdnnSEX6SzCyXpFB9EzYuxTpKxrjPQk8Lnr3E4jYviV0//83P
qwsxvZM6WvP7E5BU4juae5RH71Q7qaseORfQeVDimpgdvsWUmusAUnHfSuIFcPmMc+OU08DzlHl5
+WMPTmQDseXrfRZCSvl4aV5HCt555yvfSFjDjT3YjaD9t+ncfLhEiOeQLDYy/mUJgs3WteADLOh9
sIPsgJFqxXLsPzCmTe8BcjJGIdqF2jjAiPVSeWEps4JUETH3erHXPG+pCUqaRq0URsGMsEAg//kz
HdsCe08ASe55SmJy584qx9z38vqM7o1s+FoyjuCHOnKEBzkNPpQeyz8+JWKiN/kRAYFPgfunFpFg
WMeG/EmelJY/dAC3EPow1iphaas6Pemkh2/EOUV52rsJyvUhueQZe4npqwThW0XfpPTiWLLV6X0k
ynATl2RS58roQ9KPYHEF9V+bXOPL7D/LTQFgYD4hJMSlfP80WB3FVKXpj8hEuv70uYJHF5t1Qepy
PZD7JZNi3P2jPJKsGozCTBQSXI+9ig/UYTTL0CICq6z9U+68vKbLqHirTHMpSL4vzf1XAG8yqiPF
mraR7j1BaKGjiUn+1qJppD/pzhdy2c+xpgF0qAdvP0eMx298yF6CnnFQgA1gwoNr6aBMqz/7LWS9
duOuaFjp1eoRNeKvKvmNuEMBEWrmWzegzj0AaZ4CS8Q/fv5GRbr3Hn+xKxyTcTIkcdnurKMTxWk0
q1troXiEMCeFB4dCaeR40S01ee3NXjaE2B1XGkzpEzk39n1CngLtiHlHbwk4CB+NCXYAuRfVyclQ
Sbt7WpoFAdrq/aYsFvlJhNQTGt0JGCSdZAHpsWhJByIy6N8YFZlza2GKlImFajeXB8JoHedznpQ/
jZjd/Ti1Msn/V4u7i7R5yQ2CgV9fZjbTUTWgkxLZ5TiEIrmkadFJ3uGJ1OJ7Y+oghldF8PNdhovS
rTRc4fZs16uQQrAjBOGAxGCseIE9IF/0G7oeg6+6qz1DxYhdG4lKBOo6jo4oaeW20qXVyRTT5/nG
kOfQ0A5aEisHpgV68UcoKD2qAR4Jd9GdQB7q5Ch5ZHBlbXsL/bvHElnIm+kN/uwfr1cqmRDWSLzy
qPB491UBtMoXH1fSWQmaIZHHbrTMUDNSIgLEbcuJifkq/3iZRy5oIev3yz1Igu1rm4r0eCLC2aOB
x5uKjmxj3qFN2IVcjyl79AhZSEvu2LRjPm5Y8zOZeI9LeOSUCy3ehMlpEi44kwnQNC15XrkcbQIo
egdh+DWhHoudNZeCh4oVjm4tNED2O0aU/3Dm7mmeIAGYHpHoVuZbTXAwwMcX58/mDhlpjWjPkeli
q26Yzx5xfwNFNNa6yeZO7T7nDVYTqogeatD6duttf7SLn01EaBH4bKh1QHcS43d6p+nyRAJxWkX2
d9kQxFa63e+LvGOx1fl1j7/HaFR6Htz8Xj5AoEuK1uOXE+laiG8z/mNQHwa0y8UBEgR6+Wc79spa
DLGX7qDJRQBJ1wUcLmzNO+/QfBwNJga79UP/uRVSLCOx8yQ8WRaTOSt4thzm1MwOXbyMUuAjpHVh
21udMdcnLu47HEthSmtN/jmydN8sKtDNepXipfnsgfzD7Nri3WcrP3Q7N8XQ6jfK22Hf9B2Ct00w
ee8zkaIzdAeN2aLt+xzQ33XuzYvy2lrNmj2fy7C1Z+zmYszRqv3fPa1GKBV2uQU4+/UHXJ7BiNWY
2JoFO1e/b0k3scXXhwweXvr83HtRvjO884F1vJpWzHihVU+zsz0Hsukxdzj306UP45z9RWE1Dr2u
9IwZYWiVHYFu9A9LrC8gMJ/Ua9CYUJYB/S1pAAGvb+79fmxqdneb5snGNZTv7vt7RVXH0Mbts1sk
r5L9aE+GSJj/cPCDKtJI1by8ycSBDkcpEpyism/0/YualN4CiPWzFJKrqEQRA9k+W534dEDAnmV1
M6SRuMYx+RU+MyoU91L455/La2OLIZJZauB9QlMeoqO6dsdhGuxxk4btGUKCdjLzhn8CznWbeuGI
NxxjAYcYF5roOnRtYml+SjJpDm4QMU1Nq1ifQhnDfaU24Le0SYxmNFg0VHq3eSLFyz8bpgghM8cz
pAA1+91T950LkLXJbxl1GjF7ajwaeBe+rL3mgfxveTvTnX99XPHZAQlbQOd4w5AdT6aR7I6Quvel
LTT9oPbAzjKJE+4k0p4uNuN9bTPE7IzCvS8wOcLgCJ6CZblaozJ723NX1M8gLYd+NjvgvTxJrF37
fhwLY9AUxgwuGK9VYyuO54WR1HlREsM9vMPm9xZ33SgtHOl0KL8buJr/lGt9zhhj1vznUREVbuPW
hMF7dZIJW7/2dRdBDA0zaiHvLI2SdbPKgiwV0l1DoGtetq1FhHJNUAW7dhOSQlJi5OYPX0Nu0NFo
ZXy0aoN7j/HXpqGiIN6Yh438KPi3pItAXsAI9d0wkyob8dAn0bJzNaxppPy9ppf3cabBQYqyb3t9
yjoku5c8ljIUh2vbdsjB7YRO2dgfkts5juYdlQESYkXj9pg1ob+NdTv/mazrKoJZXLKwdt7tRlPY
Vah/inQVNNAWWMYAKnUdGjQmvpDy7jD5c9bdHWOburv2N6J3vyZGDQRtetIZAWRd2sHl5dw5Kxpt
tfm4tcYqyfmBdmVevPhrspZ/r5pxlgDq9P3V7zNRG01vBhqZgW0Aq7plwAodr8Y9YQGHrxJNOYqV
4JRKymut8NPI565WZpsX1ghFtrW3U0SKdcVp15e4lY2B9Tpy2TGXkv1Bx7xADCNxfVmf48D6ADoC
8pUm18UZKcmgm75nVr/g+WRzwJAhM173vb6RcIrBR8nxsQ/9eluJD/PiHgTGa8t++F23oRDQXAE9
rum/+UjeG9CuaD811QFNYbD/bgvBvyw3vProL8O6U1UQqfxTw5JaPCJFS3lcSZN3Hf7eR4KpoAyo
+8F4GylP4bW0V4J0MjrUOyXXhTb7emgOZ3AWEBu71UPE99y3/iespXFbewSH1jruwuFVXNg3m8S5
bbZ5jpSYhqSIMIj0GYAdSEh6rdvFfKICUadgqZzXmbe7WgtQymMSCMI95AXaOuzUl2IWE04uOPV8
AB7DPiU++jaWmhOIcHCkx/rEDQClAa09GytlCtYDkD1iznQ3geJGTTp05qexfldt0aAGJMEleBXb
MsZwK3428AigixBotg92mH6z8+rPcOgDn1Mth3IKzQ1hMGSrgPClZtMNeezrd+MzwBRUfisMddTx
Zr0Bm5Mj/VUCzGK5DYGojr3UnW56EX8Gua1juyDO3tNthi7L67l88XCXQmO6U8X0P8iXu4rFxLiv
AJ+r91WVNUAvcNFVPFchv/xErkqvVjOVHZXfzYGMSUXl6fuNu1LDM+MK73okHeKQWqeYFCmyhB8T
PzxstRyxSQooI5OZDFOojC4hvlIl33G5mOb3WjNKf1yOY+E1L2VNqVeJ1uP4lt0OXWhCtMcMaWhl
HGMyv/y/POZJbYo7bx4PG43SIvSJqenNa5XSW6Yb8S4pyvhxMu/QExNo/y3rI2QC9slWc2Lilb29
xUWJeQWkW3dBdvRcVyfj3895JQyZSOSyG1ATAQuItHr0FcGQCnBzqi4M7ALR7OEKirQ5QgGSr1zW
xrinFlYwHmL3gxb09zgoEzRMSXtkKyN5cH/agHywRDb/ho8KVxJ8Up4q4YXg+lWxfNWLX3rgxIVG
C3m0+PTk1409gRKJgRlgd8YrqWH0vSzJ+8T33jSX7u0/Krkdb8pDQpyGpmDAjphO0urwX6DKDkEF
QvLz+ZhWvznbfmjTbSNFtAN6ATHQYSat4+Qdl6F3+ahiTO1X+7vTWdFzbvuDus/ZBIsDWCXLtvZu
xBoiAoeMhzJwJ1ia9qzSFjsnwmcaq4ufTQxvhrfGmqalC27BzUIIWHzzcvhYRXSXGsTuwfw6VsX6
Zxf1yDbYQ+DDh/ISDl0CRpCbCNZZoKOfB+V3acOT1ln+hpwvkQEXHeGT/kPNDwwMpgGRsXG8H6Af
r3jkoAVexpIJk9aR2gAif1Nkv2pQWHa/mkVBrK7nYh3iEuzmh/2ZtmhYDFkApJRbx5f43DzRAS/m
8cADTmokYD5UPaVEZSOWEqnIJ2dA1MreOQR6O/sheKfqP1jTjMI4iw7rGzTK8oqQN64ZJXPIAZFD
/rP9L42z4QP1nSshui3Xet8V0hivUZPVns3iQm5NJURpBPiEBx1VcAI5xqvWglRuU7HJlSA5N6Dr
tHkrx1JxJEFOORqAmR8xNLeVXaA3A4STii/cNixYEHz9VHsVT57hYFvYRkd0nOqsgB3r1Sa3B+Bx
UZqx+gp2xmL2/qgu7Hf9Kl0wNZB2uMsJh7/3zN2QAPaLhvcYD6SZXIYEuJQ6TsG28zWCIq8PXwL/
3VYCLJTQb94TrNVqZ1I/ncpzkxqnjRabYYpRxuqAJTry3dTuj9kWVsLZ8v4bOE39ZzeP0JbmwrfO
lRnWxxQmUoWa1StjAiMf8YRX1oq1y2QQ7lxcgX1H311fOrMANg/uOW/YHEdELOn1GozyIufE2lS/
C9D6McSSmLvzSQnzW0IYUHSev/enw6ROYdI0acj70vTE6HsJGo5IkVOpgqb4cL7rGySsE/F0DAVl
6icJSkFEelupqysTgSPbm+gYX3k4A3nMD9ib1jLvzdz1fW0pSQ7my7YWNV0Rgaj9xUOe7OmUjoZ3
0qjSSnq0UqlfZx4Eyl3cAGdCF06U7myKCJmzSO4nRquHU+KmbOoCMulCkA8u221Jd4nAHN3g3L7W
JO1TUS4dUVa9REYR+cYAUne99NH7RzKNcl6R7Y4ZCHX7xlfqWopObAS3ysAsuO/mlXb2F2+TPFzf
beh8j4EeJ79ZHze8UudKrT0AxRpJ5y1iC13yl1BZBVKmZ7UHIuR8+vdniXnrC+ZeOwn5cAM/LLTl
8Th9tOqj9pR2DyR2Wr3pMVUgr7C8729JN1VNRQYmQvs1eZuVxssoQM4RMRpcV6HGhiGehGU6nrjD
m6KwRI9R5q6jZsdKoRvEtkJR2cWOLEKNsXeOrOjkt7rHmh4zsdXdGr18rmEvIbHAwwNA0OvYql5z
G4jB16gWFZJIi/Hx8+NVajWuarZfJzZQk+2PdmY5jRz6SGGCDY/Tee6YgnNYQxV2GwAiTueVTZQu
HaiPWarjayyjYJjPK/65BwuokHynxljpzkMH1Wb57ncV80YbexCXCg+X66sM3lV7UZLY9PxZ4UFY
Unt/Wt1dD6q3MM9L/zJdk2uzQi1kijZRGlqeS8bqBuS7Zd0f36x5cc5yYXZwxdTGAeBrCYQVFEVN
X3/Z7ZkvFl6AbF3SOVtF9bUBz0GlaJMVrz/o2ScMgAQ37XuUysyWLizaLH5H94ekvQcQl0aetYal
1FPAZNhL56vURUaS/RQm7M7hLHt1pF9krlEUYjOsjVbETFwicB25DksvtbrE0hXTZDMmf6RqTOAD
TeslTKPvvdPXg1ttf73j0uYgBwfbzYj81wBld4x3cJwOqoAxnSJ+e1nA5rfuQYlZnEbQ7lL3Fnkr
IAWCrVnmP+TuLjVahcJEkc1QnIVUMraak2xND4+U3jbVw1lyzXC+2hUbgWOlJvzDpW3XmyE78JZ2
GOx3xtmPYXRhZuamGM4qRDvxsEvmqWL6ZOaLii56REhAq8chv0IRXY9gzhMzi8KVHzukZWO2/suv
QsTjEEL9savCZTYsZJ1nyUeT5MocPZM2CgYzvFy8iCpMcXUm/e2uczX5msTlea6ViztVuBdL1rgq
JQZjci//ZnCoFgOxitxCXARDNeXNiM8F6BahzNyB9k6QmcbzVZH1m6E4+UKcfM7WnhHqlF7+PAyX
PD17brnlutzBSLSKN/eMwGN9e8YYZLBmJzmiThenzM+vDQoKU0LJljBQsbPHBTmMotI/TeAByrm+
uAEMBuOfY8Od0Ifqdi5pPW6kP8p2PtMlxSwWA3u+tyuaazX51OQYV3jyeX8jvJ665Mgv15HzONfi
R/0UE+pnDbjRp2izLYrbrov4PBXlBWSZYA6ime7sk01EDV2h26M6ByyUdJjJffa8l6SnOREpfSZS
xdWun0luq2mlclT2lC+74y7GIG8q/W5sC0wbZqD7oiI/+DLvY2bc7amgaRLO9jq2UpxgKhhA7WqO
OrtGE4glqMktiDMU8euk4bFzu1zPBZIng4VSWJypaMLzKbGLt48c9GgpdiccFmyaMzhXgnscm4nS
r54hqt19wqKAavmuw2r0BHoU0fCQ4dFZ2DFisF0KYXQW0F+0BWsdAGoMuWRVfnvsE9nLiIpT1EdJ
IJuHxmCitext+IWK0h1jYN9UM1yRRFeanVXA+aSX0F4F3bkERcME7F/aTiBT7lQnu8XFNoTd69LD
KAE2QtX6hucaoI+XG/VliLrJ2QNfrXbquUIoFe38VdYK9rYo6Wzx23Lt0OUrPAvoUvqY7/z8Hyl4
xu+Zvc4ecgS1aHC2fMwcWeDrV2+zDrsLTArkcwESXbSXJ15hHrCRxFXm5Qv7wuEl2Fr+Pu291PQm
maMxGLroHIareX3pnwN0vPXgltN09XmEYIiMagBryIKRS6Tn8FAhqvtiL66QlVuIsFLXZf+lVy76
9cGKhsZbHl0FxxNN4l6ws7BNgkksMjdvirdhydnIbKcVrhi3BUej2ksTIhHs45BrAjzattmukg6V
wBMvoS6yzRFY4xDcsnXhcW2GsMwB608T+9rxdQeUgN7nGRN+GxHS205WTHgx9OLECUZxRuBR+mRg
7eV0zHI7T2yUejMs7cd0yd2WvJzGljh4rNkDmwH/wy7Bi5Mym9n1zDx59LA539RoZPg0v6HhIrsW
U5utFSgP1cM9UYzg5qLn4SPXeaOS08ZoTj3MfpgWqfY0WzTcDaMgGwTbtWbzuN4BeUGypUvvZFix
Ck7BiljBuZPafTsH4WlBlfZ5Xs25VF6KXgq/hM4DGyCCJkA6dIXx3a+zZv14XaVrz+1b/veYgMaY
PlQf2q5WTJD3evyIMFVwr1zWwnCQ9e6YdyFQZol5jXXad801wtZPqBcmAf7YL8OjyD7q2xIRny4N
OTJbhXJL/kwnG5EHTy+KZ9ubGlTy0FwmCnzwr6aV5NI3myFajaCGM146zvgiozKNOswZiWiVs4pQ
iyUtfzGWuX4akhYwzTYpo5gkXk1rLlxUa+JxlC/bxnhsBO7B2X8Zuvou4BXu0eOZGhFNBD6oM5a1
udPUf+M72vOv7LSdT4SgZ/R2cd97A+w/Y9ub18YQVNMKr19jZ7WdQ2GdfyfjlUytNGNXKhynGBbD
23HWMBGJrK7S9GaZgjr74z/WaT10EZCtB/XbcMMdcSHpVMkbl1Yp47sHSSZhM+1XMchMQoEh/78i
S2FSvozTK8bvvGQQKUF5JMlaMj0X7uTyUj32xbVmotc/XKaOYnPMcskRK7qsQq+nXFNKzvDIMmd1
dwVKr/VqdPGnFJBZDHdcYNYj2o7fFqhqef1vh+QIk7p/AhWG4WuQ1h9rCia3a0XcIn4ZafevU3Y0
njkzo2mn/Cl+lz3S4Vlv1OflQRt0CaNQ5lqqKBo4S4osKwR0zu+xBhWdWx7GU76a10v0x0pUN0QK
yayddAOazUprAsu0Ojt3yr4qohXjbrQXpCMX2Y+PrCa956jDQ5dYW5/lHaOMG4odTzCoM7xw+6r/
cs9NVAKc6pTH2n3Sy4xlHGWS5C+UuHfyuZMZm+T2seJeAJz3l9LdQW4jGiohHJFb77c+Zjb2v+Fq
vARmN41IZWxySIzS4wp1x5sgcue2i82n56HRVXOtSE8EggXJCZVmMd+oeCfvdbKgMPDJS+H7URCn
qME0d3zljJgeHym/Hzn+F6Ki3++LfFfy7kXmI7AhursHOhtEXQKdla4MDMgzMuS6Z2ywJgxn6f48
aPT+RWdVwx8cTNDcE3E5O3gc4jKnVRpGXVabguoIhDPL37FBgnXBssqUExq08dd4NBk1dGT3udEA
SXWEzLpy5mZP+46Kvgn2Fu8OaTRUdeHXrO6Mlrah8FAvsIU1A4M0l9DmIudohk3LqpgPpbzSmmXv
jTm7uqh3rJ/2cgxxJxeL3aYoArna9d0mp3DRtsAoMPq7Xsmfs4FE5n0s6iFQBqW14X5xY2ThrsGQ
QZJVbIh6JouVLGc1QcwH9wyVjDCezdEnF7VJSxLRBgXvWqb+cb+cv6hLFatonqQsW/m4EIiMYEvJ
wPggZEnzUWp7YxJ2PqAIhaL0svaU/nqa1h/UJlp/VcCLlZz0g47jmELFa15veEaiqJ9XpwWga6AG
2oOu6+iO/Ne6/TdRF7x7KcAu/NhQWcGXT2topmzW6q9DeTaJtEN57Qa4xYPlD1XNN05EVE4y1aav
kR+SLXLmlJ8PxQThOt4Ylv0EasBTFnZtJRf/xpb7Abdk9MGl7hy01kZd8y44799qFO4xvb8iDO9P
ZkldRTUeFiawAn0Mm+5IU+gZ5BoQnLytamA1sCrpaTOvZP5FFJfQHow1fjmjFYBoAhtq9sLTNFch
2+vzWBgo0babxjV+MdB/PCyubjiqNdnp3MoeLxF25LjaiXk9Hp+4LW/nQ9yiq5UIi4lp/K8mM7TE
K4fAJ44vcZhKOctl2QfpurTV9mGbFT5DRVHgchp5/JkyJjGK6SITT7gpQdVP6qNCE7FcrMsNbMbW
pXwN1LdmCxE87ewB7hqcNoAbiUPS+7NBl101Gyx5ZQio1+z4zRFCrL8/GEYyY6KjfuSBeqDkNuH1
ymRA+fsSRGbgiuMPNZwuvYlfJq2fMEGRkOCG2y/Lv9gRHTa1sMqN+2CsIO/7g5fpQDMzJrfibFMH
ez0cU/kWJZgZKPok8YT8eFcm+lHH6QUxjwXxxxrYlehoge7vY3c/2hUesxGxYWTQrVr8hd3cZ+JY
27sUm0kG258XcBLrHVghxewJffEOpX5IF1VcfoIk7vi8HJwHa+lSBAy2BQfjCFlr/Vbcfw6/Q6ZB
iOLLtZgzxFM6Vfsq7KdAwcVgwrQNvwsYYWVUmzeOVwyXirf107CrMZ4scqbRVB6HnNbu09K5wa0F
cs6xnWacpsfLsqobt7jP5Qd2/eaJ/fZjA5tgHfcyIf1bSYiTdMlSg5vNzKt2ky+4XvUshul5YxMu
euR3D0it0KNWlOfS+Gve4A+pLn+7fMe9ZU2mQiGNx8p6W3mslwRhEdhcH+8xHXziTS32htg+3UVJ
g5Wmf11xJAcoOLsPdCl5SHFfSS7xCV5maOTKgOUiz23iaCwh2cCmDT9LJ54VOA271s06AvrGJV+7
4fH4pgPHPM1LAyYTJbmOq5YLhhKYdCNHNZBlcn8P8wSFtiR7324lTBPIK9p3obTdfHYs9toKm9FO
5b6T0Ewulvg+RGhDjYXTm77Tl7xBFGvB27ReZQVYdKngiTvV+cdb8Mvs7PxvxxmXxIfkrj6shA5r
CC0PvafvJdrfN3zuJLauAnZ/0Spo+GLpjfLZ6jEHXvyLxuLPVkOFLGPBeRNIPRg6laCNcxsU7cHh
5O7qVutseKvAYRoy9xv/7vXvoCfah1SKcDiYkCNngyQUFumO2SOirbcV6f7gI+QpLt60aXT8Ixyb
RiWyYdLSZjk0+WzdgV19OtRIKSZM9k3aJWX0O1LsQgPqwv1isMKgQbZDS461s17sE+l7OcJ1pLRr
gDsa6kRH00lOAo5HXaHWhSnlojFL6+7bc4UABOb2i70ZYeWr5imRc4KDCTozL2JFOSCX2Di3Hk5E
mxU365D9/O2s0g9pWIfzqVXQO8FGi5lJuE2MOE2rNMlVsQLbLxADloh/IObRsErs4pv157nGD7rh
/gwMxmJv3ZhIFFxr1guaqpoVRdR8GH0kAKeaDeg1USQlKiBvqMK9cJyH5f0vcj/fNVGtFe3rFPo/
7BQzMHsAOJZdLWNfWP+WEeX4Mb+JmfthTxz7v2jRtdGcy0FxXN7353vOF6vRCYv4le1ayyPYH+k3
259XaiCnwcxaTG60+Wn5xWBJWpFdo4sVbaJHvQ0ek5Si7k1FQgiO34JKnNtiTajJvhg25mO7Nezw
o0ouRp05MVF2VI6SF32GhKvsEaa9P7lLNQccdTZcNo/f7ujt0xWg+TdtFJFrJu8FfN7BfvhJpgrV
bKRsEoTaDuZXHCGt44u+bEBC1rsY0AQjo0n/JS+KpjlVgyGZfsziT78UBMeGUpx2icg1IvMl7B1j
SowF6nC8cMHnEfWMBVbnLzK2/ZWwEvJI26bcJVjqGOD0v2WBuZ2Z/W5lkn5YMIoDedvvVlekxIlE
ML+jilqNCyygaXUcECrXp/qCGqyZgfklhkOn7hW5oB53fLogUxL0VRIjHgMRVBpOT0Up9NkUXAjJ
YMimnC3+AsXRRcK7OSlq9249GKcCYX8j/Lwq4TNB2hjFR+I8Kjgud0iV8uatNDA2pJDfwbBIXo7Z
14mlLum5WHVCuOZ1GICWQ7BB0iGxjAu+TVMXiRU+yU3nRKDPc0+kXE0RmZSGZyGBSoyWVTREUiAA
1SsbXXhkodt/tCvARpaj/IpfipiDj1YSNvPyHsj8SXsdOKxhSvsqQb88ue/OQmLeMRYxLA5gTMzg
7C2dgVm1hJTFzHEwMSFlmqyIsV4uA9rkTFmpPW9Meqn5Vzws8CmS2XuIPs9WEcGQGHF5MC2YT5Ms
AX+Lf5i6MdeotQ44Ed1pwm5/J6D6fQpoz2rEaCJp43saNFR+6U6LIQA0wV7BEH+/zFB2cLrQoNMB
egZSXSQPXC4R3CkXfRxDsdha+c+KGu+fNvb0iv/wwahVLg00AYoMK1hRumA7Vds9whUB/78MmjOs
1X6F4aAEZ24gijxNyVTitkeoG+sWnuAs6TpH7JpKaI2PO99FqY2MqvOs9jNEBBW9DX+Skr9wjZDr
T9PKS60FnIRxIi1SmCj05Qpw2AP3G/MNvp1RR7aDRIwQdT9PuImIOAj3mEzKnoz34xXUHyvgAE77
RX7gcjEzxf/HldejhicGhASf4BxL2fuflYsDVr9m3wVJR8jhBffhaq5zvmmLwhq5PzWsX4uHqNtk
zto/gTssN879Ku0UVsLlqMMkVlVHgJj+0jKp8WjpjxjF7mum+K4pRno20BEIsw1mx7SOJG6POGzS
+OZUznWffhUa9oD+G+6dc32n9FHr30VmD4RD75wFzeZRCmrWkAMFY20nYS72c0mSzplRlOe+lqIx
d+DMa3bxMnngCOs+aYX24rRCjbM7qNGksuc8JKj7solOpfwx3Yxe6vDAeAH2ZrBA0tjPJlJ7d9jP
KAkpikAsEWVEeje7FcTXn6rsrAlFYrXJQBz41vVUMwBbgi1tG0Kfir1IvzpYXQLgddWGVXt07gPJ
8KHDv550H3atSIYVMhBxlHaE8a6H3ir2jyTd5sc1fVstFSoTC8mnmtc3WPdIq2uAN1vuHFnL+TB9
YpftIcTE0Em/bKLP5nrqwDdPQTdm727a4iRN+tRP1sDxJ2vSTwEGvfxIX9iuh53IKsCp78MGIn5e
xnPzvpYDkFHGRJ8yDDTww07/oeLF7Yf+4jHDNxq4IwitEdi9Jf+K1+WQ9+czOlcLgqjERY5XYj1J
SCoAC+NlypwHdzIVg6Ey5M0V+ciq139x070jCMHpRzhC+rpJCEI6zjjK6OXEYTIfrOo0tLtMm8/4
adSXXNbHD9Lmv3EgOEv3YlgiwG54lqZO3PGNUi9Ztqf2PyZIS4Y4FWpiEbhRH/pidNzwTbEH12U7
coyaNCQ0zTsE9pykR0YFqslTw1gx1UA6ufMv1nPwVE9Jh7cygFxrbqpDvvDvE2SQFMRR6GnFAvtW
0wUBtZvne3pYgxhCE6vv/KS996craYXlrzZsvuVh7EQThu1rn+pQz137WHy1Ec8jlUtTrnHGKOS4
9nD3xU062EUVWvKKgs9aNzc+eRbDUGWAzcm/pqNRdV4YdTvok1VsXedkCTUMYJJe+isPwHz1OQyi
Atl31PQ+fNJXwIsFzC773TK2yMYZo0YRpeG5k2TZ9Z46PN2T8DUlJLP7oXrUmR3uaR4WZSHWLTSU
79ALNC80ybJ0su75dmYAvfAa4wrICfoCLhDqj3j1z4wFStcjks0GfX6egCcodb/Ip86n+hBZVCc1
jRXGt3R+HYeZisSiOhm5slz1jOTOiIRhjppG8PbvnFnQugEs50YePKUUc8k/VlMigWxm0U0Fr4bk
Ed2xGr25XnOFEIUBbScaSRoF7zSrPINeIVMhYJvqXxHtVLCIw6CH/uqwEnaLyUqNBk94VNW4hjfr
eqnk6jxBqDvlAA94q+n5H0b4wLrLlMxPEvzp3yF6Jak+ioVCi3BnRTRIgD1+864PUWVyavmWQqFL
odyfUoiyQwMVOoY/13+CFYKomD6hwi/hgkJJaT0sLhyhcVSLEnGaw3/kNbh2jOoVGNfv9bu2GOi0
dpx/iciMi1sQrzTuegUpDIhamiDtrbFx5vN9cWxMkMSh9fc1CTJBg9wtpbrCyllbp9aCYIfkaX89
XrcMFweT8xLbu3MNtn1KBqsTjPckQNCY0qOvggDQue1qhtIq2o94vxpu0M9GiWwcWOXJ/x8QxaBT
eYHHwnMcGADPTOR+aM6XkvS2JR2DO7l3issisNmd2xHROnLN8E+SFr/EtAudXVxc/JpWfoEr/U0m
lzHg2Tzq3A86J05wxOMRwdl89ZTS4/s6i43z3sbOKEadwkgUZ6BoWUjSNF/8oFwgJe5iZIEnGPqL
NHRxp4ECIGSnBk2mnT+Q/Xibj9I849zEisZLdsFUem9KpstyP1l+TGYRg55X/Mnu3Z/Lxq3ytT/F
42un7ICrC7BGUyrzmrc5RlPcJL/0l+hQxTLFIkE0HrWoVKUFvd65HYiRb/QDBf8GY+ijluDoztm8
c8VOLC3TzGqIUReu+5ELMlmOTQxLxUKE48jID0+gaj8BZboTamQHXLeax2yhQC0EWPE8WKw/0zcP
DFAnEuLUWAuH7Ukn2fwD65OYNJ+APYbxqXlRFmNu2DxuGaDVzTS1B+sM3HSY7h6K9wRL/YiaIzYQ
BOlnd1lvidHcoK06+3r9G5Eg4+y+2EpIwil8VPwqR/tgjq/8S+6LdbCDNRTgBPpLjeTrefkMT4g0
2gpsqruj4dt1NuQk8XAoQz+HF6LxmKq0/OtcksGaTBcTQ9GcTPoCFCYZmf84NzQzMVTFOyi9bkP7
eNEbaVQbo+Tv6FUis3KrHu6gnl8Tnv/bBptTkx53u1YotZVHh2b/fpZr9uOFautNy+G8tTX3+k2O
r6wnQ/anEZmJNiDP93Hk5+uIu+2ks91Gk3+s4vFSZeI4/vqwRD4H4aIE8xWj3uVimEzHY6RgaNaT
s09ATSIi5Gh4m+VvZPJhFpNBWGFN3aYFaAw0Ic2eTfj7KarU0WreCgT3fS8A1/I3/DDaTxnF1SEH
rQKdYHyM3RWmEG5BEKqMAZGpC0BUYSIu6CSoHfKqCx1Fm6cRZ6X9YugQUDfjpggfLnqRvfBLWg==
`pragma protect end_protected
