`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1568)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpIQNTqQIjsL5XELrUPeApEzjuC0XgnQFFb7CcP6LK5zSGKYsoiJ1rHHtB
8T/WoKjB7ef3FPY8Nh/CijGHO6L2Pxkc3uM7tqr5N9JvgLqD5feK2ZHrqufiKn+7gtx0WXDfrTon
ML7pXKoh7utjGVcQ7uR/RIZ2WUpIRHDrydPRsUu59mL6QuoxOYBWRG7cwdoW89SGDRPjV6k63QzG
4CBu/CRbGZf7yYKBupdh9Xa70rep2AJuhvRoWBv+EzCe2Aur2mDa+uJt4DTR5pRYTfUXMWTwXSJS
0rEn9PZH10Rsjvi1yqSfdQaiJ8qhOyhPHj2KK/1PrSPsDwKXpzZ8eW5LPQA2MNK+TEBWBfYzpqu4
ShFoN6yDw4qrd1eIS1ZnddMnYe1OwApZTOUSX0AoikDnb0ljNLUVncTqz5GvNubgUwMyTxK6vT2m
WIzF2943PJ8vP9LVEhxvBSK4eQU++K9OeTJ+qRwJjTy2MdxBAUSh5cySsSBIWQJbZx/5GDUu3g9M
VXrGE1Fq4QwigMKq90Y0tz9+x1c8WdSvtdGBm4OhHK++64m1kFxkPo2cRL0T9dHuZUlhjp0nXcD0
hjOSaeUM7Iyj/6lZiv0H2h+yjs/6+80TWML2vMl32+KzgF3Zaoob0xRoHq2LvBYLHoTqtjujTuud
Ip9hZQ3PBHT9ofcJdqRC7BusWEpG9oBe/5FINNhRDPanztN8ovMvfUpCv1taYzs229FmU3PdDcSt
COsGUz1KdOXRj8PiKkg7l5IAHtXF4LpvC77HZd6FVYb09ZvivFcQylIlqWYMQa/Qj9dgItbunCL9
Ywc7yRD/JP0zHgpnxbASUER9fcHUzDtzpf/HAt/eiQYNEqpbMT6vpAu0CB2eWG3HpQVkCFvkig7J
OqPhqsvR4nNfYEYrzXaIXBW9fsJGiim8QMKIbC3IIy88gK/GCcxqxTLjA5pKxxv0kWcfTWco3kU3
D9EeVQR8x/tgDxCpSOG9s+U0FhwjgIrWAZGzDMdrCZ5Oeqifji+ZqThGTN+kvhqIwaa+kxxsS7GO
0cGxYLK4A8z3SAhXGJGBNbAZ2t3gkh387F2ndgn4wCe+/sl6rVK5dx+gtPQVwOdIs1KGFqlEYo8O
wp6v6ZQPajf+kp0GCGiW/s/d1OrllfYf0ErW0sva/SF/TZzH1XiiL/nevPnM06ivR9mJfqhKgaiE
P7PjIgeeI6u3X4GXss3pk4aejC88UrkiIsnQPg/qlVn43IgaiYnTOC6/jmp3BhIXiVNls4WTphJH
nN+QK6SJ7DONrz/bcoinU3zg3nzhX0J1ZOzRNO2/ML66dKWpg76D7UPMANOdEiSQ1jMoE/yo7ekP
u1B0zl/bvNN132ZldwF9rjiqbd9y6EKz799ErV+ckOKtcIxzJvqhbgemSrCER8qczO605fX52yXm
ktbRhb8ysGFX323GAZk9GRhmJvwYLQY3xilPXS2fcrjP1OuNCYmAbrSG20kDyM3b/AbVBFNw1q2C
6eppNLiphOdT5avkX8zBR5QG8AtyUeCCo8r0+KngNpTKWU9GreTUwf2l3+VS+dZduIJRdcXi8SrH
r5bxkXdDV8ItyVVBQ18TfXjVNObgJb4FX2UBNJ+mzeDyu40RKQlb3Xaf6+SCDY/ri1XrEOE8vZVf
SWxE1VJvOrPlOyYIZk49/c/9TKsfDZSM+GHN+SLUHjIpbrs/M8Ihz/SJX2FZjj5vNxcPh6Xq2pSZ
bCT+ZAM/s4bcSos8CZShMIaU/BZDPkJDBsd6MY8sPQMtZKNsRspnlL6xXGv/xxWb4Eyk+dsJ4hJ7
eQGJAA8rvv201N75j2VCI0rvuTEsEaMLHAGaDJU0ntqbVZoYjI2rCcNycC94QEZmAKyGYWIkYurE
Z+E3Crgm1Djs9+cYs/ARN18pqqob4X1RNNj8Ofyr5X1CQUdF9LFFr9KqHfGmfhzamw09sX8HHBuC
VatsuX0fGN0cm1I6D+aZndUPyYn4N1/3Z2XJ7ARjVEdQ+2ruUUewtPaqHeys7OcbEZ1eA/DSsO8A
2bydC3nfObm2hgfNo/1MIjgLJdGZViOnFzLAC3w=
`pragma protect end_protected
