`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16736)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpITs1XQmPpnjP+M2PQhx1wDEZBlms4d4yz+GTfY5qh8Zf7n2wQdCYmxD7
lTW5D8DlVmRGQr783/BdyWZH7To+1S6nKq/sublxYH9ix/a3ny60Y7QwWoZSBS+S724ApNR4z3xD
BEjGP3ItzqvW4AL7y87OXqAZCuiu3IjK04Ww2XyPxnmdoPjst/lIYw0vHMotZj2/QgxdCTXUlLrU
UJzPPUxmDpxAZS9ReUY3j6q7/QE44w6yhMlJkfX0dD/DUB/0Q2lz692SBfGvLVFnBBskbB3t3N7N
L2bnSkxlW1cAQWXRCAfy0CnWbA0/SxPWeMGDM6azgC934JG8SoAnxt39RI6VD/XE2461H0RMOn1H
Z7scT+hnjwizSh97tJMm1dmBIygY8oSinTJbas2wB4IGY/5ZT2nAvRearx4iUl/PyqetDAB23gIW
niVcMOBKKaSzZnrK3HNArGL6WlKvb3L2paLK0A3GqKhgLtJN2KOUuAkKFBNB7r19C9hfB0Z9QX89
Z16iHd0W4KR/RTWMR4723gGeZ23lpd6P61KjV8TiWVX7W9SnjxqK/0eXp/z5cP0Ti/YuWIGnH+RA
d4gTjEDmbkpZt2qqPCd4poiU//ZfKGWiisUe1Dj8Xn3tAigvvt/ZIxMBopW48yQkhzKSCSWPJJcM
1e8rToG+XIHMHY1FcJSKSV/CWEloKEed+xex3xQtKVGXp+ZVPNce8t6YdI4v7YzLLB1dZbi2/S7E
fsZ/iioWBFGOjYXp/cg91iW5TGV6QV+njsSL4nZ50V62+tvMORsqo0y1N38RjrsL+Z+Isgl2ckWP
9NA96OBkBsYnyO6H1ybwqIAO77DN2yJXe0ng1TfeDqtMWUHl5xAV9KnlXl8tbz61eN5eEneDKX34
vdvCR/b/20nrr/2oUI9MDItASRg+Q7XCFw5RtXlXu9LM8Oa840JsnuK3VkcMlePturlEe8JqNX0/
BAjlfejiHsEVo04xFFMAlHPhmnzQxO3DuTAZkqyl8yyQoWfgE7QQV+owaUfTS8hkW9EukSugL6Mw
IANkkNeGLtijI8/lFqhrX9hPiccpc9Sk7h3NqC9p8VaILUt5fzYSNVWBvE3UT6yPiKxbfX75V6na
Pw+XryFfv2RTgUqyeVOtPo1vVgCF5Hn+HkKEE2vGJVQPDlmOIe8s2g5vHhEp4fmMEP7IyfeKxBfM
lBoKVcPhJPNUqTZ5uu/YKf7DJ/wXEQZDzAfC5AfNmpMUwrE5K7/qvBlOuRlZ7GiIm64Oi4UIefpt
iaQEvc8bFyX/Cc1DNjAOIupRonz0JvBh/jvso7s2eaPuDwQvHHGt8iZjyHqFGiCaBnlLWPZ0EM1u
rCVITeuvi1odI12/wj1TFS7ULFe0Zus4l9WaU7Tf5eLHqh2oLABD2GXn49xBQDvEV6goY7GdvaLj
GdsMZQKiHbM8xvAsQpaC3AMTezjH4SPhTq8mgGdN11va8UsV1fDrqmuCTY17GpXi//wVsSDCicdS
u1GLU83lVd+S7aOZZOHVFJN6m9wf04jXsI/KvketbrYurGWw97k6WCrkrbJpifOf35QxEYbFS63g
3TcE6YZbbAgf5dRmr4xQrDS0c9KiPTvq7Dk0UONuABvBwIwhdFn/lFDs8vSeIMkJzJbp3B6VldW+
qADbx2lbdpXfMvPX721Z1yuG+KDpE+58RWcHZkcXNsnAc6xftyypKsNO5JgqbAciy7CZMiGTnIRy
OXm4vnqKa+xFPKnqGwvHObowAjJ0ewRjyGpPtHfh3vjCmgiXrKn+XHkmFmQVgUEn909lzcQcF4qD
uFw+rsBGNToymxdmkLwCiOgO5yMLeWT552lrJrK9AbeMZ4iiqRnkxDFzz+GOE1mrasWdeBPann1B
8diAiXL6rxlAruvKTqsmSZ1B2Q9AY59ROqelGVsc61cj6oVfBVyamRvYHydHLGrxywRwHUw3+rtS
TcUNVog4PIrfDjzKnrdPEUHxXDu/GpyZQGMzQaz1vteFr/E1+KnNNRutExkOMrSkfDU3MpBLEwMK
e4WMMRJZJW5bJw6dCo4wFMs0Nwzcr98Fik22uwE9rfh3ysJ6VpoKFXtRWdR24seCLfiUr1Up1mpG
flsBlcGdP+Ww0Xi6p0pkh/9R5MtaHphwFqea9NztvldLT02DSZk23UP3Rp+wRdrkeJXwaD4GuzwV
UX1OvroZ1iZ2GOSY1TZvkpdBFvN8g4NW+PZnu97LfYRNLpbpSREiEZ+/QMVOeqchkzG5IkVEjjKJ
tLohYl1ABgqHAG36Uljvxq9Kf4Ieq/AtNXQKhVj6GZoojZ7FsQAChcE4HqqM4jP3mPf9iNYcfrXF
5Q5ivIiP+C3KpwkET/PfDV1M8+g1kvS+MtvjFQrfkvM/UY4T8K3HDXH9wvSWO1dkLBPPq7q1rfVm
1GPTE6v1mZCkDzm7Owq3EdBdumj9L2RvT/5Om5vt7dneV1Bn6th7A12laFsgv6g3PzY7O+O553gu
VLMcNYDRVZ2lRryYLeSy3uO0KdKGaZio4j5USpdAJwo9Oioc1u3fBrCKPVtJIfTkdF8jt8Aw1JR0
r06/xbX92ASBp2wsHve/JogqDRYtXZfeA96mQ3FS4ia43r1lAK8sxBWz6pMQ/rRwWLzeUfsx4yTL
YnLQhamU0lsrmJ9VmSxH/bbE5Qy/r1vXUUFws38EY8AZxZeJSYL1gFtqkomFPTZjTqBiy5SOYqHt
Yn1f8qGuoB8wd2WKg0RoSePWU9Yd6FgIuYHz2S9M7zDr/HWxM4dM1mibvuenlDi0ZCEBNbYUgKx+
mCfGR0cAG/Izx3cY+aQumQ0hvP+mIj54V/2Py4VSb8BCR0QSuvxYwWvnV9HnyZis1eUUdOKZD9d6
i9fenwJvIuQqJfvf30M+oo5I2GD5gG1H7o58xVrgZ97TpxoOv95JReJM0IF1ZcyslJMpyxON3kYd
kx2tsdAia/jWHPbA/OLx6UWCxrXyq0fqKI4ww/d2HexGpMb/P0Vp/RcLsUTiM9DJqcRAwzGtw0R5
WxS/ZzJbdhzXiTtYmYwTbZyxQkvo6JF6FJpk+TplkbxvTJc+mtnU12vf6eFTxeDBKEKjqAyUVbwN
SLtUdm42xhsPjAoaedEpyIXX0BV3V+iWH5dU4Mxn7rfhVElS5YNWnHLZQMyDI0DKK20wtdzjbfdu
k4JG48ZRKkOk5mK3VMh8GDx79eTNWRcfWcsEhIkWrrXJTgvWrKut8AtshawXkV+eN1AQCHBaobya
PeZkJnlQL3ld6WH/XPzEgkuG/B+t59RrihZ25PtKkdkCQJEbzcBQHDMfQyGBbnLvarfjUA9PF0vH
RtTHzWSWn+ZzfYusFGsH9kdLvv8ro8Uih1VzoJiv1+YCSukKfUbTTQnAqCfS9ta7HM2c6nknSh5s
c/7DuG/NoFIhxNDDRUoFwIjve81UyEjscYtYYabS1IPpYlS8CrpnVjvYY7hyAOELwzfgFflmdcNx
+JiuUnuuzE9yl1SliAxLBYi8EBkFKPu0AU2+2w3JNIGM+OtEYb9Kb6JMCHphjB8wOp/Zz6MIrBIs
4dAic3XxnD0i212T2P30ipYGxvLwZMVIRZ21GG2M2NnYc9dwwnmZAfVnpKB3TrCzPGVDpMFaFl5a
LwEQSpvAZtmuqr2k5if1eJjbJY54h5OpJ+RP3FBCaiz5BdnsEJ76TQhOmFUYPzn+iP/h9gR9n8wb
UDLbA3Hzu5oK+CgZvV3pat5qT6a+Aur5UwgFEipu/jqE/HEdAyzz6x2YKZZxdiZqOTehZ+29hSkY
1gzp5zEhZTu5Th3sZ0kT/y7KNycybWh9jThZ1F5v7yPH62YOnXcyKw26WyfQrcW6ELwGcqoz+K5e
YDMLx+Jehqtji8yEPTEsWYcTpziB4Y6539HQuY1kLqIN+xGS1ab+0w4lF/yyEsd9ZBz0bkbRK4Gh
r5H8nJwp7LzoAtyDOW1zQqAGExno826g4icnAy0pAyVcHJe+NFRM+3Aw9qr7CP0FZ3W0M5JZm9YY
l+lKFxH6n86r0J55GK+e9Ng/ptfDkDTiOYfKwxO21ERrpjUgoAsY3R2alg3w9CRf2/HCDBds8WMt
JC6WQ3m9Meci2kmqecmN1ZFDBAlU9KFd9ZPOvd2X4UWvFFtYUX1qe1y9mT2GyRmr0U2hSfLXH03x
HSXTe9oh/CTXuTNnVm0OXEQtmvz32oZyA02ZeMoxFJ1LVKGTWy+TplSsrpEA6Hg06iGeti6iQcQe
3baE5EATn/2eEloWcn/ZUUCeK/ieTPyTtDlbfXSuPXRftk8+n/xYVLUhUrQV3N49JL0LV5A8NVqi
r3DWJYfX3TAn/XLgTe5uSjd4wcmfF4fzCad+FiuBiPSpNp086oaKt1Z+KbeVQ8lYDYp4lJkXN899
+sPv595HkFymFSCDSw1dP7GnP/2Pvsnh5vcajyyfbrlmp5JQo3RIwXBxfrF8FSHmz2UaKWIjwTA4
cSpw9Jn58axcqKk8WZI3xlnIOG214SLMQ2D35RUYZC8bMfp3wmzTldcl4RdD6hayWrnkABhPinbV
Ypf3DGQlYKszrNrMtPUYYvfTvW8G57EvbgFQuzu6iHVOAIO2Y9NJOYO+qOEGBYVPdYJbvtb2QZwk
OZfWQwQXVHRutoo5gzyHEx9tuELwT0qgIyY+chWF/68kLGyRCAVA4iTIl8BLGvgjsBCmw1c+c2AP
H3iSWhnv20xKWxagJVveDUMe1SJovPzfWFPKs9O1pUyLNqquL7fW4+nkCugbgMGJk3XgouNgdLPc
OLnSvCYpXYlq3F4ADJsN+mD/JDwLV3J3+Xi2rydnjNWlNTsc599+q3RDU8L/MqVWgUvSn/fk2pda
OCGbVIun2uXgpiPnwaeqGQ/bNsBIZB33NmZhb/9hvzN7W6SrvzYCjKadnxuf+nDYic30B/3O7gqY
+zOY69GMGO4Ucaw/pafnaJKGzUXBTk3gRVgjahfpOIMvGuflK6sCxh8r+AM248o7zf1bn3OyWtNt
zqei49p1QGO/nw4CbIOVdLUTWo2iSy9zaBQdyvgyXtKSyoI23rQKshatzlxHX5gJUh9psGwrcxLM
WjTYUoyVYokT2VrRmyN79sfOiw+AXa80HAtEGSpjAYOFRKyEvjTgJtwqPEQRg+ASr22I4ZBTtcIV
ivBEQXxuBF/aaEz3Q2ZpNEDqFLd6VLGki59TbNuPNK4S7qTXO8jd6c9blx9wQho4Vd5kh6unKRzS
7LC5e6LRepBhpMIoB8fSoaCuLSGBEu6nLkGI6mHnLoJa3escuZNeCJtwYX2X6mvwIxIrDIBFNl+s
fPxZJIOGUK9RsayQgVMFMMgNsTFgS1OD125m57HGWKGzb1+RLAMRjc5Iwc4n+Yuh87CGjprXQzS2
i0UGBgCr04VrVUkphZB7pzzsM9LOEtFoQHZIzaYs7xON7RI1E6UCqNFNQ5eInCwl6rZxc0Aa7nLO
O+aKFjmBqV75TEOQ6f/CX/UJL74FPjTeIbWed56v12FaGibfKVOOOfwBs6v9Qw9E1GxpLemdNwoo
IDtwhp47FasgPbn+hVg0vNDkV6gH4uq/fA0CtpVZWdhkA9hie3dm/YCVMIpXMc9euArRCF6h/Lpw
lauarOnQRSkiqZ0B4vTdWWKZsLzGKSF4SN8RQfl+HNLGtDB7EHm4tvYEiG77Zgalig2TPjuRoc5V
S62yrMfKux/EK0BI6bMPshMq3ZHD4TngFTXQ9sJvZygQVpeTZD0dvNCRzRPWzyW++sri6UWcyGMp
RBAxjTNrV2hNHp+GPzhbsPl9B6MCe+Lpq8LUMRMvlUU1k+XJpmHjENZNhtWPixJovzoQYSQgVSL2
L7c9p7kdlqGd1oSgh2sbCvffVg0zuS7Rehl5IB8PzihEfOiYSqkVCZ+RuNgsIQpgW3bJ5wUU9ELZ
UyMy6EQAAugiHlwKKyAWceDeWMtvhJF8g8/lIbNTBVJ7v2fNMPIPBFkNEnglD7TzpCBJAOy5B1vm
MudkFRrhEMmWXH6YFzKe1T5FfGqDmucj0Is7gPIVJ/6MiR/g95r6kal9gMNrYq+92waFwZMdqD49
c9fCabp9gHjy6wOTNbR22VYeVPSPBAx1Hmerj6pv1mLGUMkJ77msd2EE8P5ZxzryC4ElTUVHx5jL
zZ36O/bxPDvGrtcCaz8UYSeqPz7qYVvakG5FP8nXWys+7hWGOv3AoAUo7/NjzEWDj/iIGIFWbU+o
MpXsVRVrW0dRrbq7O+y9es8kaoGOHnpIoTgvnsMkhBo8LbZ8o+RURvfuFc6Qu0MtwbCKO1ACTWs7
Tj9ZBWflUN9Y19cG7AEFe+CjlqRKGZL1D+rLUH0UIuR6iaiDnOBGo4l9V4abBZfMOwFGWGTgVlq5
fVOQAw89a5leCVdt/fvq3+WxdUBy8/+mymLcDZ+dp/Xsmt1WNXe28UE8b9ngXK5bwm7hQRLh4HKW
Ez3v6rnLrGv6mOUnioXg6wLlSoHV76PJsEZU7FVdAmrzYl76bD5DLeFv0IPEjLVm+EiWQLwiY6R8
CAN3vn8VQjvCP2Io4Bds+8p4Jl4dwWgVlV2tqaj+dAeMxVsn6S3aMqCSbJLmG+U5Yv5I6uNc3YfD
F6GWYtrVF3xN0BsHllEbrq9YrHPzAqBSZbHpUHtVBdtqmxtUr8oRJ2cOhLQ3aQzqBwux4LPnMj/l
SHwV519YQhuuIzTDVlcSYDiJlKR/sN/BBesQDYIJxTFHUYrtww8lOCaN5alCcv0kqZ8VIe9jYMK2
LZpHqlqvl4PMHAQjrnrQjs2Nr0jLeYZOgZmdmazRzeuUv4XWIQy16rxPJ8NsBxC/423EziF6Oajr
QBZpHUyXdKgpIs1KDYCxVLThUbxxNs/rA5jJIGekDcsfIzWY6pYy7551hy3znOC/NyX0hQp8Z31/
5sxvzOVmBmf4EJ/CJ5PqGlz+wfLFZEzzF7K59inShFPf7hz4N6XCk+MdoLoBkynPrE66AJ5u0o9P
RKelfULXLdWOeg7XWL5+CCGrzYkYxFrB2OnBGKuzRWzsZ4jz/Ip05wc9cWXGV1EGnv92Nq7MKDFl
nwCLwbvVA38LuYn68PkTypX9MB+FKKmSiJYlRpC7cQyNSyKfJuJ3m2aphuGAtd2ib4TbTNxvOz9i
KrvhOrwKbwCU10ShqggA9JfgRxxlGFwxxtMV5WLZoGbmExXEJnJOa2BwRt+Rr7KwpRTiMl3Rrqym
4tKrcg8x3qoK0VPQoELd7FNps4qvoyId3aS8D51aVhTc5Ir9NOgtgS2j9RRhwVkFUyxE0nCZV0CE
tR64OKvGATMvljbhMju7k+kFLNsC7oM1j6EqlWjCrNknABMspEZSG7g4zNBXb7HLhKRb8Tt3RD6B
m5pqVH1g5JAIhOyIPw4papym679s+86eexIYwhPSBCZPdDFAoDdNFSrpX9iYiL0RalZqzTUg8StA
fYt61T8wsAyRCgqUydCuaDDcPnLNB3/Dqb8YAb/vJnb3wxzeWLf6oCb7lLGSA9pD89ZZypABQ1Yi
Thj9FJZEWcfhlEYVNtY1yZrZ5Vym58e0bDy24B1dX1CpS1uAthV5DWDww8zmfjmPLh1YGxrCnoT/
lmz6edna+oFcCIaWJlIW3BALHwJN6XR2VMscqO95yKB7xB4WhmacAUmFvQWoOMvlGzwCbFTa+vS/
pRtMazI9HWetolnZt0x+jjSjenw/ml08TJq56P59/AnuziMFAubpD0kdxhSnPPNwpT8B8tt8gjSk
CLtTolBFNJZpqICERr3zejNxiHxviffSaLk6gK9KqS8yiNb6CP6JOTNx3LCDoMshz6CZXJdNxq8B
jv1kccSOKUIeiNMtxgHjQS1KmRgbhALfTUQamNhZaBwO6/7udoB3/RPyaXmP24LEznmAbcIL5g3c
rJEYBqhvPis2f1FuAUP11gIPFDWbMC0J2fED07yWcd++8R+UgEvVDHcJul632iOzIRMTPZJOP+Ai
5bONyu1D5Eos38jdtOlzPgRbYQn/p3M8diR1xWen51jCPB+Qey3FnxP2xW+boyFZOYrgSMAwzb78
6UJIXrcg3bVPfU8sL5GPj02C9h2KppNg/dfWPh/ks8wctfW2ptmR6Bk6XtoyVzw0GVhQmqYXh4Ue
D7s6XpD0m4PGjUv6UKIVyPC+H0vGdkQeJHb/JOTswEiNjAiZcR625TMwrEwMl2W+h+7Gt6CSf+4H
Iu5dYU+a4bh9n19lvyjgAdEBt5KcfGmKIyKDKER2D3onZStuR3sWS8SjI4k9dIAOEOg4lZ+yA8V0
qwiIlwuZ0aV6Uq9X2iT+GiU7i3lc3Usyl1Km0k96r0G4XHfFubFQI7JPK6YEFGNWw4oXFmL0unlb
I3yRH9z9Uh+CCLUjU5BZJ4FMiWq8SXVH2VZHK8a4psr+9NTRDSD5T/0fg1xjyLkomdPWiVeqynVJ
bXBduK5PYH6gGDynIxYqvZ/YMJqi0oTvCKvnZI6qcnhiuQ5QZEI+8JEkDaQf/WbptW/dF+0VAHY3
N2UbjvZrmz53lAXoljRhoCuWk6e55j3G9QvuvZVRm9snaNmQUICWoxNP7uez43OimpslMADs1ogM
ff/ttCxwToTv6aQqtqjR/NYIs70IAiEbNEcui8DnsJsIRApUAONGll2/Zbx2gEbr2DFacaeIh1vQ
JgSTXaGq4tTfNsfrxOSy4a7e7xpnJfQ03JBDZ3vQPW1RbW6TwtY0gs4v1CObDj5MIm1oml9LWBE6
jOAx2jIJmZokNRJXEcPpI+Z12H7doreysBlJPbZfFLD9DPL7UZYdCDflvS8jusCJGqELmjptCLcR
ard42/q5xCnHyiDvBNHMGKbJWk+dcR71IUmjKasLkx/AGjw22iXiznA/XOPFhsNeT6DUdOGWnPI4
LSZm48Vw9BlRcrgWSTPqXOYTm348fUZutKeC+neNJSgXatQTdfc3nDq2lEK1GuKkgjZKOkjRglHe
3BWdC5t1MtUUSreyvmHUQuIMbQjkHhNpc/sEjKu64SdbdPzZWnbjGcJJ5MjIsD8o1veiE/VT/tXK
dO0iw913o2HBccS/2P9azXdhh8ucWyqr1s+76eLrzXFt46A5EHdaFKijc9cAC8woMgeeanSBxMsx
B0fpJer21sCAPh/ENyMxxOgR2YUA0CWaKpZbO3//LLtf2eyxVP4Ty96alN8hOHenNCS8tBcCahZw
B6uFB7fVP3qVZgCnfQEJkB9yUdYcWUhtRfVGbDQY/ebbcWPFZrhKdI8QH23JOY+7DPOo/z/NIQ3o
mYl4lWOKyuToYlVTZk6LRWXxIAUVliiGFVo3Ir7OkFt58YDZY+mCFhLrY1bCGAM4UUix1LyjV10r
gO3qvkBng5e3qj2g+UraTAFUVJKim2KZAHEhRIrLHKpp52FDDXjBPz4RUEvkHfa7giUS9Alxg7Rr
tc0Y3U9fj2KLYrrWkpqTVPKwVNzfby0IgDA9AxBqGTMV5MeokmGT8bn3/38VgHvBTeTA1zS1FR86
G5HNJQ5fqVMxw0mLi3gRczMmvnrcCzM2O1xmp9aBVfFaCMoTqdzUOSxEEiNVFXqSa5l182MuROey
hGhyMoFALOZ9Fd/Fs+dXQNcF6/x408ip0dMl4zHh06yLKNXjD/IMLdxjSVf9RbHfg9XOrTxoaWOC
VMmfv1yYSEXQNa0gTKXu90kwpiVrOIEIo46z7taa5ypbEWTvaOU6HRYddwgfEHVa+zs1xwRe2BXR
cdsTTjy8l0RNzJHwnGlJwoTikuCAGVu+XjuNE8moYJwgJ5IqGKITu7O8s2RAVLkiOSNVzE5GcrVS
bpb9K57MjUukTRtpZ7yY67PlTYQUAd3IYT32xkfSfqgX6ZCvVZIASFUWMsZLPWGHYl34pu6AGUFb
8nW0v4RQSw1e9GDjnf9kskTbWbIYu72DCB19cvNK6IHUhclLgG82al9LtmIPXLCyLFPqtw1IDK5T
unJ94gQSV4V+VFBl81VY/1bynDBEt3gaw4ApONlwSTuivmcg9DA7Z9ZtdCQ2DJcU+b1TNsbiBQ06
mUiGvenQJc6xcLn3gT388hWlDAbYbMWsXv8r/QeG32R4JgAPU7xb8JkcB0yy0AMVX4hBJbSiwy5Q
k99TznuFEwAdAYtmlZl1Wn9ORwNhPY7HLt3u0Vw+bIX0oOr661EdRc7+crQ9RuQ9+M9HMs+9ynvu
SHqHiBX5IvZ2vkEMhH4njxvLKyzyYQfYAsq9ZEBco2BIQUAgmFejc8CrnRFYFNzzfRo1cRLegAFQ
XjE6YPzovPOeaQ9o/RX/c3I5DPXj/hM4t91VFjx5qCaP4H+l+LzceyMGi69/8qvIM9ASHzeT03Mn
Izeo3WcNahhE6vkI8reuY7OyzSupAw4GsJgYRYEL5LHURYANkQkh0pXGHz+f1328hTt0Si09MhNB
4mT32rzJVvRbLV5paI7ptSE5tM9qZeF+hbKOZUfUX2wooxDYu6CYK0mLb5wsV/+W83IiXdK7irLg
M/k3dODiXRQDgPr6b8aUk3+ZuJNgitH3nHcFe2kOcOSbn4IMbCH+ic74tq5Ew3wGWrmZQKE239nt
l6xia+mXKIbdYGXnEy5EjDhBFrrE6EGA1ismK/5B2jOgMfD0Hr1NfsllRsCdkQKbTFxvJ6t3iODC
z1PgRCAPXNeT3TMUyEzN5ewDTV8NAt9y9qRNM+zSViek2tTjj9/S3m9bKj6LW6zblyePzDxNWUoa
HHtRTGJUxmjFRw3+D2XN3EviOwnjWDKrs75ZEfd3cvxRCr2yvrEfrg/0xK2QSE+Xe5Rj23AkJY2q
iSUHwDQMb/S9nZlEQ5weLMTlhvAa2q35+IE/w4sP/EqeA79t2AEA8SRZZsyAWgGyCJ8qD+1g27i3
O2t/z9DUA4FJFQ8cyGiyBiWwd+0nTEQLa4XnEMAD1VKLrOnnrAyWUCtX5vVw1KYuiMmLDHaotW99
R4bwhZhZTRwT+rmPmekB6RFQXtUpSUv8WYRS/oQ9D9bUdlNDu+lVkLMjkV3eehnAKJ93ycEukkNu
XTTlcxD5GH7gn0IrOurdTTc8d7SwlNgXEX0UjrEBG9CbJ5CFUwwZwsUsUTf5RZwPB+UytsKz/zHE
g/JN81WkjJP5AYswywluBQIqS2PiCnnyxxXP30iMyZ7KrWaHn05DMBenmAZfJ02P8BoRbJVqETDX
mraWZLXlKc2QXPewB35Uili72W+RQvQdtegX09BaU1uylIGRY0ZjiJs8NhpWV2h0LYfzAUOmV5IR
SSYfV93Q+W8Bhi09N2gLfSLBt+lKQD28AO3lU7C3amgg9/+FZ+wEhGrBZVVgpEKhNo4aNIHHuzIE
ZejB/WguqmPqFy6yRFYb5AJ540+jSl9LvSqBZbBSPM73gu7R29WVnK0uLeR2T/LzxbnfHgvqmW6/
H5IXeMY//V7h+JcxxdD7X4piYZiFPMR9JFHACtSab8kiVErvHzZT3gLkRg/PgtSe9PwaNbARPk/v
OlTdf9u60QwJGGa1Cma7jUcGLSzZv6u+g13I+t7LHOfvea/2KSyNKX0IzplXTyERzTx3LET8MFIv
gKX+fbL4Cz2PN6/1jO1stc4Z89ytJ62/gyC9vlWcIL+d6wov8CMXS9YkOSUwDoMekLD7XF1CpDiN
x3zRngErxe8ImZvfpWh06As8kTIgvBDO2jkxXnRYs9FZ7vdKh0pYZeVriT0HrybtvhfFdk/TvjhY
6RSPpLAqA40sLa16A/NG8K/1i+sEIub1fNPcGEI6L6s/TithcPtHG1LADbzJwAU42tfPn0/BPVaj
UbUn8YRdaTMUXkjV2jV74sTPmQ2wbTpqpBRU08H1rZ83vOuze9eRhOHURhCVM2iOvLeVOoNnuMYV
81Uv2HTroNB2TO0zEOrJOORukx+lShEF+UCq3kkAo60jHHDV/llDHic1EIHJayMEBKG9dtyOMgKp
/+zwEIyQQgSAnsGHqCOZWNfv2sLwS30Bbe81X6GSfvaSTiHEhjn/JzS55HXTEyf5OFuc4Rz61iqj
uUHwiOxci5bRUmkBRTqvpNXxDBV0OAviMTLBUwncaOOhFS3p8kMYAjWn91Y+PvtYoXjeiiF6fYiL
CNvudLDvxvXaRFNpNxu6BJyzjtov/O9ua8jG+2KusVhLhN5mHK8K/6JnJRqC66uBw7GTK8WqynO0
6lnrQmRdAP9yG2Sg1kZ3rz55mHf7Fr+Ewb0TEGSXrloHVRVT5VmqFsL0j4ZSimjQdeV6qqDf26m8
ll+yrSBwCb775PSa6rCcv0zGBilsriXXfKGC7fj5q0uvfY5IvJNGzXg7S/iKGVe4lKczkI1T2QS3
YnMCWqT7acqu9Hju6R7GbJXn3azdgas3seTNRFHH5YhN0FZWe5qbUXC2Oz0I2KZpYzvRzqM+PuoG
cd4chrvaVE0rQAwWRpdb9GQTDuegK5bcklKMdTNnWxoU1hzvmYNNPrqP3LoUnUj7FyGdU2abPq6t
9rMRtBxl/fr3zhNg0ALJNr2JUNQUS9gQAaeQJsSEjUwybf1H/dZacuQPSpPPJ9d5Ew7HkrY/t2al
Mg2L0uNWy0hXZwtve/FlRsibG6mUSiZlFum+QrmvLXsmxRS3soB2m3gF4tSWuVBZEKGH7xd+L5wR
NeBwdANCcIxvhTGgC9RSr2iGddcyKJqrOkmynr3AT/iMtqgirLFwWy3MkvRq/cUD3InNqQd+3d73
65JGX7AfT30OPkZc58mIErPMxnVd/+MOjdjeDwzUieU3J3XSGt3joCnzWjoA0IrbbOtoxXBe1kcE
N9fDTlDo69utEsuIWJpe9VsnpL1B0wKAFquQOxGupwkf00DgQL4uNEXwWlJeojMTxDY/BwU/y5AB
z+kpX9/2dDte13MSZk0KZYn7Hw2QLUkzUpPaK4ZIlS9dJtC2A+o2Yt46NKqcQUoTZT3UHwrmabBg
PZNp06NN0oLWi5iHE4DC6ara5ikHSUpUAIdbrm8v5XQVZ9gmaZ7CcRCPuwWqgloG2cnIubTC1YM7
nGYCAPZXRMPNyuJlFpcR67622h36fywZH7F5riabKOxYoRuPL20EuZGyhcm6XZ3gmVXuf/3ro+1q
7TjZPBc9z/ne0RPf7myRtoi5HnhF/0r35tSodngh/RX/m6xbnDKm5IjtxdsCL09J2efr5R1F2uKT
dSHzmASgk46aZxdQvELbsDSsuXmFMPJvrjkrMZeLc1jBFF0KKWET5zG3zHP+Wr2ARyBuKSVoqX0D
CpY/defKUtavPKljeTd7Yq73Nm6gB8cHnYXq6lqVAreSWZ/CVwhsNca3WdHgrlaAskbaO1abgA0y
c/sUnmXJN5jg7YmY3pne/9PnzPXXk2zYsMycYLbfY4rU89EN7tE51OPLfxX+xbSHEq+7zAmDMUh6
vcb6E4lG2Q4Et4lolQIj7c+n3MgmF9AIcladLdi7LbnqpVZeP/kzrok9nmVnvspHHJ+bYWWTVSTl
qJ2p+Bptg5XoT6aVGjOSnczg0hlByFM/LnD8pe6YqsLaAajIiSdHG1vRANda5GPEx++xvB0NHBDf
wyUQLTc85QECPJSnRoBvnS4LvXtXxqCtztLiTaib3LCBanhiuA/6p+RJQucqi2VlgCM2Hk0XFuXn
ItRgKerVzG2KwfwGFo38wsOMOKbwPEkAyv++1vpVWzucTD+db4Yd9cHQ6dHRYpLgBFFVkIcfURMp
V09/428Rug0EwJm+nWTtEGLeDmidlxhTFGm6pAIiVFAnF5pFjzK6tGs86pcuFPjeYt14Q4mpMHtC
IYhOXw8Zek8GjtNv0YFXqB/gvD5WHUcxWdff+C2Oe1tRO3N8nZmHkuSSOFYU97PCY4idhLB3gpR0
+HAewHggTgFb4xW8MVvzxLon9yyF3rINLMOahe34Tv1pj/kwRvIJNFOrOlXpRZukyD87+NIAw5oQ
9b+2R4N6+h5qrSciSng/brXhoXzApUftQLS1jKeIwWUC3MoMlu31UGMPhMQ3wpM0JXDHCFj8uX7u
lw12zxWJEQQZ3fhhnQwQybIElcKMF+vcDdqt/IOhkCuMoOHCxR4rl3f2bQg2i/DXm3Kjq2KGV9dU
qBaqK+SqSs6A4mUuzGkn9paT6uO0V4WKLuUuEKiYKXGrujOjN32nsOuA9nWBOjnq4jF7E0n4EI8t
6sdDRTP28wapejaR7lUrcyyqVZqF/dDUOt9+6aYtZIKRAhip6eEkBHt6eGJeYhlOLwoEHDw1i7uP
pR5bf7FNUs9h5GUTDRzV96ts2uuFT3BKrGhxTH7dhWWjls7NDvHtU1IAncZym/ZXXdoT2JCzg3hl
bU2KiTgEiaPcXcIerZr+uned4dp9Y5vkhcvhat9jgq8BXjYc7WVzlVcT6oS0j5DM2/ENtvKvkv9w
53crPuGsBxm2fQGOBXl0bNytXj7KJ31dxNzw2RTV1qzpG0w2owFKozSoAemIw02B9R7uFpC4epX/
QlMfWgAGqr97nAJULPsI02BQBH20oRvGUDFm5CHz/UCbqNqLBDNU2QYRY31rggWhEAfxzeL60o3d
E1NOIe6QQg7N+9lfbORmDZmHObLoQFo5wG/pVGrRP5mwhs1FiVYqMQXl27prZgVvvybbHMuA9Kca
7XfaPv+K0knXcWoo2DgP/52cPoH6Vy2xJgTNWxzNXepr7lAMDmZdER4s5/N3c8wA7TdeK2DM0su6
r5KrcXQOfRvaXOKT9EduDnfV8V6F275r2SEnPG5nzukuijaxgbhnjakaXcAKU0b9eUhJcBXcHLTT
B3Qdim1s3USAAR6elUnEjrucjEY5xUos+aOjEJygWP0OC8n3y3/xiEG5l8btYmTyZg2v1zkHWen3
nM5ZuYXLReAdm0RXV+Z6D5rKWEtDZft1QVeQCafqIyePoUrV9z/XKw/TujAQo2Ek2iqEnLNeteqx
w4qDRbD7RZ+t7q+wK7YX9rPw2u/fdyRAuMhSWMGi/v8GSPvHHfqtmTpDj7aKpSU0K2MJnjzp3885
p7WUt7MeDJJHBNGjmTWp/6SnKe2WFFgEKRV67HUoCAYSyJ59u4tkLDGTno1e98fKZPT4kk91pQvu
OReycwkb/qAmWhdJZqfwvaHHx2podblh3y/sRVH2jzYcoz5yV3dsLQ966OgHvkoDzfwGYrI/sajG
hNtLK6a2nfuSZyeuO+dO1fBS3zVvlKr+cmgDUsnGfgIGN2+HaxUc298YI4ipePFTVQZZk/pkUykq
zxm+Ef3ITmOgV+7vgzku/Dom6SeMrsLlO3N73zmhGQ+YM+RcfmXx/QCx6GHusQNel/igb8j2z4TA
WlAk5If3Ea2O+2j5g5v7PZRr3OD9uR+k4GEgrtVSTjTqUPuvnRmKAIajidXL0cGTmUYUQIyP9YFK
Gzfgp9zcXTLS7n1CpAFnnXUdOH6NXp4Z+cI+sXD8TWEYplu4QxESoirjzxczUtHo4sne1+zVjjrZ
9TK1jGA23R/8jNeIiXmLdgi8rCiuuscimCPK7i635sbDJ0nSvTzWnyv2IfNBy5Ph6gG+f0tlLEfv
QITwxWHBnK0g8EwZ5kipcdAnqVNY8ZXMoZP2krjR1Doldvt21oqAf/f2ziEmC0J4OjqxiNelwIoF
rHwarXF03TQI/BPv4GhgfBNfvqyOn/bznRNR/+Lkvm75qdEGbCJDcUWHx99T2Eltgfsn4XtBHJnX
PMma1HOEEpeVNXJQokdfFCqr5LS/UIw/97DKDDzavO1+bzmUaZkY6Y6Kn2u0jQJ75Wx7DVXK5D0n
Uo/+V2mOSXn5XVtMSULF/kG2wwh1P0r4DCprbvA4/CRYSa8c/IKS3WijDRXCiouOobwHPGYCG9Vu
PCloGn9yCzTWZplLxkHjvMT5iMYUHbSq+mORKJl28VX5lazV7HO+06vD0KtnSbD7JHuzw7CXvR4X
v+CkJfeIUr0V8H7+VdycQE1toAiThVsNuojaXQlPMGLKAEWvrlck5IwN3m3KmXIziC4SS2ny3JuD
VwXKuBxs80OkAgBecfScYPygkKMGAettMe7QFawA/K2dPmyNcZhSQbA/iei1V8dp6bckal6NTVyo
JsY32eEKjipT6meewB0JC8l4u+sgNooEahFq/Jo7N49ipGm98DezA9dlrIPWPxTMmQvBqr4N5bdC
hfrkqtJYVRO9q5mz+tNGO7Zb7HBlU06R/j2Ar3ZP/OM5rrjCQ3sqDTa7v80LAWhXOXjkTF4AnUD6
zMsc+8nR7w7dM72WvcxCnTbA8BIbPHixbRMqUnf/IOUIBJ14OK5/yetNSuOrZWnsjabmaUrE1iPa
CFnU3OH87MVt18Xec6oWPxlZzUyU/s/q63Aw4raO4K0FibPYqAtCVlEW61tU/amm2XPpwxvRMAEz
9xybl9FTL9VoYaHCqzj9IexQmlSpcKGyY5Q5JYDlziBuFAGqHjl0OgEckfwjwoq/uOHX5nsTnH60
ez21bdEUZWa3q5D0QvEEY/vkVRAOySow31OarFR6u3OLp+e7k8I2+Y3k6fFayZFtM/fw+0xmkilB
fTyIF6uT4feAsPLXGeUkLVhA1dYJapODVGVriG4ru3LfCrhnyN1tOrQ1ChgsiiZX6cnWGlmP3zYl
fMmWXSmMiFxFTjWjzqUTlptI+59hY3JZ8+TIaSP94hxKRACXs49CCo4eGJI19Wne8ral8bYxEtpp
NKTEy8I5YXdbk1hU6sCQ1um6XE6QEgLLjIcFeAT4OjstMy6cLvZqGMLrTnOa3ZaH+iqX3s8Rk89A
+nM6rPfD3qbYPnuyksqjwF+jao1wYMKZ0lQvB12V9zNPMJ7SSbR/2wwmDoMwn2LvBRGSZwb8XPOk
fBn9ck5BOmaOFCOmIAUtJfpB+hkMDG6DZtjwrSWi9MM2F+9EmZUx8W3b58S6D324WFWfibLnlr34
SyTG6KlH4yPIjzlh/ssbgqfQzF6rVDzTaljMFyU1zH1MkWHnun4UOwYGZtQPO7Zlx5PGV/bkquGs
necSTiC1OEzdRESxZW3UwAgMu4jjfzt8CQzcasSJTfhmU++i13SVxKprCvm35wPgtMwt6ZRC+7rl
aJWyd1KPrtdiuuaPfOzXOvGV1mqpGOrH13XD9zTDkrzK7ltrUfeIAAw/QOZiaOHUcnroCiJ4Kb0j
nGZVq3pMzHRBZ+l3ByMTEVOk5xLnsm6RRzOMLjqPUlY4Gs5cO0HfNGXaGALdMsfxPcKWc+178IkR
OklbIt2O2U5uJPh3iJM5Bkyilsy2OjaZMakCSii8yQlh1XQ5+roHDAy79UifAUujUqtRSY3HpPEU
H8BoG/6eoUwH/K/w4r6IEueReIfePp3hyCooexI06MchUcUg0dO9tpDoA2OW49fAFkRhLDmWhIDs
uEQ6y0f8IubO825ekE0T2ZprG629VND07gJLevj5BV7HsSbtIvWbh25Q67nOsHleTUMXK4diU4Pj
42y6Y0rbLICUDbyMQzyjOdLapWmm5KSVPsrv+M6DaggV+d38TxS4jzn4pKqdvWOG2FmcIDJbblgh
mF8re0ezJ4hgClKvntqEb3mynfkQP1vQzCzJcVkcyzaRZsS4OIRYoA+R1pJBelcR2P7wdgD8I1J+
ENNOLcoyPAZbLPkpyk23ZpJwmfZGsrQzy0lCBEZN3KiO0GRJmDE6Mp3C5rRQ22R1qZrIBa6+qoUW
gYK51uM3KOMwHMMDjMMF/LMOwUAJtwtJKmdm1qeli82beZMsHTS/VRvvyJbmWUKRfOT2icEKhHP+
4XE39yZBf3JRBAPOpGZGoOdGhPI4T1qMHBgIdbwXbnrMnyCWnoQo/knSXw2wLydXWchAnRzEKctK
daiTTpOlUlLnF3eBSRYhUET30OiWvGZqTwGXK3ZY3FVEbCZJBrXzm9fLTKCb3abKxu3UmnLjxBvI
nQyNdXWYPrxMttkMBhAyDJPjiec/Mf95zeER+911Og50jlIqZkcYqNQhsSkJ+5M8rMhIJZBwe7PD
ZK77KhxifTDYNnBX8wqZKm+0Pi72vMmFHy5PttMnO+6YM4WwID+DhkZw7qK24udnPjyWe8Kkrwrk
hgT0uVbOfYm8/rxcgyIqK4LIewCheT/++rB7nVT9v4geFqrMtu1FrSRmeRl5diQV7uJXZkQ28JvF
n6ILPWyosjuA5P0qJlou13WI+YB1TQmybjicWk7KnPBihcyH9y3oFQhKIN0Y7Zkk0TaF/bmWYOOJ
CzUsJAN+Yg9a49dmhvd0ARIb+R7yg8AGYpSVsUeKkDE0ixpJVbe/SZ2hOZq64H5bNUmL1k1WST7a
1zY7y+I0UpnZjEamObCqvEbceXEUZN93Ow8NAEuK3q1jeEqjXBVLVqS3qKrcd9+p31jaVhhAV1x+
xjj9jMtEQXa/79jFDp/c5JAp81i6ghl/Immi0NUZA/BeWN3B0cSinClj2E5W1nTuCTg5A0vUEVGG
mEEMztafQmU4h+NmqeM7leZ2+lls0C6FL3pVQQVyH2rOZkxI2lVwHQCcSve4nj74BwT7RaPKuy4v
Ewc9eSA+meAGCe+2rS6LM6nc0LDsoQCO0vB2Ttdk7A1L4CQHUWwEXaIF334jljDNSi11C0/x0/To
vs7neW9RS7sF/0dbIqOVSWvfGLbcXq4Dquu+w0Dym+zAslP62valnuXnBrfGk2cGqk3cF9A5EW+h
Ass9iLBT8HZlT96dDL4oR9L75dbcfcABznF9OILA5U1nwluWg7NKcJ4eTWbxJba2gq0KXeGo9PbL
jKJR+mIdEH7kbs7SszDcpqdOJuWzFE5Xq8pp98/gsYL8dN5OYgOgZkWe2/1T7Gl/wHngrXFD5AZ1
391M/bKmNFN++3TT/Grf6eZCnXy0bilTtmLTNpkd5WiD2O7zC9Mz5CkwSd0Id0t4Jz74Jz9qhAWx
mCnibnSbDXNYut97Ep283J2d4Ywae/evvZMvXfLANprJHEf5/0X525qOQyfkvN3sPzMih3WemMeo
IxL1zRWfLK/mkR8IfVXWrS4Rf3uXQsGQNgo2GM6PArN4jPsNda3CkyNScutFGVdSzJugkPwOszAE
mhhxsEMiKEqeaSJwc7KX2s7+v+07v4kB7lN+hPyHusPJTgfAIkRxD9076dfmgJx//SwlsPPXHDbf
0221H6yTvQnuhiehco1WYGfyJUbgHfGgJBnYqGn8PODLl5/azpUrrg5XYYFlfyAZim1gAMIUrIu1
Pld908235Q6YoZfHZ8QA2+cfIf3tIGkn8kftdN+gGMrw4rR49zRhdSBovNtODMzwnDIAEdAg26Qk
Gq8BxDRkjlr/cjlIKVe5WlpoOfy04M57oxDutPy2+UCQyMHLxCkp4XkZwbn7wH1D0k8xqNN3RYlI
dZPwP1mL1B4FWJ2H4IRCc91l7TsILmiRpznaEpTLrhDf6kRRN2I3Zrmr8x0cYNyNsvm/FG96Qnl1
McyhLtevIh/LrJ4MylCtC42UA+HgNJ5uycdF04kHdB0M0Ex8wIqc3Z/vnqlqAXBI6XdpHzXjRw+S
k2eQyHwCt3lfG0/0VYAEHlidpFtqhvdxdQoDudC+zt9kLL4N+mcrYdCg10f7ysqsyUy719BAJs58
qC+4h0YhkY09L8clsxoGKu3mMTZSZjd2699AMAURbLR7VeZ/Z8fpsXk2eydSLC3wBAS6dweeYiTw
o28hT24AmK/iYjjaViL319OelHkWK8CCWxfuS2gsTmvNVk3WD84ABsX1sNKxx6SNIFZiqQFy+sN1
k0mwQFgDcHKfJ2R39pRPjgvnIRP4cZ77nKVKQUbXx8OnusgZd/3RZqWLO7sE77ZNhbvgnglKrRw+
Yk1YXQNOXJUHXBB6povTLiu6PJp2E3sUb1EZGqbNFCvhUNIkjZzOFc4FTZigL1v8SSvJYDFgIvlL
N0rvqJQzP8zEBOBvffgYoIRt9EikY2MWaMUbJznPVaB6Lsv1ecHz01oitReGQar02OH363IQbkgR
GQbzHUrhGLEDV52Y2S+fyRRSjrx1suODY8XUfaDc0040o27qkGJsHLbqBRLVLrdpdeeRD3wVrP2s
4OELjLj5ogJM5xRjKAyGIElMtkGVL4BCTuaHzQJHhPAwRRM2uh37MCeJYBgK5OGjL4SecJlXYo3f
X91ZVpXUBT0cCbGWa0EkOtSjsRSW3jIsJKNaK/YzZ5idTi2gpMTRwoibF6bEOlu7yH9HV9OCI3QT
SN25BkI8D/lbBDqYfjZPndKVNad+kin6cwXNlIbf/Yttjq34Bs4dS0wqOFlK/XOjxe2+8i8cr6BU
RRqe2fbxTu/yXTFHBqG+mzegoDBW+eUR21DaDZvZVHn2e+h+o62BgX1Y9ufqH8v3b3//gHn9IYBZ
7VU++jKpa6u2QdI4OK5ChupZK8bb+PwwgcOYE4Tw7svJiC6PF76zMOUUu1uKOsqiR+9+VSbhE+ti
kH/7zJyMnxLp7WYarwMrjQNURi/bUguFVXlHlE9wx6SKsuyiWCb2YtsUoBSCvWRnXnWsdR/iJpRV
BahAMizikWfT0E2yV4XiNkmA2AbniIwOrExM9VPrG7eZbTJ1u8i6Qy+e65CvrOwyeUacfYrf2Zj2
ZMCPrJhqgXS9AvcAG7dKgOFqmQny1iMO1epWsc9hL+pgRr5Sr+0J3i6OraJgeqh7v+v+qRqbYDSC
v4+XVCwiiN2aUb6jBFBWNgO3wDaIJu4FLoW1cjLDHza0nP08ngeiR0LMm3gKvRJO9UXTMANAlmiQ
llEwO8GCfi7niVYkPflizO51FC0Ni0qXORZquGSA9j6e24Yx6dTvxv3JzTy6PgP7zej8R/EPRWKn
yg4awtRrlztw0HHDoiTAdYtAEouVxDre2aLZrMfFyMDMeki6saSM4/re8jkhgyahsDPRjB90NMFm
z+CQbDLgdfmBbet1n6vwacbhx3vcihiP18dPe3A23w53DEmY/r1qhSDMAHiyGoKnmbX4OTC+Oehd
y5EHCXmmsEH1YXk+Em1qCQyuW+nkmNtoDj2sE7vl4UEcdHuVH7imH84CAACpNnGPzyYahR4EjHtm
EojgSSW5tI3S/aAkuj8QCrvyqeW5xrkVCSDQYjMpvSstppZMskWbMfXM0qcnMS86Bftiv5zBUUBm
44dspXdcTQajdL9J+aWS7FAVYcduFzG09vIGyklwxGBM2Di5587PV7fnNDWJNvQygI/LCVXxSlJ3
S6qLU2D3y8QzClFufOjO6JW5QLjsdl0sDI69hXRJLbs4S2QfrivjhGYnVfrhwQqcRuh11MGckYt5
R+rJazP508V5dyUY2lv1LH5powYFrqI5FM/DBDV1/gRdVIukgXWYIjpEUxsCp6A2auFuW4/RHQsJ
aKjlmWYxYvg/wNuLL74dKlIY7COsmLmtLMzf2rnAz/VBUNz6B1olQB+0SBYoATqbrBA7wrbzCkB2
jdJNptCqoPk88SeNBi0kkU+5/0sHU6xurDHk3f84V/O7gnYNBKZU409+zuRuj++NxpMap7cUQqlA
T/kYrla5F8VvVBUvMZiOlmw3ln69/jznGrT4sH263PReV51egDtW3VFyYlLs1A4BgrTNGPpiriAk
lfKlWDpIgXj0GJQ3VICblENCxTmLhM+0Um3DoS6mJ+dSuk9qDk44X6if8SSN5J65erZ8i6A0UIig
u+ffj9vfAutFv32V7nKqOv+SMK8m4b5Glkym8AmiwSYkwhNlysCuwutr1D2yAk348nt06mKUwTOf
pD3eIzPXqbmkgC9kgUG/76ca4KeajsQlVt3SQa2AHts1Nm6F72NRm/Pcfmgy0W3qx0ZQfeU+SEYE
KeaRvcQFlIYLsiHXselHHPe/TQWVO2Q9TPVH68QyEIsLAozqXx1hZJk/e4KUhjSCc64OA2eSeIsS
T4F150Ml1i+vAbHKwgZoQIdMWJ980Ha1xgq38yLSKxvF3nrDZVcuvrrwmnrgo0TCWUEfQbAiHD3z
Sq+pnGuKiMohm0VfNS76z1sVYNspqgaKEWaipp2MymYrxWUVx26EwlBEJvoMFkkFrorb+yYMy7p4
QxDXzyQxztVlwIWldkllk6P4F1moXWLGeh7GeE3XWT0YyCoE1TZGkxIZKQg6PgCdGKYH8gT68ItA
mRcqFFGopF+UJJbEsisCAYBBxq9Hyu6ZnUko3q98ujNbi+5x8QR5g7qUWihW/dZ8vCIDE/LSIB+a
9SnZBo0xEUJBN1rpnle88xWhPP0w1nwb/KaeWRFz7Fm6XrMf9rAork4LrFgtLEkVLT5Mja5ECLDk
PSoQs8DC64KpSiUn+aLQwVxdgV05GteCCx7pDUDR51VjC+r1XwMfvElAsFjhgUWKCeOD+cFjDZEZ
kq0D9B7YkDfMkviXZV6GHZ4IJu3tYfXIX/i5S637y7FP3Zg=
`pragma protect end_protected
