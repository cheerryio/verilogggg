    .INIT_00(256'h0206e60b12101f010250000b0202ff0002dc082063e01f0002d0092068728000),
    .INIT_01(256'h0206ec0b123010010207e104010200330250000b122280000207e8040102df02),
    .INIT_02(256'h025000050402df020208152056501f000206c43240d32077025000040102057a),
    .INIT_03(256'h0207c02056e2202a025000030bf2202a020815205652202a0207ba2240f28000),
    .INIT_04(256'h020815190012202a0207ca0b01f2202a0250002f03b2202a0208150b00e2202a),
    .INIT_05(256'h0207d80b0022202a001100202c32202a001020202ba2202a025000364222202a),
    .INIT_06(256'h00bc0c0b0022202a00bd0d202cc2202a00be0e3241f2202a00bf0f1d0022202a),
    .INIT_07(256'h0010802078028000020809202d52df020250003241f01f010208061d0032202a),
    .INIT_08(256'h001100010821d0040010002f01f320770207d8224501d0010011010100220568),
    .INIT_09(256'h025000324412056b02071d1d002323b50208062200a1d0080207f620590322de),
    .INIT_0A(256'h001101324412056e0010801d010010600207ba32441322de02080c1d0081d004),
    .INIT_0B(256'h0207f6050402053c0011002056520534001004364332057a0207d81d0200109f),
    .INIT_0C(256'h02080f1d040200370250002245022bfc02072901002205060208062056e2054c),
    .INIT_0D(256'h0207d82056e09002001101030bf2500000108020565200630207c03643a2004a),
    .INIT_0E(256'h0208063602a0d0010207f61d0800b0000011002245032046001008010020d080),
    .INIT_0F(256'h0207ca010020121f0208122056e011ff025000030bf010ff02073a2056536046),
    .INIT_10(256'h00100c0b0023e0400207d8202941b2000011012028b1b1000010802245019001),
    .INIT_11(256'h02074f0b0020d0400208062029d090010207f63244b2f0000011001d00201001),
    .INIT_12(256'h036849207802b00c00d008202a62b00000900e3244b250000250001d00332046),
    .INIT_13(256'h03284d010002d01000d0022056e010ff00900e050402bfff025000205652bf7e),
    .INIT_14(256'h0328510900d2d00100d0022200a0300f00900f205a8090010250002057a2d011),
    .INIT_15(256'h0328550900d0900600d0022500036059009010364530d0200250000d0800900d),
    .INIT_16(256'h032859014400900d00d002250000900600901136457090060250000d04022054),
    .INIT_17(256'h00100c0b0142205b0008400b2150900700095001300360600250000150a0d080),
    .INIT_18(256'h0131000d0082054a014808143002500001490e14200090070011000d01009007),
    .INIT_19(256'h03686b011012054e01d100030072050a036861143002053e019001142002052e),
    .INIT_1A(256'h00d508224682052602500014106205480018ff3a46c2054c0019ff190012053c),
    .INIT_1B(256'h0018ff2d2092050a0019ff2d30a205100011021235020550036871102402050a),
    .INIT_1C(256'h00015001a000101903e87e250002500001d1030201020506025000090082050e),
    .INIT_1D(256'h01410e09c1c2023301180114b06250000018ff14b063e0740000400bb1319001),
    .INIT_1E(256'h00190b10ba00d00101180809f1f0900d03e87609e1e2022101400809d1d2023b),
    .INIT_1F(256'h00084013f000108000095013e00206cb02500013d00206c400110410cb03207a),
    .INIT_20(256'h001102204531dc9303e8872049d2080301b90501b00207d801981801a0401101),
    .INIT_21(256'h00018020453207ef02500009d07010000018ff20453011000019ff09c073607d),
    .INIT_22(256'h01410601a731d11201490009f070311e01410620453001e000381f09e07208a4),
    .INIT_23(256'h0011020b6121d1160149000b511320a20141060b4101d11401490001b0132092),
    .INIT_24(256'h01400612e602f23901400612d5001220000a9010c402202a00008003601320b6),
    .INIT_25(256'h0140063e49114008014a001bb001410a01400619a01001e001400613f00000d0),
    .INIT_26(256'h01d90b2049d1d04803d00001b01320d001da5d01a741d058014a0025000030f8),
    .INIT_27(256'h001104204571d0b803a8a12df07320d301d814204571d08803689f25000320d0),
    .INIT_28(256'h025000204572f23903a89f2dd070122001d808204572202a0250002de07320d3),
    .INIT_29(256'h009508204571400802f5032db071410a00950820457001e00208b82dc07000d0),
    .INIT_2A(256'h009508015001d08802f6050146c320d302f504250001d0480096082da07030f8),
    .INIT_2B(256'h0095080d0101d01802f6310b014320d802f5300b2151d0b800960801300320d8),
    .INIT_2C(256'h009508142001d02802f6380d008320d602f537143001d00800960814200320d6),
    .INIT_2D(256'h025000190012f23902f606011010123002f53c030072202a00960814300320d6),
    .INIT_2E(256'h02d5091024014008001100224b71410a00160714106001e00015ef3a4bb000d0),
    .INIT_2F(256'h001300090081d0980250002d209320d002d10b2d30a1d08802d60a12350030f8),
    .INIT_30(256'h02f0162d0081d0c80208dc2d209320d000b1172d30a1d0b800b01606010320d0),
    .INIT_31(256'h00b01814c001d0d800130114b00320d302f22014a061d0e802f11725000320d3),
    .INIT_32(256'h02f119250001d00802f01814f00320d30208dc14e001d01800b11914d00320d3),
    .INIT_33(256'h00b11b14c082202a00b01a14d08320d300130214e081d0e802f22114f0e320d3),
    .INIT_34(256'h02f222110b90100302f11b25000220da02f01a14a082f0020208dc14b0801002),
    .INIT_35(256'h0208dc190112f23900b11d390000124000b01c190e9220da001303390002f002),
    .INIT_36(256'h025000190f60120302f223390002021d02f11d110072f00202f01c3e4dd01004),
    .INIT_37(256'h03100000c000100101f1ff250002f03a01d0ff1100a01000001200250002f201),
    .INIT_38(256'h014006204e7202610140062055a20258014006204f12022d014006204e72f024),
    .INIT_39(256'h01400e011002080301410025000202800140062055a2024f014100204f120246),
    .INIT_3A(256'h00b224141002028001003014c06207ef01400e141000101001400e14c0601100),
    .INIT_3B(256'h022bfc1410001100022bfc14c062026a022bfc141000110002500014c0601010),
    .INIT_3C(256'h022bfc11107206c4022bfc3a4f4207ac022bfc1d10a207ef022bfc2500001010),
    .INIT_3D(256'h022bfc2055d01101022bfc01a0001080022bfc25000206c4022bfc111302077a),
    .INIT_3E(256'h022bfc0110401004022bfc3900001100022bfc204d320803022bfc09006207d8),
    .INIT_3F(256'h022bfc04a00207ba022bfc364fc20246022bfc19101207ba022bfc204c5207ef),
    .INIT_40(256'h022bfc19201207ba022bfc2055a20258022bfc204f1207ba022bfc001002024f),
    .INIT_41(256'h022bfc2255a206c4022bfc0110d2077a022bfc25000206c4022bfc364f720261),
    .INIT_42(256'h022bfc2255a01014022bfc0115f01100022bfc2255a20803022bfc0112020280),
    .INIT_43(256'h022bfc2255a207d8022bfc0113101101022bfc2255a010c0022bfc0113e207ef),
    .INIT_44(256'h022bfc2255a2026a022bfc0113001100022bfc2255a01014022bfc01133207ba),
    .INIT_45(256'h022bfc2255a0b002022bfc01132207ef022bfc2255a01014022bfc0113101100),
    .INIT_46(256'h022bfc2255a206c4022bfc01134207ac022bfc2255a32173022bfc011331d002),
    .INIT_47(256'h022bfc2255a206c4022bfc011362077a022bfc2255a206c4022bfc011352077a),
    .INIT_48(256'h022bfc2255a20803022bfc01138207d8022bfc2255a01101022bfc0113701080),
    .INIT_49(256'h022bfc2255a207c0022bfc01141207ef022bfc2255a01008022bfc0113901100),
    .INIT_4A(256'h022bfc2255a207c0022bfc011432024f022bfc2255a207c0022bfc0114220246),
    .INIT_4B(256'h022bfc2255a206c4022bfc0114520261022bfc2255a207c0022bfc0114420258),
    .INIT_4C(256'h022bfc2255a206c4022bfc011472077a022bfc2255a206c4022bfc011462077a),
    .INIT_4D(256'h022bfc2255a01018022bfc0114901100022bfc2255a20803022bfc0114820280),
    .INIT_4E(256'h022bfc2255a207d8022bfc0114b01101022bfc2255a010c0022bfc0114a207ef),
    .INIT_4F(256'h022bfc2255a2026a022bfc0114d01100022bfc2255a01018022bfc0114c207c0),
    .INIT_50(256'h022bfc2255a0b002022bfc0114f207ef022bfc2255a01018022bfc0114e01100),
    .INIT_51(256'h022bfc2255a206c4022bfc01151207ac022bfc2255a32173022bfc011501d003),
    .INIT_52(256'h022bfc2255a206c4022bfc011532077a022bfc2255a206c4022bfc011522077a),
    .INIT_53(256'h022bfc2255a01101022bfc0115501080022bfc2255a206c4022bfc011542077a),
    .INIT_54(256'h022bfc2255a0100c022bfc0115701100022bfc2255a20803022bfc01156207d8),
    .INIT_55(256'h022bfc2255a207ca022bfc0115920246022bfc2255a207ca022bfc01158207ef),
    .INIT_56(256'h022bfc2d106207ca022bfc2056120258022bfc2255a207ca022bfc0115a2024f),
    .INIT_57(256'h022bfc3655d206c4022bfc0d0202077a022bfc0900d206c4022bfc2500020261),
    .INIT_58(256'h022bfc36561206c4022bfc0d0102077a022bfc0900d206c4022bfc250002077a),
    .INIT_59(256'h022bfc250000101c022bfc0306001100022bfc0900020803022bfc2500020280),
    .INIT_5A(256'h022bfc09013207d8022bfc2500001101022bfc0309f010c0022bfc09000207ef),
    .INIT_5B(256'h022bfc031602026a022bfc0010001100022bfc250000101c022bfc03007207ca),
    .INIT_5C(256'h022bfc20530206d1022bfc2d100207ef022bfc041000101c022bfc2056801100),
    .INIT_5D(256'h022bfc204df207ba022bfc20565206d1022bfc20508207ba022bfc2052a206ce),
    .INIT_5E(256'h022bfc0319f32187022bfc001001d002022bfc250000b002022bfc20506206ce),
    .INIT_5F(256'h022bfc2054a206ce022bfc2d100207c0022bfc04100206d1022bfc20565207c0),
    .INIT_60(256'h022bfc1d001207ca022bfc0b03232187022bfc205081d003022bfc2052a0b002),
    .INIT_61(256'h022bfc20506202ba022bfc204df206ce022bfc20568207ca022bfc325a4206d1),
    .INIT_62(256'h022bfc2050832191022bfc2052a1d002022bfc2054a0b002022bfc25000202c3),
    .INIT_63(256'h022bfc2500032191022bfc205061d003022bfc204df0b002022bfc01002202cc),
    .INIT_64(256'h022bfc0410001002022bfc205652b02e022bfc0319f20780022bfc00100202d5),
    .INIT_65(256'h022bfc2059001002022bfc010002d010022bfc2500001002022bfc2d1002d00f),
    .INIT_66(256'h022bfc2052a20851022bfc2054a2b02e022bfc2d1032084d022bfc0b1322d011),
    .INIT_67(256'h022bfc325a41d002022bfc1d0010b002022bfc0b0322d00f022bfc2050801002),
    .INIT_68(256'h022bfc250002d010022bfc2050601002022bfc204df20855022bfc01040321aa),
    .INIT_69(256'h022bfc2500020859022bfc20506321aa022bfc204df1d003022bfc010200b002),
    .INIT_6A(256'h022bfc205422b02e022bfc325af2084d022bfc1d0002d011022bfc2056801002),
    .INIT_6B(256'h022bfc205360b002022bfc250002d00f022bfc2050801002022bfc2050c20851),
    .INIT_6C(256'h022bfc2050801002022bfc2054020855022bfc2054a321bb022bfc225ac1d002),
    .INIT_6D(256'h022bfc2057f321bb022bfc205061d003022bfc204e00b002022bfc00c302d010),
    .INIT_6E(256'h022bfc20508207ac022bfc205362d011022bfc2054801002022bfc2057320859),
    .INIT_6F(256'h022bfc2500020280022bfc20506206c4022bfc204e020227022bfc0bc3a2021d),
    .INIT_70(256'h022bfc2051201100022bfc2050820275022bfc2053001100022bfc2053e01010),
    .INIT_71(256'h022bfc0bc0520280022bfc204e0207ba022bfc0bc06207ef022bfc2051201010),
    .INIT_72(256'h022bfc2050601100022bfc204e020275022bfc0bc0401100022bfc204e001014),
    .INIT_73(256'h022bfc205081d002022bfc205280b002022bfc2054c207ef022bfc2061601014),
    .INIT_74(256'h022bfc2062801018022bfc3a5d520280022bfc0d504207c0022bfc09502321e4),
    .INIT_75(256'h022bfc09e1e01018022bfc09d1d01100022bfc09c1c20275022bfc225ec01100),
    .INIT_76(256'h022bfc14b06321e4022bfc14b061d003022bfc0bb130b002022bfc09f1f207ef),
    .INIT_77(256'h022bfc13f0001100022bfc13e000101c022bfc13d0020280022bfc10cb0207ca),
    .INIT_78(256'h022bfc2fc34207ef022bfc2fd350101c022bfc2fe3601100022bfc2ff3b20275),
    .INIT_79(256'h022bfc204e00300f022bfc0bc3609001022bfc204e02b04e022bfc0bc3b2021d),
    .INIT_7A(256'h022bfc204e00d002022bfc0bc3409002022bfc204e03220b022bfc0bc351d001),
    .INIT_7B(256'h022bfc205082b40f022bfc205282b20f022bfc2052a20780022bfc20506321fc),
    .INIT_7C(256'h022bfc2260a2b10f022bfc206282b08f022bfc3a5f42b04f022bfc0d5042b80f),
    .INIT_7D(256'h022bfc0bf3b2d010022bfc0be360101c022bfc0bd352d010022bfc0bc34010e0),
    .INIT_7E(256'h022bfc204532200a022bfc2049d205a8022bfc01b002057a022bfc01a0401002),
    .INIT_7F(256'h022bfc204531d002022bfc09e070b002022bfc2045320294022bfc09f072028b),
    .INITP_00(256'h23695ff88b272931c78a2eec66c1f6657667c8e7f4cbf9effd4ac7d9f97771f4),
    .INITP_01(256'h586a7aee754b08aa799e0fce5d4a74ebca0eb6f5020fe369e3677af2119fed8c),
    .INITP_02(256'h98112cffc5ae9c42f22ab244400c97454b97844743bb90d3f8d152899ed19a01),
    .INITP_03(256'h311854ae3c1ef6830b24a03c8bc90fc6a53b90619af81905edb5fc28aa9e9d31),
    .INITP_04(256'h1be09ae200c6b6a0a922bd2d0709023c9fb9ad01b49a8323a765b1b113cd81a4),
    .INITP_05(256'h23f0e443411e320fe544512c17d7e50f0850d80d96fd512397ed126072fc28ef),
    .INITP_06(256'h57a007bb7ece6eee748cbcb3c5c6fb61002d33e07c586618b5a2c157e7ff1708),
    .INITP_07(256'hf2fe46d2c3da5a57dd74fa70ea6df4f671d371da30af8ba8b50205b5100c8310),
    .INITP_08(256'he35ce3dde3ca654be54069cf6ed569dde64ce1c1696bf4c1e3c1fae8c140c879),
    .INITP_09(256'h6e6ee877e66ae1fde872f4e2e366e37ce3f7686a68fe686068e16152f4c5e8c9),
    .INITP_0A(256'hfc654e767dddeae7eae2eaf8e7f6f461e8ece379e3e4e3fee37265f7e5fbe8ef),
    .INITP_0B(256'h5778de41ccecfc77cd46eee97f75dfd947f377c3cff169537761c2f8fce44e7c),
    .INITP_0C(256'h474b73ef7b4f6add4ee5fae75250c8fef4e1caece1fcd3f5764e585c44e3fb6d),
    .INITP_0D(256'hf8f5c9fc64ed4ec454e14bc0ef45d37172eeefe3d2d4ce51edf9d8e6e0f55a52),
    .INITP_0E(256'hf0d6dedaffe8c549fd784acf7cc26d4b78f6d4667dceeac77a4c7f7bff6c7be5),
    .INITP_0F(256'h78e9e2cffef5d6617e51c06bc5685de4f36deb78ccf6c7685c6b56e6605251e2),
