`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6576)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpIW7IlOaVi4Gc9uJjkE4D1tIJkwlSaZnRXnKIleWYEAJhCJPcVhaBFv2D
8juyufAPDrKCwru0h6czlVo1YFubsjOw4JbXvtllvl1SLxgskzj/T2OD08JhwDw2hWK+jkudxUNv
u0SA47oC1ER2f0gqFtBe3YvAO/Jl9KsvzjRczP3ibH4/TImffz2apDUv3UAlJziYyU5X82Y5zDRw
ByxMvQ6n3ZwgvPhqmFxL1d9Yn1t2t2OeFfYe+hfzDBndwd60UciVi6rObkL4HhBSVkd9SIGw9QYr
RRozRFiFNrCI28aFqwNb8W49Ee6Mx8dIia3xE5RuaPKfWz0MBwartSRin3/FG/YGn498Rq/R+Sch
eDus70eLfMql/IOPWVUdlLu4m3SuDk0vQtcmQilZVWavxYFN2r1Zi7+6kzxBDCyKooa5Z5RXdO0n
EOrp5680odf5vcse/APoQzc0F6MXsJTwIUVTC96hNHw92JjLUzZX2h/NHdCZAYxIW75rxN7Smb7J
NF4E+/zneX/Z9bC9rzcCZSzMAN0RGkCaGofioR872zua20Zr++phsTVXXxkeWCBIzE1PY9+hBse9
r1mFtpBbhZ68PY/fZ59v7wdVy0b053u8m9W1CTLeAh8H7Gd1J0yh4MhVoaofdVFYPKVYU2SXUCG0
tck06/dfhvLdFIoBDM1fsviPX4Ts82ZT3F6rOJULFHPT5OTzD9FjL/+9IbKgqiEP1xRllCrVxxBb
iuHEJWrAxJGPiLIhUDRpIBgPZCjA0LT8AqG1ZnNLR47aJa1z8lAsN6zdE5H2HBV3c4EV/+2fEh2Q
Nw54HkvFBziQ2e07Qe6hnk0Z/aZ+8atCE9nTR64KcpiPUY+dcg5cTtXWIOrqwtOHBnKhZJYfCP7o
/pFGbC4XihQKi4YrrkMssv1q+jUbOfqG0zDDUL34x6zdPPbyAYVmyq7CL0X7hSjD86owt/4LiRAl
fQpAI+HyIFyHVmfhCcQ1YS+G9EB13h6jE/x8UZh/cE5r/SnLKIDHLUl+VL86ymiX0x5QecKAFGad
BIZhhhqAnXOaTwdC2p4iQtQKTx8LvE4ZHgBNkFBv24G7JT5ijJxxAVu8k/9bu/zpZ2zC2Tl+uzXF
KFmclPOoq5T6PSQDG7dY3w0+pmxWSxJkZewFuVpB1w0nFbjV6h8IjnWT/KTZiPtI2adiJP2MMc52
MMR3hOhAJ8870Kconwwghrc1IHNenUQdvW8Y6PSxGuSMcroAtAkNwrIdMnqCpq9CsOW8LFTMYUVb
jIoaLAyhWPaWf1eRRBU3IZglPaxikRRMgCXucfAZM0nNh3D/7NdMQTLq41p3LiVeQI06R1Wvw11S
dpt2itQcx/2V1m6PJMjx5XVbG5jL0Hqatuw0Xazx0mD6iHKubJI0H+Th+l4gY0NUpy05XuXjZtGT
rqhk4FKmUyfMM9BOrBEWPzRfMtxNEgbbdHGL8U6QhRBYMzfRceQoO17t8k493rQRaLAo+NsUcqLY
ad+CjHKr1XleUuzUw5/Mde275z3oj9n9Ikr2h2BtaLay2Ql+dfdxOx8JpixMjraI7DZbvb2atRgv
wQcEiEsaEHLR8pI96qnatFXZ6A1Yk0t4BoHPIBuxfg1/pDWLt+9GJv/z7SMIiTJ7wHS85nQHV/AN
38TehozlGl7pwMYBHS0twV0QiqUNtUUlG/fGpOhRdeqMxgoO2GgUihqTkV3fDRqUQG4l1Aha8vnn
97shCaWAEkPCU0wR4U1NuMwgfHzWFXLBAAZMQAkWfdburlmk8nDLU8ae0JdYr7ukUt1CdDR76oUz
hwfhaN+PZDB0cf5utGtXcmsgYRtTq56QTXrcbiTYS0DtODB3h8oFBrOZELPIWBqq7Ekac6Y2npuU
q7yvjZ0HyDLJopnGsR8pWXWcmYIccoOlN90VhOIjtH8lyf/LhWhNTBIGGy7sEUPFjbn3U3BX27/a
Bz6UEC/MKBbxjrZSrFIUwLkjhIYGJB41Zc/LgDLBG5bPC7Gz+idEVsR4CLcHRUcYEh3b6OqvLTnH
yMcDOlz4zqanPrIqBGR69c8gb1rrhnGtaDM0Bfhs7lgF30C783I3hFXRgF0rmYmfpn2ZimwJp037
HprXU7tdez4tzkyfYPzKJ0buCw+ImINGuuxqOUUhh6TjwKxzuat5JBqeJZEZNlxJ658qpbI9ncRE
shGvkdsBEzgy0vqvMN06O6OS2lbOTtHxXFN/9Nmd4XHeA2y9qTYGvctI7IDmi73Lee+ZbpD8iAgO
iUfvT/XAKuT7OnSfJz2LtacAwToprLk4p5evBxyi2d5o8uEXJALexoe4fe0cxG8ltUZf8jkUOpok
Lj+1ddBhSf2VXajtWIct/SQ2VbbRIlKrpVQx4G7FsaRNb2e6HcCkkkhCdgwzJtL8VVn8sYmXf1br
cqVMCewBwP9el9FroeGlxAZTD68/rTF49YJ7zDjSU7WFop3IThTv7nmHLECvXqsVOFjhjShsgTfG
2dCh36bF0mVuY6SNoOx5uNMzl4n8VhENfwUYSvjs/uCposYCY0Y8BGpQ2g05C77jjz3wIWGt/kzx
N2qe5AcVdOhERPvRh7hTg8AtOjEHtITMEgwa5yKY226uhEd4jMOWRHCyxHjO5Ilb9EOF1Fn/HC0z
sBJ+uDmJSkKoeSKDYizJ2XS0CT9CXJi/vSXgeBib+DP0IlETFU5yuUWR+pv+NOFgNGxz9oulhWCM
23oPCp4Nw/vQw0Csbt02RAI3AJHmmRqa+5Yblh78yRe+GO2oL1rVtY18XkJteozyQ3eB2/W79g2c
jfEH5OsVCAInDOHMPa1SncllduiOe6oC+ChYPOSkyQgPvZC3iIGZjj/r/ivzzBq8Yovq+Dp26D6u
Gwjw2/kzmx9J0+j1xgBqbFPLI5njx4TWIUfdHWuRy3p0ews1csa8NDKDmxMAvUmdvTA4BYbhBku2
K8xCNIPBphQOdD6H9P6ZJX7h0fcrZ5zYTVE2FXoKtbUKVz06dc2qNYxVdmmFR+W0bByyqwcTcG6z
WQ9URaACl/jD0DGZDR93kJ4oLxHzfZYh2WTSKNKl8DovuYpmogp2RmOHEIt9rFpCi39qiySpnLWW
lnfp3AiA+uojwRtV+deJNEQjYURVG/F3EZ7XS5dFro7idpemWXkybO00y6gTePChRaxiGGy1XqO9
00a0pnQ9778msVN+oqkyYF6Fc5tYaScjU5qtNnjPfcn2JZYyPd/2bDzXSvhQhqGTVYg3+K5teqW1
0PYZf/p01aNfWA4kDWgY+VkTaX0RBtxC7JV7GmbB9YXLN+UHYrqRgHOTzGnEe1e7faYwSLhjVdrR
auUrlyaQ9qjLvfGLWoW+F9VA10BXMfk6FmHPXwMCnYNNr3uqS8+8KQvu8l0PXPllaqF0h4KWqjSU
h6TrV3WDwCYAIP90BmW5qn2vb9fd2hOJ487sI32iuQHEt78dSY2lUt0mLToTQC87WRXwP2ekcg/I
QZz50q3NJux2idSStA+pXe/103YCez1F97az92FzJOV8ZJhUxeU6jzOkP4nJvTbjQCwjkDkutTzY
H5QAdKfMLdgZ3X1x1dK8O7mVU9tQfNs1X1iec+vS3hFVC3GlGdfAIWMhIu41f8+eQdr2CL4MiLNf
9T3YA2UJ5Npq/tL2eEzDK6NwSR/n7EaHeGOQefpBBWOjfYe23Qx4fPLrqgnVoIK47tBD2LK3Lp37
G6r6ayaW7C09YAw0r0e6v6/WWwHDMqMweuvq2G9VUDAEmP0pfQqsvosfW6SXc3pHMDJ5ApkzH0vv
68QJ2SV8cVy7p3HiYpKELKHXk2vdP73DVBGZrg59NCUg08kIvCnmZEZp7L8mQzYmBFRzyvuVejm9
Qr/8rQat3mCeo7E90zCILlu1bQ4CpyFrodxIeghpJ8gd2At9lj6X7KpoKIma7vTXj93Gpb1xB2MW
TlLt9QNqQIf0qtwHp6+D9CgR9Ushci7DRw8H5sB803kjYALaY8iFQfmK+RdOTWnUQRDO/COnptJL
UyqaFyMYHQjqVWy+t4nVpZrjPVWvayueJcjzpuii1UzEsqDScJYF/lJjE5tUSe97dinop3Ic+u9A
VoEbncHnqeiIUWFCRawXgBUn5JWv7T0nQcNz6dG2IgUj2cEGLIfJuTutvrgTn+K6rNWpiae99DiD
C1B6mhxwMlNbNhmM53nmC9oUgbqaPjzbUfN6aFkY27LE52BuxjJJfDyW4BcRSwOYi8ZWM4/AX+bT
Xk4rW5LA+aWlEcQFL45N1iqS5eBY/k+0QHfP5vhmNzIxCgQ14+iCsKgTtNGgB+Bzti7hsPJ6HhJ3
7qR+LokeATDAACXCWRu3uz9AnsgteF2Y8MlDBkRDNbY7/v7Guzr4XbGkPuLrb2up20IsY8q/W5kn
R6wN5k6ykYzvczwQvsc+v37VldF1T1vhkcK34GPp6pYjLERN3TZaeC6enJ06PeQD7ss4kacwUZx7
rhNG/GxquQUvcisTKjSvdhwBcblx0m8SKCliD8zXMhfQZ1m59NM01owusaK7Yu/wD+wmduOD+c3T
f+GENO/aCek/QQyH5JUmLWEExmXUIYs9BVmBcyN8ltE8vasskM/e4A92PjfqPvPVU0DtavWWQoE+
++D3ks8YsK/BZWUHTHQJ7ZWJf9OzStpLIq9yw2VjX6JDowGvrt8enUf0I8F2NshdhjpzIN6BOjFv
MvhBwdhPGSxI3HaaB6QwrYCf3hsT9H7f4kmwvNoo8oXP0XEu1V2Yk1CbvDQE0O0Thkld7Gl+VDQq
39gpRBpwU8iR++kPvSJUo2m/PH2b36NDC8pUmMKybRsBeKT3L71rDK6c8KDENPALRcgHTD1zao/Q
Mqu1XxhBA5gdl4eDgdHNGk/nMZC801D01bcysiu9/yFbwsl7N37DmxyStdG7yJx9gtpmTUiw5PeG
H2i/AF4wUoA1qcIZXGz20CXcTyhm7HpF/Wez8bUq89BjQwMEiP9WmhxE8Vme9eSwXEEdhA2JvRyV
Hp5Fo/vSXd4BQZrqvd4XoMcWNx3LH6Q7+YMMLkZWMOay0g18X5XTtaHQhkqs3TtC0wEN6kXwlaAR
eICeD1s8uVQ/K92/gHika+rPdY34dDwyq81cMYclHq8XKRt0VFXuFP5uzRM4CBG7SvQRxVz8AFpq
2Hyb2c9dwjsfzfm5yN6L1SIsK7msb9PVfqBK8wdRNxoRpiD32q8eUH3QiPwS+8OmvfL8Ckdm+fde
FKs+wV3C3W8UnFfddtQsdg3fdNz+Tuq98behDnwXETGTB/k5rl0BiU0O1e8QslJ7Q5AEGF7NYDza
aFy9UQOi0msJxRDq1N/81yk9EyJ7Smhgdn37gd/KPMgBRfj+I1CCZKgUgDD7F48Qy5yyAOTCMgss
xv8tuyquYNv/MkTcw+PsvAVzfJBI9UBK/AOcjkfm3j3LRvwJisEBDIrBC+w62HQQy3dY6U9f+EGM
15RtD5v18bAni52pQcaiRHqb5i2uLcnJebZOw3qmiuZ/phtDbIIpwZh/YEo38xB8l3sFjjzCqE1f
2caFrzhr4YsEstuyTB5iZLQzC8ggBKtsPp7D69mdpWd3PwvZFaYP+XvU2vwWlFyB4Ixy9UEAdysX
UGNz/20Is7Nw4RHlXJMM+qrQcFTIKRWUaRhIlKGVb2DpM0AI711rkimbSn98JPTYbw9M6hZBensd
7e/w/a9jn1ZrDVeb3rsFmb2ONnpcNfmzBiPdQtqnq07w0IeKYxrRYDTR0+iqgEB2dBgUquqi0owY
qA8zbNKY7q1X/KGCzyZFH5FssCCnBNie+tRnAt8HkgG8AtckvJPoTfzGor5cm+3Mv6W4/7jFGnoe
LCPXvmxe9c+Qf1treNdQuCnpJ3AjvpEePG/6syFd87+1Yr33at33LP3lPUxTWk+RxESlcJJmjcFt
B47xGf90h+8B96T1aVGUYCNjKEsfUkVxybvNrpewpoZdlvtxUFSKsIw0S6LznceIXuuKFoqKGlZ1
lLo5y1IjzHMsPCHaxf4pH6dM9C7TGDRt9keWsRcI+LKUb1r6y7BML4qNnk1bYv50KZpWjgLHUT6i
nd4LVK2zg70VneftocVIL403bEp0DILrhyZU+6AwogCr96hKH7hhQlJ3s6fPcpgtC66sdrWKRCpm
T2iH4yhcgil4A6N5nSfq50p6IsSaZz5//POiZtCpOpQlyZ+pf56SewgYZyUi1ARXDYLd6W6Ylxek
Y7VBq++xquk1grbry9rG9qpjKJtlRm6NszPtKNt1WbINDWXQaUA94CzWfQLaDhYaxZRzeQfVrFUW
TERli0pSlCj4TvS8Y8e9c8n4WGOB8GrlkWXuXAqbFcC0CQ0fo3rc8u75vpGnDNkRR0XxVR9Hm8Gj
/grjYflFOmnaoHGS3BD7ZChX6oXbRoWqD6nfCl3gvOo4qcU6a/KD6RhBiEM4+yeoQbqFPwQ1tlA3
r3PIeZglttz4fqXBRjTPIym6Ypp7dbMRr2Qode9qGsRXBjUzbbNECaXS5NtpM1PKfQNOZtnAWvqX
9YIouPJXXgN3af1JIsbB5EdTKfcrF3/VjySS9zkCXL+ffpVD6qa82M5n0kYXsS6+a2nwzIeFRJaQ
gC8OafWRCMuqKF2hPViX+NGXKkKSkEJbz+/4jWq+TjIzp0gTht98p9ZGtr4PIng1igvK1UYuRDlJ
nWgsO0xqPztOo1dxHQ006P54hGhDH+LO804IlvQn7lrj5AszY4OuSBgn0HYhWNfm8YOaNCiH6Pon
IgS4Aq+v5PyUg2qVKuf2GEkiMIa6sSUngtqgGxCI3n4UeiKOkMQHup3djTaT9IccRcZ1xp6MzEFG
MmbqlmcuB7d1WNjt0mNdoVSdCtpnmlEjWMm0AkHVJgZZIGb0nK5bpC/x9fNwTXXscInDuPjRSpyS
q/xPcvOlev5ulH0Kl/21E5NaCLcVYG4Nz4nj9W31swSE+FpUdECu6GeyhyhkzPcmE8M5lPZm8RN3
yJISU/xh9K14M7WMby83MYRD21bw6sHQpkrMjthl7MczFa4S1Gwfe4oo/8unScpzHI8hLCcb2YjH
99N/IyOckkFWu7DlFal23gCtaJqXAvga73rQciiEq0bUGuwvoLu59uA1zmYNUPd9LVt2yBilLq9F
y1WkT8wCKEzntauvkWjgFKRY81KtoUOOmaxK+XoXBFWiybFjCM6N5ax2ZrRx9I2Vkvf5JMqzMBN6
jrxRbMGVNXnSl1Ho5pyCoq/rfXX/gT+WjVKlzqRhqCZsm+HPq2tRkBchrk0qtib64ohmg0xVnOo4
qH1aEZujlQLJ3c2w2pWLSRehKc8/wTH7Mywu+czZkbFKGJvf8m4EHU4/u7lr2gjJEefch5zsX9EY
uTb/Hj2cXKZADDqRWdstqywrEsNO83xALS3Nqzp4hEs0JQlO5/j1jMlSPjGI5eCNxVKaNHNdX3NN
xklndRo3VKlMV9MWVFLI0ofSzDVz4ruZiJDKz8i6t8EFjx/QyRc+gyNXbYGZlinXKg8Nr+4FHykL
g8SvmN2zXAYOIPz5fe13t1Kij1lMMjuXPLQ6AZoP7sFm/ABCZf++oTZgtLCOkQP0uvy0L21u1/GK
3Zx7B8U/soPQ84ORLrMejnKIVNZ2tTFEcvWcFLiUlkMEBwZtA2xW3f5WU/YTdVw03B1jtq7hA+Ik
4OKyP6091xLRpxxHj52FX7FKIwyw44uI+dZaRVIpj/Gs5XQ6K0kEzymtZFPQCcQL2SxusTUorfPO
A6FoTjQcuimVBuT/qbfb2//Wzw0xYOGr9btgACfKK/kbojSrvAvMMSbdxRXxHDw2pF1ic7WyEq4u
DKljrbvDZmvzc0bpQ37dFI+XA6GV50Lsysk0jf5+EGuSDlbD+DYlQFHrJJL6hrGO7b0xXwaTewbn
BLDt4VwbUWPYB2Gehz2Ey4l27vHA41AnPLUnZ+1qYoqKxXQW1qR6H0a+Ds08xQ4AHi7HIcdNmIIW
yHABcgDJywAktmU6rSmKqSGyc3h0EZnQU3sI8k9mOkzbcn8eCOc+/1kgu0YTe9W2cDtfCkDJNhUX
p2H+nIbcE4b8iMW5bwnSW81Wyg00Fl2RwMWgnwcRZILccAsE344uB0q8L6gx5GQrj4EeBmBSo+d5
2w7/iONYxtGwCJqxkIeajGub6hYvbjQENpK9TC8qzxEjGLaQNXfo0mc5GB3PRbRlrmAUEKGcicL6
vpM+5QttLZscEb6ewc2iAYoTaP1HDiXvi8IgjiTDW2jRUnpbP+K7cdqzAOgDKu92wvAC+0BEf+Be
qTkUqGCRhJ3wTw+ZnyXkPjPDS5CKAa+ijc/9UUdo2JzAidf3eqowROKMti3gNY8J51WmBQHf8L5o
a7J6sqLx2ZSdFKPjVDZgAD2YwQjcT7EQmjbrqVDQBN73bAiO2rS5LdZL7UUPcTym735VbNLtk3Rc
3NkFWDWXrLpuRAQuXTOU1rQCpt/BdCb+Kzd016OhoM38okfPR2pEWPPY+hP2naEFIa6mmxdSRXM8
7SlnwIRoP9KaDa3P+Ac8YbRWbVFjcNplhNl6Wp1uzqmZr5tc2071ueqSwifidLsBvQ96xOnp/eIQ
3NPXuLaD98M3uoNsSerj5PkhQdCibi0lOzq6x7KztEvqFi6JdQCQfYO0CqV8lxLI5j2OhgMac37q
ERJrRnrMNwsXKDmD3joP33gCOgO4MetvjPQGeHOB/AWNLKGWVoHj+swiyj9KwlHYEIU89uE5ZFlG
mZ2ECOBwmcqsW2Efbw1g24Y+2kYU
`pragma protect end_protected
