`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AbtYS1qx1XJQwcR3dK2m6fwJ/a7l5k36rhAN0/BjjLJRPMA822p2APcpp4urXF6tbFoVheprueT5
yQVh8aEvQg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ewCvhMrI444gvhrZL5UedycCqCiQi3V/vNjUJE7QxihIJczzMVLYm1Do7aLvyFzWqwr5e8O1wfyb
8jiY0NOjU/LVby2XBpZhZWio3i+CBycrjjg85VVtih8EPG+IXGxg1DV9xJAJK7UZGb/hOxReUvKl
WElSKN7ydE3n7vtHTWg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGNkk6nsSre4j//sB80wqoR7TZaeXiddvudeaZoREY4KICRbZG0SUkW2Rig3UgE+0fPqB0MJaVNE
4+SpGpMmCQ+uGH9njocLfUgRCC3cVD2Qw3a6FdHmnt9w9TO/UYsErwMwdcPkxrf+qVdcsgLiTeG4
ML39a/gbhALskzVron0Ad/Ga+sdixRx+OZCGskBMwckDsJ7TaSnRrKniRVT8hqeeNB5INEpMZpfk
aH47TPXjD2ZdnaZRPUla7vQ7VytXzHf9ikp4IverO50AxBZ0cog9P7NnOPQduwE3iBhhBmG+W5n2
EblFp+iP6F21UCJlGNuyMDS0nYgq/kM8KT+uqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TB7LY8yNOc6mHyZZUKvhqMOOyT0ldzV30WNMBQGZ+smXGgUrX8kzuWrijolM/1mGcZgwfkhGdMXb
SdEjhfYs6uYhUnLRP4BLcpGj1ljMYKUZTRBg0PjcQliL5AaoSb2H/DTgaycnzH1XfRviEWaUKNqE
ZVevI+zPtdsHejN5wRT+Ai6qXlIpeT+vI3zsLdBeOA5rBb1VO87DVvu8Gd2mFd5e7JjBff1TQh3U
OdJn+LhPGAT1bmysYUiFIIx6pE/v0VqBj5lW56zweJem0GYP/uU0Mn84yONLf6seq1GNk+k0l/Jo
vJx1croNrp782+PK2Ku4+GW1cOls5vPOqi31oQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PrBhLPxaq/q/OLPMW58IkJt5Hwr2qplpqVZq91e8U3ZxED6RHHvJMV2zzR36pMdLY5dwyfM9SVYe
HGBm+gFMs4I9r1el9KLC1Vjx/wwyNS2WoYjDnRjOGGo+sD4bMSdcJHhNVIVqo+VhOOT0g79jHuWj
dd5+Xep6tVRHss9ayck=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OjXmzsa5k96Yv3Eghykbt5VUlQDs2uQJjEilki55kJT1q0sjGMZHHvEMSfBUTR8cneKpM7Ous2nz
Pfw8N3gMAtANYPDdsQ2FWVhvua7JeW1WAbU1KNU2fodreJ0uBYXSnK3zuI91D+yLwAhZRWYySp79
K89nt9adiSJUq72gqg1VmCppQrU/5Y/h4V/V+WCJGFM+qTpQ+nJOLzr2aI2OC+41kRD4dtHLhXIt
4oTZx7ieCgpPg3pIQRXdCfYFuChVlZi2voUXZ1PKbkScZrdlsVkIAW2UiEeUsCQekFuYkNgGIHP0
2QOtwXq5z3lUEaH/qgiaTJpWDEIPEUxlxAjMuw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
4xoO1c+NqtrYkzaKKva5WUiBPBAvX5ZDv9gZG6cM2TVk4pyZGwxa8tPfwUDV3X4JepXH73t+eHHt
9TfBtbUn7/aCur4FOIs7Ew3WtzeaKgxfEtSFQM4l793hz5aLiC0jclb1H+T3bXqb71bF/REXtu3s
nGR3OBC9DBNNC+AjjWYEujLSCKGYtfsM2xbJAJsg3TVm3tt3/bg6AYniyygbhNZ3XMDHAVrctWmX
I4czC0ARtoSeKo1F/tG0Lji52av2udl0AcvMEwr6EZOKfYZkLgoC5W/Om+Uw5/iEBobM5lCOLgYK
xVqExrZxXCMLpG89d/9gjxvzfPaV9pgrfF2+Qw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J+ykBy4c2cFt5c0uQfHFxTcxdU1U/V3YIloigBDJHrY/jm3X1GW1Val9trwqRdX79detroxFZwdu
Wpq/vLPPFSLW6XzzGMUR3eKiBnm0h0kNPKfQmQDthOxq+4halnmf9/cBIwwk//F8JjzMhgLm0CLf
a0isFV43mKb4jbI0dF3+9tFUNlXwt/vSbrCs9UHe7xemalLkuTdsK+hWU0CiBdVYCveo2bheXy17
2MHdBMHmtBgXIWyZ3l5YvgIM1cEsnjmHOex4ytPV0GUoUBzpcIg38KVuxzdr2/ZZzMsU8+CwLkYQ
iAlUM+3fVJ7g3iff7vtcaPFuqCdyESqCtTVjpw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
n6KlfsfZRlFriW0+hYvfoK8g2QUKaJhv+j7+ATqBtJbN3ZHLiI4C5PCqyevgC5fhKq4UGo2gG3+c
Xw+Y6onnRga2Kn4rKiIV7qKgzMusoSNFAm78D09SSiYNQ4CtEZLr0uA1DsMMn3w7wYYiOVYUzSmE
ZeQcdi3qNlZ1Q97MJYQOGrH83eM0TEuOEdqtUj2gOQcFoCPPLyC3OFi022m0tVD/5Z2J/36SwgCX
Erb/tNDb3IkzdiT0AFiG+3WP1USP8F+zdXgsziqnN4Ewf518NsW5WVTw9l6Es3xmVyzebc6d17qg
oz+nKCcR9hyxI3t7ppyr7ZWRK9vw4c7Ij0d9Jg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2624)
`pragma protect data_block
B1RBLrjJ5ienBeH+s3hpIaXsHg4Qky61BuTVrHwgMJ1PVik0OXmq3Uyf1uvv0O1oXqA8jQP62/iS
xBZeSkLb0NOgN3a2JxYFRubjzOQW6sjwviYxJNwB87sP9icx/66Zl3vUC8jmBZGeytYLx7xqb+gI
WYMZD1acSB0Ld7uYCKol8YQZ0H6Gte5NNbHvmVwZIw55bSFxpJ9L5CygaWggZ8SygYiGpKhhtqMD
1flbXGWf3sdq1yaLXjamFVzzwUpx9/8jyuwM7rQUBVL4jyK96AqiBeKv3jFnHvJKrbmfeo4R1MoL
Eu3J709qJxBYLTH89MEfSwkz4WDzXly9q52FzDnsVA6hiePcnDDa3IvaKvEh22s53TxvTm7E/xXs
N47Ruox6cqiCHDsRrsuLWCVr6992ldpr/11COHBU2xmb1MHKzT5ZB4Atx9+TIB23SdMASFALBKbI
FytrUSF06JdN2z7dDAd/9saCKyI/FF0fNWyJ/IoXs9h2gvwGpO2h1+2qHFtjB1HPUn2zcfHCZKBt
UECuuyY8S0kY5apPJsclPRfkJgLPCf9y6EIZr0wcJDR0jaDsyVY+7PMxC7PgfqzybjF8F4WVvU1Y
yuJuXLNN01uf0uxadUllmcYCqZYWJDkKwtAgbycPOqQBFQEBaHvyzRo1E7sMq1E4ziaQqNVoF1Ak
9zbXOT6VvwhNlsK9N1DcpK0R3dO1YaIhyTEprYRlUFNdCAwud2kIXwLAeo1qVl/AOhPvQlqBBsdn
kcNB2DDv07pX2epMapa5+bePWLPw7i+VOmxYuYnhWPiPE+3AmMG3RxNdBW2jxQmKtkcwkTzy/IVE
p01WQQQNtDgXuW3hRbfjz/uasLi1s00LmPYjergm0ox+ZqCx4ujK+Kj2OoM/JwJwqvups1cKyzZ2
llKtB/nD+RK9IgG1/y6W+ooBINOK7Oob0nd3GR1e0D3ylofNohi1RzcZNYVoFnFyyLBVx7O/lIcF
zAPXvlPe4Zn6BpXukkHQ7RVJtbrCUfacUjSRgv2vp4jLhUAAyocd4zBrWsECWfR2jjqqz3IKv7jv
nZA3yKW0OgO/6antb5Fs1OpvwmP0x8a2Xd8eHKeASLWzt2pw8Qhpzihdop4irBtj7na8dd+n6N7K
7w+elI+O3YJ+rGvhvC0+oHt5dujBHS8qVjZpXUkembZnwAmcl3aYQm/rs5R5nu9UMktizXwZuGze
zMiYmCazww0h8+so6tH68w9KXQQ3PSaRleWF9JzZ07a0ahasTQFbUe60TxGkm/2f9Bqu/Fwjvlzz
T4jqy7qkjHk28+i+YEg253L3U+PyYz1NTLL+qxbTqhfVPd+2S45Ooht1eE1tbDywl9xDirDJOmjj
0yJ6L2vHa+6wT7ohCiOB6Opt70b/A8pGv54ergRVSHCnqVR2TWLWS7KQtbMIuRLzR+CUBKWuHMsE
JE4qedYbZe0OZ9ijoFUpWF39LKnXjbGfNOJE+Z7MqETXOlM9/sp9v97FPO3K7yWX4fHuldJitJkw
Oje6Fc42Mu42yoC7dxGconZ9g/j09Ng0tRdJ+DZ9qcBlivAQcHfPX3hTc0as2LTQKv/ZL2ow+th9
iexdssrEr41/loGoNuDMpv1kUUffFSqm4syl8zssc6JCBDtmnusx0ZIy3DiRX98MSMdhSDehouKI
BYayMOd65BmH8WUETPx/BDnWnQ5rUF3dsvRSWj0lYGGPHjVePt+odY//ztlrfE7Ch2hW9P0xN45o
DNLSJNLH2iNRDj3jsNryfO7MizYcNqHUPx93QPN8NYdOGQ+GfGWiQxubbRRUTrOjNnkpdgIKA+1z
VW21tmzbZMS/PQzqrKDMgrHVAl4MkGXcBP6lLloX1Fe4I3b2FZ8jLbjBY5iBB6F+7luOq4xADKbA
HF5TH37t6Ywjg4Svyk4nuRbP+bKZHXAGQPqc3z0PlzsE4UD/qKDcfYb2Nf00XsoVP+vTKiJy1XFe
4bThBt8uzr8SDg7y1J69Hnggy+sCIdGH7Nvi6ts1A5mGZJY4ZwX0iO/NI86uzSW/12VnGmMMegyj
cjzbrQAieGRighGSteKPO9xEhh2NW/BSHz8OgA0JGjAELmDPZaSeYQg7JkzQU0i8lBzm47x60bsb
jNdTbV2fsTlpLUJZ+E+0WMNy9xLoOP1gsJyWE7qDKxCh1ZXnlykC5fu1bN5YbrtuNYVQ6cd0QGCT
h+JOOOEANqvZxT0p9yLFnIEA6GHMnToSdgsWKDGGgtvEVgdBbwDoRgQkXK8Sf+Acbtk6ket80Sc5
V2aqP0FZS/LLk+rNVOkEbifPTlZ6U90CjI8u7sXe2Cnk2I2Lqx2MVa6xmCHxxpViVdBtkdw9ahaL
r6Lnej3D5PB02xAcr7SPAKRWMTeY+tG2rNn/sQJa1ItdjFBMWi0DNkbouOe8COyIm41R0mmpBEEf
YFQOSOUFUp0oskY+hEezIHZ8u7a59so96hs1/0DjCc0cIg2FjCWCJb1VUqICXLEoQhw3hf5Lf76h
a6mvMCIctaXB1KDpTHjcoyXVZa7Ko9JQKC0augh9s61RUyn/LP+LQpxP+ycc+KtDBgbewtaTcTrl
MJL++zLyU0pkB/tjVhRwT6G4h30u9m2Rb1a8/V0cgxk4na2OBKf24KxXRwUU07MI6lJJqJyBh2Su
wvlf1CvgFEgwpLn4qJa2TU29IeOTjk52kn6EGdUJZMZYq/pL9YZP4M58GIv8ofjRVYtQfgbBc19a
bUOTKpnNBrL0P0GoZ1ttcU2pcEr5YCgYNsx+22pOcbt9zAf10fyrKJ9jo2bd6mic2WCkruOE6lAm
7WQp4TAPQaHjuP7QbiFHtyoKBETfn2ux3cog2nE9duCZ8JeDzJljtxhunrjKIjvdYxD8qYpGPSXf
n6hg0Kqbiy3woUoHcCHgBNB9COo3DO83/43pxQ0gVp2ZoUZrexb60dMD53YNsx/Yq2vosUiW8Q8P
xTKeIMpQ40L4kUA4ei36orebjb5xAU6kzbPi8Q7TfSPtJv/Y6lIMeZZMKBhHqRiH2Z0WKi/pRvEs
VDk/qhfDgMvBfH+PvJmaWBsx7JOEO3HHV40Ztls1SC93Ec8vd35xfjWHbIWho9Uizpm7JYqC7iSF
vi1+bFTzOPQuF11McADQPPbFvgktwevFhbinGwb2Z3FosqMpSLmutOwu+uthpy3ZwvEuGTiq41K9
N8KhiNWc5jhw15oYoXhH4fmAFSkkh9mwlisARn/ezEwqqaCOGtKM1Sx3syRO/JwjDX6NM/TAF1/h
yI7EMPHFLcF5fvUp1oo/xp7eUGCd8Jwizeh6C7NCfwF6yg1JZoiNri26MtSqyUu6feZDErGilp3A
uyO8ADxw0TECQfm2mMeO9l9MbGRJTDmfRlLP8/SIgO5Aw6wifcuV9+PHCVh1O088lcdZeDPRxYGz
PwyRRIaXUbl9Gt4Zpf9EMdTZZ0s91yr7O6aOCA2BdBAPPz4F0U59HlQLUklC5le/W+OQOGl9g/Xq
Iis=
`pragma protect end_protected
