    .INIT_00(256'h00000006b202089d0000000b21a206e300000014b002200800000014a0020782),
    .INIT_01(256'h0000000b92f2b40f0000000b82e2b20f00000000140208ac0000002fb1a2013e),
    .INIT_02(256'h00000001b000100100000020a582f01e00000020a3a0100000000020a2e2b80f),
    .INIT_03(256'h0000000ba26206e900000014b002070900000014a0e207700000000ba252f032),
    .INIT_04(256'h00000014b002089d00000014a00206e300000014b002248100000014a00206e5),
    .INIT_05(256'h000000062b0010020000000b21d2b80f00000014b002b40f00000014a002b20f),
    .INIT_06(256'h00000014a002071d00000014b00224c200000014a00207700000002f21d2f032),
    .INIT_07(256'h00000014a000bc0a00000014b00206bd00000014a000bc0b00000014b00206e5),
    .INIT_08(256'h0000000ba270bc0800000014b00206bd00000014a000bc0900000014b00206bd),
    .INIT_09(256'h00000014b00206e300000014a00206bd00000014b000bc0700000014a00206bd),
    .INIT_0A(256'h00000006b202089d0000000b21c3242f00000014b000d00800000014a0009002),
    .INIT_0B(256'h00000001b000100000000001a002200800000025000207540000002fb1c01010),
    .INIT_0C(256'h00000014a000ba070000000d8ff2200800000014a00207820000000d1ff20754),
    .INIT_0D(256'h00000014b000be0b0000000daff0bd0a00000014a000bc090000000d9ff0bb08),
    .INIT_0E(256'h00000001a001d0c000000000200030f000000025000000e00000002fb2501f00),
    .INIT_0F(256'h00000014a042247c00000014a043244000000014a000d0800000000d1ff32440),
    .INIT_10(256'h00000014a04206a900000014a042f01400000014a040301f00000014a04000a0),
    .INIT_11(256'h00000020a4b0307f000000022a0000b000000014a04206a900000014a04206a9),
    .INIT_12(256'h00000000a80000e0000000250002f0150000002f2263e47c000000062b01d07b),
    .INIT_13(256'h00000014a060300300000014b00000f000000014a062f01300000000b9003003),
    .INIT_14(256'h00000014a062fe1200000014b002fd1100000014a062fc1000000014b00206a9),
    .INIT_15(256'h0000002500003f0100000014b002f01300000014a063646600000014b000df08),
    .INIT_16(256'h00000001b003647c00000001a001cab0000000003800bb02000000002100ba13),
    .INIT_17(256'h00000014a002ff0f0000000d2ff2fe0e000000033012fd0d000000032aa2fc0c),
    .INIT_18(256'h00000014b081df010000000daff03f0300000014a0014f000000000d3ff14e06),
    .INIT_19(256'h000000032cc0bb0200000001a000ba130000000038022479000000002103247c),
    .INIT_1A(256'h0000000d3ff2fc1000000014a0003e010000000d2ff3647c000000033021cab0),
    .INIT_1B(256'h000000002100b10500000014b080b0040000000daff2fe1200000014a002fd11),
    .INIT_1C(256'h000000033041ae20000000032f01ad1000000001a0018c00000000003800b206),
    .INIT_1D(256'h00000014a00034010000000d3ff0b40f00000014a0020b660000000d2ff3e47c),
    .INIT_1E(256'h00000025000209050000002fb272068e00000014b08209010000000daff2f40f),
    .INIT_1F(256'h00000001100207820000000100c20754000000008400100000000000950208ac),
    .INIT_20(256'h0000001900136192000000131000d040000000148080900f0000001490e22008),
    .INIT_21(256'h000000019ff3618d00000036a8a0d0800000001d1003619200000036a800d020),
    .INIT_22(256'h00000036a900d0400000000d50836189000000250000d080000000018ff0900e),
    .INIT_23(256'h000000250000d010000000018ff36183000000019ff0d0200000000110236186),
    .INIT_24(256'h000000000403249b000000001500d0040000003ea9c0900e0000001d10336180),
    .INIT_25(256'h00000014008030f00000001410e2b04e000000118012f00b000000018ff0901b),
    .INIT_26(256'h000000250000900d00000001104224810000000190f324aa0000003ea951d0e0),
    .INIT_27(256'h0000001b9041d04900000019828090060000000084036481000000009500d020),
    .INIT_28(256'h000000018ff20727000000019ff36481000000011021d0530000003eaa5324aa),
    .INIT_29(256'h00000014106206e90000000381f20709000000001802078b00000025000206e3),
    .INIT_2A(256'h00000014106206e30000001490020713000000141062248100000014900206e5),
    .INIT_2B(256'h00000036ab2010000000001d90f208ac0000000110220134000000149002089d),
    .INIT_2C(256'h00000025000207540000000110401000000000390002d0030000001d80c2f032),
    .INIT_2D(256'h0000000b30d201340000000b20c2089d00000020b4d220080000003700120782),
    .INIT_2E(256'h000000143000100000000014206207480000000ba0f010600000000b40e208ac),
    .INIT_2F(256'h0000000327f20754000000142080100000000014a002d003000000144002f032),
    .INIT_30(256'h0000001450e01e000000001450e01d0000000003403220080000000054020782),
    .INIT_31(256'h0000001470e2ff12000000007a02fe11000000036032fd10000000006a001f00),
    .INIT_32(256'h00000001e000b00f00000001d0020b66000000037032fd1e0000001470e01d01),
    .INIT_33(256'h0000001d6030300100000032af10b00f0000001d602324d4000000008201d0ff),
    .INIT_34(256'h0000001cd30221b400000001a0020918000000019002090100000032b182f00f),
    .INIT_35(256'h00000009f080901b00000032ade324dd0000001ce400d00400000036ad70900e),
    .INIT_36(256'h00000011d011d0e000000013a00030f0000000139002b04e000000108f02f00b),
    .INIT_37(256'h0000000be300b20600000001d000b10500000022ad30b00400000013e00324ef),
    .INIT_38(256'h000000108e003f0100000032ae80bf120000001cd500be110000000bf310bd10),
    .INIT_39(256'h00000022ae1324ef00000011d011ef2000000013a001ee10000000129f01cd00),
    .INIT_3A(256'h0000000b0022fd1000000003a0113f000000002f91113e000000002f81011d01),
    .INIT_3B(256'h000000370002089d0000002fa12224c800000004a002ff12000000140062fe11),
    .INIT_3C(256'h0000000b2372d1030000000be31010000000000bd30208ac0000002500020134),
    .INIT_3D(256'h0000001cf202200800000001f002078200000001a00207540000000190001000),
    .INIT_3E(256'h00000013a0001200000000129e036552000000108d01d00100000032afe0b01e),
    .INIT_3F(256'h0000000b23c2f81600000001f0020a7c00000022af70b51700000011f010b416),
    .INIT_40(256'h000000139000b519000000108200b41800000032b07042100000001cf502f917),
    .INIT_41(256'h00000001f000421000000022b002f91900000011f012f81800000013a0020a7c),
    .INIT_42(256'h000000139002f81a0000001180220a7c00000032b0f0b51b0000001cf300b41a),
    .INIT_43(256'h0000002f8100b51d00000022b080b41c00000011f0104210000000138002f91b),
    .INIT_44(256'h00000014006042100000000b0022f91d00000003a012f81c0000002f91120a7c),
    .INIT_45(256'h000000250002f21e00000037000012020000002fa123252300000004a000d202),
    .INIT_46(256'h000000018000b0320000000b237208180000000be312080b0000000bd3020820),
    .INIT_47(256'h0000001cf20324d400000001f001d00200000001a00324b6000000019001d001),
    .INIT_48(256'h00000013a0001204000000129e022593000000108d00502000000032b2620742),
    .INIT_49(256'h00000003ff00b1170000000bf390b01600000022b1f20c1c00000011f012f21e),
    .INIT_4A(256'h0000000b23c1f1ff00000001f001d0ff00000032b332f1150000001df002f014),
    .INIT_4B(256'h000000139002f014000000108200b11900000032b330b0180000001df023468e),
    .INIT_4C(256'h00000001f003468e00000022b2c1f1ff00000011f011d0ff00000013a002f115),
    .INIT_4D(256'h000000108202f11500000032b3c2f0140000001cf500b11b0000000b2380b01a),
    .INIT_4E(256'h00000022b350b01c00000011f013468e00000013a001f1ff000000139001d0ff),
    .INIT_4F(256'h000000118011d0ff00000032b442f1150000001cf302f01400000001f000b11d),
    .INIT_50(256'h00000022b3d1d00000000011f010b032000000138003468e000000139001f1ff),
    .INIT_51(256'h0000000b0022080b00000003a01208200000002f911209050000002f81036546),
    .INIT_52(256'h000000370001d0010000002fa120b03200000004a00208180000001400620847),
    .INIT_53(256'h000000096082074200000009508324d400000020b5f1d00200000025000324b6),
    .INIT_54(256'h000000096083655f000000095081d0080000002f605225930000002f504030df),
    .INIT_55(256'h00000009608206e300000009508207070000002f631207250000002f53020707),
    .INIT_56(256'h00000009608324b6000000095081d0010000002f6380b0320000002f537207f0),
    .INIT_57(256'h000000015f01d01000000025000225930000002f606050200000002f53c20742),
    .INIT_58(256'h0000002d60a207310000002d5092072b0000000110020703000000016073656c),
    .INIT_59(256'h00000020b4d1d001000000370010b03200000025000207f00000002d10b206e3),
    .INIT_5A(256'h0000002f834225930000000ba12050200000000b911207420000000b810324b6),
    .INIT_5B(256'h0000000bd372072b00000001200207030000002fa36365790000002f9351d020),
    .INIT_5C(256'h0000001a9400b03200000018830207f00000000b431206e30000000b33020731),
    .INIT_5D(256'h0000002f834030df00000011201207420000003ab7d324b60000001ba001d001),
    .INIT_5E(256'h00000032baf207030000001c2d0365860000002fa361d0400000002f93522593),
    .INIT_5F(256'h0000000ba36207f00000000b935206e30000000b8342073100000022b722072b),
    .INIT_60(256'h000000094082074200000001300324b6000000012001d0010000002f20f0b032),
    .INIT_61(256'h0000001b90036017000000188401d08000000032c15225930000001d401030df),
    .INIT_62(256'h00000013300206e3000000112012071b0000003ab902071f0000001ba0020725),
    .INIT_63(256'h00000022b83324b60000002fa361d0010000002f9350b0320000002f834207f0),
    .INIT_64(256'h0000002f30e207480000000ba36225930000000b935030df0000000b83420742),
    .INIT_65(256'h0000000b50d0b01e0000000b40c220080000002f80c207540000002f20d01008),
    .INIT_66(256'h0000002f40c0d0040000001440809002000000145083660b000000144061d004),
    .INIT_67(256'h000000145080be04000000146082067d0000000b60e206570000000b50d325f6),
    .INIT_68(256'h00000014608325a90000000b70f1ff320000000b60e1dedb0000002f50d0bf05),
    .INIT_69(256'h0000002f70e0120b0000000377f011bb0000001470001ed00000001460801f09),
    .INIT_6A(256'h000000047000112b0000001400601e400000000b00201f0a00000001700225ad),
    .INIT_6B(256'h0000000b4392df0a0000002500009d07000000370002062f0000002f70f0120c),
    .INIT_6C(256'h0000000b43c365b700000032be61ce100000001d4002dd08000000034f02de09),
    .INIT_6D(256'h0000001ba0011e010000001b900225ba00000018840365b7000000012001cf20),
    .INIT_6E(256'h0000002f9350b1170000002f8340b01600000011201225ad0000003abc013f00),
    .INIT_6F(256'h00000022bb51f1ff00000032be61d0ff0000001d2022f1150000002fa362f014),
    .INIT_70(256'h0000002f20f0d0ff0000000ba36012000000000b935206370000000b834325c6),
    .INIT_71(256'h0000001b9000b119000000188400b018000000194022f2200000000b43c14200),
    .INIT_72(256'h0000000b9351f1ff0000000b8341d0ff0000003ec152f1150000001ba002f014),
    .INIT_73(256'h000000033010d0ff00000000380012000000000b20f206370000000ba36325d2),
    .INIT_74(256'h000000148080b11b000000143060b01a000000148082f2210000001490e14200),
    .INIT_75(256'h000000149081f1ff000000148061d0ff0000002f30c2f115000000143082f014),
    .INIT_76(256'h000000142000d0ff00000014908012000000002f80d2063700000014808325de),
    .INIT_77(256'h000000013010b11d0000002f20e0b01c0000001420e2f2220000001420614200),
    .INIT_78(256'h0000002f30f1d0ff000000043002f115000000140062f0140000000b00201200),
    .INIT_79(256'h00000001200012000000000b4382063700000025000325eb000000370001f1ff),
    .INIT_7A(256'h0000003abf1208130000001ba002f2230000001b90014200000000188400d0ff),
    .INIT_7B(256'h0000002fa360b1210000002f9350b0200000002f834208180000001120120860),
    .INIT_7C(256'h0000000ba360b1230000000b935040100000000b8340b12200000022be804010),
    .INIT_7D(256'h000000188400504000000019402207420000000b438325f90000002f20f04010),
    .INIT_7E(256'h0000000b834207480000003ec15030bf0000001ba00207420000001b900225fb),
    .INIT_7F(256'h0000000b300190010000000b20f0b01f0000000ba362f03b0000000b9350b00e),
    .INITP_00(256'h08b88b3d902a13901191288a221d271ea0bc09af1716bbbe348c03843e04a012),
    .INITP_01(256'h9e0a9f13a7a1af17a6a10e228b83121a94a6bd853e8e37023e9b299ba8b80eb8),
    .INITP_02(256'h0d01141806a2a6bebd3b8c2a0cad87b700a79f1a2db9090a1d3e88888884931a),
    .INITP_03(256'h963915bbac9d363b8d3d87971ea338bca6ac2f8ea1128294aaa1a2ae253e9f30),
    .INITP_04(256'h1d0601a3279c3b9c1ab7a60cb889902a3882b99ba03c3d80a5bfa7bfb79f391e),
    .INITP_05(256'h942982b697b6b49b260134a9bd0a88b9ae8b00863b132299b92817bf12a69e8c),
    .INITP_06(256'h9a1b08943e23ad999b3b3b0789a02a9d0d26803f13002538bc9202b31c1f28b5),
    .INITP_07(256'h0da20603ba99962cb0313a30128b05bda02c2d88b31d268c97253b008ea93934),
    .INITP_08(256'ha6a3b42493151e08b6b83b33163e992005ab8101ac3010bd30231aa7ba070011),
    .INITP_09(256'h362535313e8e3ea7841602023fa394303906940c9925981399b93a863c1f9c83),
    .INITP_0A(256'hafa7aab30090afa58c8dae3c1014a2320483323327b52388b91baf143a809eb9),
    .INITP_0B(256'h3eba050e2e9aaaa793278e8a9fb986b8891eac2d9e2e310c31a93daa9499993f),
    .INITP_0C(256'h1b82aa2f11389fa3a102988aaaa4af0b9722b0043e218d98848fb138a0b18596),
    .INITP_0D(256'h1813263c3285b02d1b808d038b1bbab81db6ba9f9f8cb307059cac950c0aa431),
    .INITP_0E(256'h2802aa2d3686082302253000281da91182b9143abf98a1941f1c8b8c943d320a),
    .INITP_0F(256'hb01b3437893e99080b0d0c99b4ba08b934bc1335b51907169f89beb9a1b89d22),
