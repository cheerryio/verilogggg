`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hWPaokAJxPlgA9bHTYPq5SYL9v7ZAlnDYRWXqCQ44ybtRvru+5rFDTVwvZGQR5Vd4QOFfNEgcq5A
kvWw/tTeNw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
squNp31jU1/P7ULLjrTachISXBT7Khj0S0m8eMIyYoopREGdw39LoXRL7Fa3kwScG+x/bXQzyEYi
1ouwEorQbXJFNgNWFpJrH1StKC25vdRNNoRPGVV8TRg9uvHp426Vrg3LHu0TZ+YKz3WoNObQU0H+
7MmYZ97bIzM/HNriD1s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ty3IiW8wyOTmD9ghXL13QnmWw+sE6gQXaWJ7UhhJ+DaLCuGgs2OY636kmHlNGccpW6SvdjiyAKL5
WWH06pZrGEzH+39KPxg+W1XkFVSKVLlqwnn05B5OzK7VTt1AM0SgmqAdzm/exEiKzvoEskb2GFD3
YxAussA9bETNGCkD8kG6gVU3/zvxv6k13vLEfhBh0GWYe5c8ObaquBgYDuCCDaXdAsGO6FkXHeI9
v0pEnrunz5dQ+1UoLYhWSyRxxXwFjfiYt0W+p/u90Ng/EVoDqk3Y1xUbfM7mHEj+ta4DmsckUbom
L6KGuDHj9fMGFNag9x8Ap+BlvPqsblpK2vfTDw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NqKK6pqPPejPCx0uKTfcPVBOSc/iSai+D2/aLd8D/DyvrJ154xOVR8PSn8isM6iI4DK8bTj4iEHO
J1YS80LR5w8bVlxgWtihVWUAT5sziMJdTh8jkt3lgoCqxo7mPz6ysf77NG6Fj54F10fYH3b0nvDe
xAOc6Ddmi1YC2aFUOtmSebC0bEcVnE7ojCRlyOmvntCaY/DmYwkawZQjfuo3cod7PMgvpeXyKhd+
BJMb1Mgm2qhXtD654hURY3d1K8BP0p8nANhJiTiR6WFkMAB0jsWEpjaZCj85HI1//6BGTQE8teui
aqsno6jsbsXIMS5kxfb7H/Hbw2Njlv6vZPtTJA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L600lulbs/0HjmQDuA5MddORztkcCmciBM9cKvAo/JG2BweEmtl3uetrXhU1FMiM6OE6IR186g3s
mi8GWkYeiS9TIO1YNU+YBgJujagOCCTJprXqtXCbGToLBYKSIfmSynrp07BMxzYZih5+c6U8yOpe
0jv+v8JXGO12xqgUWfg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfW5lF4UVhGJ2N2czod8zZvPs8kMuOEFO6kJcZN7Qc88nL+QJ9IFO7L9YaWpKHy+gAqiHlnGPdFH
KDGb7GLX2nqX8h60Lde0lUZg320rfRZsfXNg23WGvWut/a7OPj8Fy3l3MiNwEbe8Vw/sIq4yaLcZ
DJBV6NrqfSBxKZOXNOd6Baccy0MEPtKdMBKJu9eAQ5tUSzJAPMoNURaUlyF9SUKkSga3S7A3Zv+e
4WUxUfMXZ4JqISIMh81Mce4Mljiy5h0UZZ8Q0LX/kl6pFoP+/Ed9nfOnTVoOvtewUe0rA/RFdPEF
vucUcS4L4GrKbku9Vhwo4WaSSrIV45X/ZFz4xw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAd9eoSMyk12JjT0BJQdJIAkopar8/IooD1ItvqO16zGSxMozSLM6tGQI2qULq5yHi+Z8H9WA52
7+yF85xvbZ0lJ0LpVLv2IHpVXgp+SQhQZMnPpGg/Dd4yWw9rba80uedrPM9QmIRNnCArZhYj0Ep2
jAhcBy648zDcHw2kobmEFJb3D5jj9L/IxL9yct0P7rPpv46r6/LYZb10zQSsDz5QKpCZkLFGvuXm
SFcF+zxvn+qy7BLY/MbAhjzfDazQBUGOc6zAQ6UHDS7XBEaLtZUbKrjk/2sXinGmjdxbvnRlfoQs
PxMohtBME+6s77Iq0A0ZPzykLz6uHbqCdAo0bA==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekXXFOqI2h6Z2daKQR4fv2JVpJQyDI2jNUZAAefKW0DIXlLVZdiXhHmwyBkelbYoIFN8RkPfaY/I
grgBUz0CTmQQs1tyu/krvHPBZ09y8/YQXs0w39vQCqX73g5hH79hcJQ+nmOel1MZx7ZlPRy1e5wM
hcN818AA68+dP12SvuSoC10GnEcWJN4NKy9i42v5mCQmR6ofE+HcaNaoGEtMCMX7kPXtPskUtpm6
YO3Jh52NZpPjgT0uiF0qvM7beF7BjIgmZY+qWlCfGZzhi4KFTsZF4D3k2lhKnc8KuCHV7M27/u71
bpieCLmaGmeQIYpIe3qPe/H5/mrjvoYgjkGNrA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y93mReaMf2axArLmrifshq8OQzoEZkJ6xlMdpV9/ZGAnIGfYjkQ8JS74RjyNsoWPcJ7EAQXYQ5ik
LrIunWb73GsnGEcDoTZPU2uH/HMPWP14Sx6WShAKe2Xz62GOorWbIiiUFUJ/fgu3GSz88yPbHt8I
Q8Yfq9WLQg+xGWWq5ogCtm2NG97+LPayotdBEx0VSstcfF39MvKSYKmfGlG2DUMCAyQzwn0F2mpR
JD6wnOBj13t3/0eF9NBX3UAZhx/hIx6s5b9yBnrixNlLn/aLDPyKNU+AIx6mLYXii2aCpvNaUlZP
E31mi3DcBcrgGtAGv9NvnaQZer/KvSS2ZeKFlg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 138736)
`pragma protect data_block
YAZO9t3rnTBw4qatOXwyCahs3fiyq/876fXZqyDwf+7hgFiHp+c2EDoHEPmq1A//rk9HUvTwg7d/
3Gf2g2OBNHxLYFpe/8SvfbnT2ApIzVcfVc6+ImCxpXOjae09k1G0QKbjpzJ0k9ugm+gl7x3i3Us3
FVlaNYbv3v7qKP/FXmOan6TbDrLOWh7Q42y3SUAf6fgQx2dks49khdoy2ftO/yUVcR2/TfUX5Kmn
qPhuo9iHsPywHZhVfHLYL5MBl3ieJIebbWqGW46WjT/DPYoxY42JmtW+2pC+M6r5T7Xw1XA5xDAU
Nis+b+CQ53bLTxzIrVeK66sT6y5Ca6SADlDZaR+GZLHNybrQiIa6m7dONqR0/UymFju2zNvwHDtF
01Wt9NyjmEVeM/XBetJQDmJOQ/2DsE4STGlzqSz27rM0GZMaVrR3A6DBZcjJAtYYx5F+eiSjc5k8
1gC5yr5aX8FRcda6RFgk1u4SkUPUYDygaJgndFokS9fqBl0c7eWFwZ1BZEs0DrZ1zd9kp1ewVmPb
7NWItnTY60kYoxdhAkf8amF65btSSLxu2w6XA6b2ZXECYpdA+6IworQUmldKB3E/VfsC8La0T5Re
dEC+K18u9sjYruG7ZMaoYWgpHWteZ7lqChfwqShpruz6iGRpf3uY5HL9d3K84JjkdmMQ62y7hRNx
JiolzZ3Wzkl2iONgiOEVBEPOYB/n1z81AFHnHFklCfJ3NaRMF/4UcfzCJjJ/PJ5XiqGodfF2cTOm
/s4rpSdUWD7U7JVGBSwOxOKHrIXRbjtyw3eajWmXAZMfbc9+zBlGx9X272BzDtJoxNuYeAN1cBDX
6GvvgD9zd1uB2ebi8DH0xSbIzVBFA2KVb50ABD5S9Tk+YyeZ+FZV6WN4gpuFC4MNhsXcxUL/Bu6+
3NJjf7/tt41y2jGBsTfoGuIFp6Pq+rmeUHjk/xVX9ZOguvgM6GXsdQuS7xbkUMJ12+poa7jTi+lx
0ImRMFgHM1md49mHXvvPdCHE0ejxCH2dKy6hJqCO+6TWiBl3F2Eej4a63tTC61TXVQpFCccc78hY
nxjqNnhiIG7n4p1tN9faViV8KkwHNpF2vx6AItu2DiKL5DTzdFprHZzDokfq5vJOyM0U/gFi3Egq
A12rml+vyuUICO2wn7MZb7E9Kz7akycJDMn8C5SuKgfwf9NDLLwi4Yb7PFTqXDsqYW/z51+JSGm7
/Y0iUxIKB+2d13bT8XVXrLxwLpqPOnre44GnDSEQ3+pSJ1gJ7C1IcuEqwi3oLbaqiJAU99+KAWcU
109o0YI5EOlpaVuK6II02+bz5CaEmkA0TF0zoBmm5xb3WnS1Hf0DEc/xBuOv1bBeSdqMWItXVZ6r
ludEmOyarR1r671SkCHexdwNzzB4u+CZ/G1t/laLsNre133xQSNsgFzu1a921/5DOnyuKqyzLSbm
Zdc7ZU29l7g/+kTHYhx06kkINeE1fe+nuM32E86bNdxj9PF6m86wmGoGzyZ6RZGxx3viCNZTxpvw
NinXvdhnKpVMzE7OoVDIbEUCzVjOuQOApV5ch8Mw3DM9u/DzZ2pP9Qxds/SDL5Jlx9IzkRmn9Zov
cPh1Vgm13PVHo5EQCs2byw9mVuZ7JrHxCBxAEooQSOgAJ8QILLrYCPwSnRaoyeMlOE1bcWXV4HPS
l/glb7rxeZn/E6FyvJlBZvqdxv//1V6mkg6xd0o3cxexBhifpDLrfl6lUIpgY0310limqQO1DIQe
hVd1YWuTJN1Zm+M2PpVa8I+hG7fpJ+kP7D4AiLC9NAtZ7tlNXwnjB8iQwfVo7Z3xj+wtarP17Eps
zIGWEUFCq49U5Ft7AGBg8p6qKyXl6s2n6VipJUDBLFYHrmUCDo4k2gMXp9MBbF0kF2iBDbzc46FY
MZ7WFLtXcrfGKC84bmqxgSvQn3ZEV7ydGND530xxZkrya9CAJ/v8KkmoyKpRvRD5woJGtN+o/l1b
idNl9a+skcZbnT8uONouW6KMF3vvECpiDNrsNSOQhWAh0yfGQ/Yl9Vq365bSMk9LVZXJGmI+meMM
a8lLSgsQTreJ7jhUPBL5FvgdfbqcoFdKmRYLWcAvQNq9TdbjYt6y6YmdajqcUwm7Lp33JYT0QMUR
NlwDnIJzdjBGH2ak0cj1px2EbHGHjGWIjo/7cz1DjJ78AhaAfX5MLyx2ff88UHXA7n95WUSr3Tfp
Pux1HzlG++eaDbDtAlgHpiu+4Pg+9Bl6byCCBJe9KyK8QIV/++RmMpkyAv/Hti/9ivOVm0GWKqcd
7JWxfLv2u+aK7v+DzXyEmBvqeZfKfjC3WuCX3cypeWkZXk3g6keH166fNzfQp4/a7SDCsoGNyLbr
Yrh4h+f57T7iGvBYdTau+e1HKWvWGqp6UqsuoqiCCxvN2gZZGCmevv2vv6+zx6ddQx5GKymL75W+
O+R4Za1bt+J5JIRHj2BLvwCo+tvm4kOy5TVbqHtvGA0aU3oVvFoKWEWSPcTlzS+UtX4uwHjQuVvo
J2eug24/k0LIyPqo+TW9/kZ0TpRu/wHgbiptq0rlk31cQeHoehQnMHCWx9l5fENVvG/JsY60Xjh5
diGajrzF7JqE8mV09v7cW3+0Al8fCqDHaNz+4LV9iUxbsZ9/o5e/ith12+Nkei5s7m3Ozy/gJrHP
N6RyUe/9sWX8qXPksdyTrTkzIDN7oPBKXUfCNFp2o14dPDzhNSyQxB6BOFa7e/MIv5vaKtPClK0+
GiM8kTJ1YqUtdg+YxXZJz2U9x56sIVvpDfMaTEMl3ZRK4o+cEFm5El6GKmfP0AboCo7SALYWP4/W
ziIA8Shv7RPKrVhE6z5X+vw4yTN5YvygnbylqeuewOPqpuCwYXR7kWI70nEkYbgQbWOQTJcMtnaB
J1bVf8oDv0t5zUxnUf7DzcRVbzDqLYLh0z9rDLAFbtWBfMKqVB9zCVlau+JOmxcMcGWmku5vQVHD
zPRKbHmndtukHacs3z5l1UMIicgTAJk/opYxavrVHfY1I+3UDXU847GFbbihv6E25KN4DCoQLpMn
Jf66P2zkw6ju46bGYrqnG+ioVGTrN6M3hoCsY68WCgFBDGlRE1Bb/EGFc2tupp7iGgcyxWc5NyaB
qzIQTko8T+e+Ir3t/VB10RLSeVtnaSEdn5yKEzNm1fP3/S1h0mesx2F4oHoiuWqUjNqqg3x5SLmZ
CpcagMMxQKxZO1xZMUWBppms4cIIL5YnIjQyKPNnyeBGnNQASy1t0KMxo4runUWlvbCeTUBIWKaP
cKCOxHB1r4XoPd/LDTjZq96M4H5UNbCe9Cs4u96PkK4nAR3rBXRtQO5ZoHpAhsLE4BhBF4aaEHVe
ulQBu5M8DxWs5eTd5EkWmg/xUcMsflnEB5riSO18RF9aq14G3BuQjTrrjV28bD7arkfAPo/T1a2Q
FSwVjmVoxsK8kPxdQkEUmJwU7Eqm0q7k072k/d3tHLlPzHdOMkgcqTrTNl2AKg4Inw2rFL4XYAP2
a3mpkqagm82dH70ctICfHPU3m3tP90xFB4wXLPktsHwSQQsT6MUj0if7QagGQ6uE7dgdXtw/XLZo
q7CQgjPgCOR19AVihxV2oeLv6Msza+4NKYt3tPv+ss2sJc3xOIM2TAXZPCCPmjVRbj+q4Fx/7b8w
8KRax1WPHtspDYXzZHuGZeIZ3ufPdDdaqo+QBWPgdhnyPOatFN5pDOWDfjiDl5jP8YErj58UzusQ
Yf52p7NthghPbc0UwCwG83bkR0uwBExAlAKPB8g6V2jvVPQX1rndPGDzvbt5CiSSeCsFcPNx7kx9
1zEYeW2fVFePBtAKrdbPAbt/cndPU8DnUXQao9U1FrmdqU4IgA/WuaR2A4GEb3y8e0+kvDWb8Sv8
20VnQs0/C/rcl8Uki+dV03dqMK5IdLNXdo3CBjsFYRULz+8LwiVDjsCc0DLI/Iy33Z5by62ylyT0
awP37hrbjH0ovFaQX/RNkScDGKhXuZM77zmiHU9Zz0Oopc5sOYrqA8WhN+2qqMOV3pClCsdw5Zx5
S9IXL/NUEJjEoBvAgDzYxAcuYMeBeBNdLrFk3ZFiJhZW+DZv/WGtpwkiyUYc3amz/kx/Lt88TZRU
Hhp/GnpVRiXtimkERBZJ3XMC5mwVNtlF005bbJp4areqBbZ52MysffzQe8ArPOA5FtSgP/R/ddd/
cftxmgpMjQ65wYDomnCzaA+lOciTxPTST6+gCZ+vzGbs/DAozUSGHKBr4KKNJ0FZdcMF5SDKDqiL
NfYeCJd4xDNrv1jyv0cTEBFp/QWyiHVkfzkYfQl7yMkrkwbSIoyk4f8oWX1enpoO12db52q8/2U+
L9Itg6tfupkZ9SOaP55/lWvNWtiflV/dr/cqZz56icomkML22W+lkF718fUcBBLFB2d2cKdNEqe/
ORZYSxiWDJTzeeTTSVNBTNsVTDuPLHyVYiwvtEteivqOGsRJfa0+09igW0IOAtsxjLwYappHR5sH
8oq6FL3I95y/Qqw2l7t40xwRfw8M2+Mgmwu7OGQYZmOikM37umkJK8n6Ez8CtvC5wrXS2XuRB98z
hOPbSt3bp+x4PlHXIE4/GmlPqC1HQdNYCe857QpgT+sLw2p9kkLHgecLMx5YBD7kuzkomVx1Tbt6
g8N/0+h1yR6aGdu7zkIM5Th1C/TGLKOFP40qGOhzipxtPu2Nl/7R9vyrveXhDlq83liuw3POxNOU
Li6W7XyBKbABGFRKyx5tj4+9mNbbauyX0r2upLW1+oSKDV8TMXRqAfd+lfdsTspz01Mms1iismbK
/d1Nz0aISoW4uq1rCB2AGaXJRDmCWwHg1ydIQBqN+t8futNs/ifrBjmoiNIbXtFENCGRaYaaJy/3
qdMIujV0KzvUTFrYs5OLZ6PNKv6EdE/x03VFogp63Qq9anQssXjq0euOybPSBckF78MufzP+b7LB
QWobXmc6NFv4zdGC+hp0tXVU1g2cky80jRne4cZXFLc+YFNxUiUKO4cciXqTe4lu48ucs+aBcY8g
wzATl5p4+4udKRruJCPSTB3OwoEphBqvp7kRivMxuhCbWAvmX/QtJ4E4g6nDvlWgs9lC+CK2hCXr
HdXb2S+D3TfVtpjEd6vafQ4C7dV5zHuLN2LirXZeB35ZV9s8LI9A+ldNiK+m0fUU9TZxpGc4uSUl
VJPGULCaWmLhUpdfDQnB7uaX2KXeMREpeQ440uLZg8RAk8U/bqiv+d7IMTvZTyAPo2mI11ew9VJa
Uj8oRNaYpf9C9nzAP3Y/StimrOhHtGGlKk+oQFeX+e/0CEquh47mpO2E3hwib8YDOewKkB7AxKOB
838N8EBiTOTxNBtp3OkW7Amf2JpwyWbbAVafXJd5oTos+imwCRD31kuj/uL6x4i9lcOaf1hD/8AH
iYV8tgOfNy6thISEhju6Qn9CyX+0gCT3kYfu3JjRbqMuaGfU5cs63C+QxSClrGrOX3IYWUXIwzUY
n/tuQa+TWmAVLE3xzmQDDCrCu05m2qZK0AKR7/hn/2GcdoUIEvH6DXs83CaoIs48f5c2gWcmoOqo
rWOf7e2ge6Fugl56t3G78/Uew91xfK8cAopeNpHaA4OpZjTgYKIzyqVFAm5iBKDWuCR0QAUiPjWW
EnwNLVGsyjHphMOJV0FrJi6sO9Uwa9s9LLcyRnQ3EON5Fx+mR936fpvYWPNl4dWfiqpKJNN64Pl6
Y4qXz3f61mWOuqJziRCDbiB8NuR5s5j5icQVOpig52Qa7uKKGRNyoD/+tv2wheqGAEiZ8rLmbi7x
fIyx54RrLcyzw9BzBehCyseYxbL9xyrMwMguuB3ZWUL2pKt7ruuqfYhSFP7CB/yvg+6zi/u6EuuM
e2AlMoLu8F1zhuIgEeUj/qw2bjwmbS//JE1X8oPd/+vKnc26QlFPl0UaZ7ErT+8QRgBlBxEWVwXq
nVeZ0iR9jOIyI61E2ZaRgZOlhnjT2ACG5xnyTxfZySQ7WISiW07QEnXjMy17PtPYPunO7WoXn4iq
V5wmLXoKml8Wu/FsMlzHP9fzFGMloJ8jIwsrL9/eFWuLV+Vf3T5L+9g5e/LWXajO/6YXiaCDzPMX
8Cj70v8a9emSaBjf2QYSTl9VVgLCBmg1a1SFiF1OJbDigKbIFAIOQ/GXEvXmm4cUjcipW04FG4gi
Fi29iicPEzw8pyr9shNPK81Fhq53vkHEI06g8BTctlA0GtsYq55ERXkSNe8teqoxHqrdYUD2TaIl
RucmeyAO0Vus702fkErNVY+OO5FTavDmS+mr/Bsb11ReyyGAn+5rhXdhQpn6VSRe5YRkIhfMIpFF
JsEW08vPcNsP9YkLaIHtwfutrwd00Ae2PlxPuYRxK9hwZWKVH1jVx9HefboOkJqELqq0efEUkLk3
CdinyOgl8qdqaBFmNJiMJ8ESMVwbiEG48391fcuOgqK7dKHkr0LWYX1N8Pd3prIBsxmc8sKMAzU5
8nvavKGmL5DDu1UY2Wjp78QOV7qe4TY7dLdJTQUEaPjyeZoDevRE0gGEX4SlLmrHw0WDFfjrEbbM
MSeLq7GMXa+nCGuZ60LN/MbhIJ5KLg0IxDfa0iQaweK1Df6zXnMelS6TRuPUmXvFq4EyXjgt3pbw
upHMHBKAtzphFnLUh1RsxfR+8PEfl4ag0RSmFpTIlLJHZhP4mOU08IeRCrcgFn55q75Y1xs0CYdg
8Tbfza9/0Uz+5R27u9/XTW52mBbIPsf/LjO5mrNEdlOCcZCLqjGfIRFBgVKKLWAkDfjg50SpYLTU
i6llBbO65zpd8I2VWPwFbyFF4IaztGvbHZVjlzh5hI3AnVRratBvJNIRrskUxrq6gVzjEQ8Vu5mu
KiebdB5VOlcTKkxu4vlDZbhUS7uDDx/OMgBvhH+syRPt5Tc+CX4YZmUILAu63GRlu7w0H71/HuHo
sHIaoHKRwaGrelWK6Sz299ieeBFgmcgkhifMSMP/1Blint1nhZXGdkQte52FmWxjuvLCJNI57o5y
pqRJMChHmjTeAEblLbAD5tiU0kCHZpEMU3lCgfSFV7Ph7XFeQC8SO3NlvbaI4aKJnKKrsXJXY0mZ
Fo4K4gjwZAz7pwdvV38/Ux4hkTw1sFQp8dB7wYHtWwDGATPcEdoll8SI4YDTqL/wY9JUHeM+Uapx
08UaBIOYRkXZcnud9KuYqh2ICfOJudm7mlP5/Q3xcutVMnhcSgUDV87JjnqARgXOTMFlhP59vcyp
AQT4dgiuWvHra6kP84Yd5/45evrast/+BWeZ1htKXvHblV8QW38UnZXEhNwcuMbcvfVH1YOUayKu
o7LFiLdkO/Py8tMjfjjzFlGOTXIi0LMko8q9ngg6xh8oTdR1Gp7kEaZhcIqI16LxSFwliXUB4vYL
OtNgNqLrC3TBHiUaC7RGRKYkY859iTe3tT02p9BTsDqKVt7lSiQLxOZqBSdgw1Vub37tUae2/t0j
USd6vcaKnOmjyulqyHlUVJzkrc4hlp7RlMVjtjTgmkglnoTVGf5odBrgP96NVdu8nfOJ9gXFt8DM
G/yOXz5ytjSZOPfyKqiA2QFfEmeip5UmnqVdLomxxNN5xoQBckVfcF2hXTAieoTLGeJ63jkldFbi
6EX9HqJy6jFOXkCaoiqk5W5DMOiWkh/mDz6u7H50ss2wRIxK3m+11rGd7ribtgR/3FYOwEPv0gd+
hOitSUjPWsfapN9aoYqlH2ZNBod2QKheomOVAZOPZaHAuV1EKKDf/0rnxyyJMlAmGXRAupVhlVah
VniTGeypzjcXja/7R5oRwmIkTB8jfZEkfcuEXXdlXN4BCLVQXdh14ju4dd5W9vZolGqjHTF6rQHB
4mFYWhH+qZSj0eRt/To/pqWzbvqUNcgC9gLGc0Yyn9HfvRRogzijoI0hlt3UsfKsF3XhlbiFlDFS
mQydmchCaUry8uqTD9JfZLzzP0ljd5zs5c6PyJqvUimgmw57wQWdCt9nZZU+d4f65tZNLMcKdIvE
GVMz/tMd9TvQXmMNtU/SenLwrMKqg24w1gO78JG10nxWti4+dGB1aVHwOPH1+NZZsmPsRtF6OdzR
358RKmfZN9ewflV8STkLnYvSXkh+6lg3+OWCmhcVdP9CSFOjKiLSf5DtwnDI4VvyrB46FN3EOQ/a
kUR1D1J8mh03zFONXliODoprLrJzOXM3qZW7spx76F0dmAhi+0Pzf9LLc9si60+P66hVCD2uQVjv
g0CFsl5wa0fDXzqP2ZHxqk179cA18ZX4ugicPj1nCkRUf/jwFnziLwG67BIPvDmzUyr/ovnHp+hu
aLfXUSenZulIvoiryqAWMNpeSyz4phxIhVipio9fLgjKbikkKnuu1VTcKl47+AUPC/Ea4wZeWr/0
qRxZ6Df5bKfX0kLABa2XeUup5CLCtttt+TOaZcA9f+1pKcmRPh9UeMCXKP62Gx9lnBlqZgDwK1x7
wqpdk0PWM7WMcQ8kwVtnkgp9R/pvGxllWKCyUVKbYhAWM4PuGjy4NdsVccautOCiDtpPiGIDnufp
7q6X7AxExIflrp9tuMwQ/yXfTi7U3bK4RdUQpFKDlvKq9M0xcOZKEmRafhASZdTME6sVdtcHCNTY
Rju0AbCP2u6UcA49KvapY7fg0zpqf237ZNTLTeOczSDomaTs1wz4VQDeYCclVxEb4ptq3lspSiCL
j2B35Bj7CCJ4QjVEp+2LHpXDQLxBqiXbnR1oaQTwFisauTuJkBXvMPv+o/7Skzb/gK515H8C2Xsx
RxSSVbacDQwukGVTg7HxBX+ypTP5lhdgz6k8NgWlb4vgU1NVGsQPtM5NK1CzVNHFtLeE2rdVfQHV
YKqtkxn9tT2Cban7CxRdTbxey2UwTcx127/LsNZXGDkClKe8Ezcf9N5IFlAc9++RELaHXq/2BWFo
GATV2az+avY44OK8VSpJx8iUgWqoESmw4iSO7sZXURHtqD967CU/+QH6yxHj0JK+nF5s1vdsxDCy
98po7zv6T1nCLpx+R5QekhmkvSJwo0wiAQVr7iCH64HZ55WX9oxwJlE3MnVXY+gbpwGrHB1XdFll
WYpxPg25kfzCFeROyCB9wUpdP2F+6hPooSVFfPcNmmLBtvkuu1Ozm/+JUKxSBUr4k3f8JL+Z0Oim
HnCZZdXZZLtSUParJC3JLXKggGlQRHIKqEoXWsyeAWE0KbM0sCF0rsQS167TBSFcP6A4CrcBghC7
XaITEFLDfDZ6xuiDqlVb5YCSQLUecIXx3CVjWKOivnu6rqcBfVIxze8NgmpILo0cYkqJCznutpsY
4BLnTnQXY8MGbejHjk80bHafEgJrejj6q8DkTerwq3GMa1DGH+orisuoT+R1uW5PtE9T9basSybO
IRcSoK7hNgSQ0S8zxOpBqeOVGprn1+CR0sS6eJnPMwyLEMKd8a5LOU5XWWZ4hb6eN6BilAbjvFmF
wCpBwIeetOHb0Yti59/GN1JqD9ihj+DI6aqRODLSAdwJz3RtZBgPUlEbFf/5Xet7qGN8ROMNaEso
ZXKi4Hj2mBUEfCszyTtDzf3sXXdlgE5RAzydFhhsdlLHgiW4JtPlOM6S20s/5Id8/7CEoh9XuoOK
WjQSqdYYxASiMm2AU2yE99cLMeqmtUKevsNsMCG0mO1My4FUrKrCoXO+ElbQ2VGU5fCp3tFMDNSV
yG6ESwjHRqFhlki31dQGrj/lLPJUHhI4YPV7aY0v2/2MgYvLWcSbvUMESPnhzwAp6q/3ooM4ABqf
Et+JA/MNrkidNBdlm5XfJJz/nRH7I+3JBnNUxNafsVgnGLeJTUTMdQv71j0osIGneMtpRKIZab7b
o4s3niGHGDhyujrr2gOyUUXkc0r2GkmoqvCH8YT2g4dl/9ToMfkUl/Qghhe72wz9Bvkd5e/E2Pji
8ef4vlrLP4lGQGgFfcRF0wrHO1EYpg4Pd8NYHQMJf2MeCN63yBCUIne72c4WJ9KCeHpDpBOoFoEU
B97wZm3g/uqfEKeFSzglXxyrWYQlc+d4niWhOm4RV6O+xNkJJMRIlqi5BZQ9yExxhr/Nz4tXytDf
DZ/sQtZnEXByY2g3pvoX1lO9oOR4rdpuigRPvieq0t4AQCy5kbj662pD/2L6KGV+BL4R3cltp2Ua
8QRqTGTV/1Y3zx/CWEsryqcf0i6ECCmfckPUf+w/XFOgXlwZQYfFqMP9abYv6jbQaKIXAMr4aXx1
9IoT1Ipg0/oiCyOSF09FLO7iPCyDkN9KW+JQeTyrlEHCjHosMpw7oWN0iDHJPX0Aq10cwW511Lvs
0CChnYcEWVQhB5/eIOKB8HL59aQjH4OLEGecSmVuEVXK+W2Ad31cBYiQazEB2B8xOgp2vL+/yByF
2MaxzdjNxTMryRSUGRpJeKJZbivxk258bsk7Ux8RfhVM/TF3bXKC0B0Ksup46QoG+RQ9lVRWqafF
1SV4YnU4XgB1xKlZBGr7JeuWo2Mydgok3RNcLpSY+i6BEjwPlM89Qxq7J2SoaKsNySu2B5OK+CxW
SCRq2stOWBT0BMD3pGyHCr4cKM+O44uOzKKCRClt2WagIT3gwlu6Hp6I0m37YMApe6fH/euoFzlz
qWtEzX3UdKplO6+orvruX6Gem16c8VEIVZHQn3GJPXnQQPPiOyuHU5T5pWcDcXFe7c1FLy8fmgfk
7ZORV3/u5pK7mD6rCbDjdoB1FeQOR/NOEORYtz6txj5Mjejrcd8L1CQroVkrD+qy4gTIIjSgKnH/
pRaZXzMpZhe/aonbfY2wLUSckpCuqkfydQYisHNTJmJ3fRpxPQqixnaNdbBwUTn0X8hfFfQeh+/0
hvAxjQJfqS1/XAJwF6ge0Iwjy8A8cqZhulB0nBcRNvSfCrOVU8vh2otimMWHh3k2g5hNmp15stj+
YS0DEDUeS6Yf0jXwxvO7BrIgcLBuxxXBVhA1f3BOc6k/dGe1DXt0sL3QFDV4zSBYDXoCSuHGazx2
DZoCSzPDH2/YtJNNUDOaK+ZR7iLRxDvA4dWP22TGBJy8wgQ9dfPmCXyRzgen4KmqEQiwg0CDWGFR
PnaNFBYDnanW5kjOU2tw0Lzn9CUTk+WNTad1NiBooBbWubFerjXiIMM816+rylUXUR7ANXcULu2+
a0luiIdNJJmJgC3U2S8eZpF9x6blCJP0iMoasglNG6wGNsgJ+R5z5MgJpFi02TiDiNbHBMuy13fV
LLHklxD8/QwLnU98PNj4J6kLRoozMGmoQoiXQN+HNuWgOPOM1npqzHwfddVyJi8WLeRaqtDKBLyn
kt6CQOU43FSPppZAMM2ozaPWW9GyEVrirtI+a8qiiKfosnB0lJC8IWQ6ApjLG+QqHJ5d2M3iWZxz
jMu9rlK/u4NENZUkmZkfpqb2Ytl/O0t+fhZDa0j9GWMJb3Bemzo4QreC3lCTsUPT7quh65O9ABHP
G3KNHX2zagQjXdjJOQxO5+wl+1KDbwx+6ARsX7DSEhC6q55VaBbSysd5CvKWBPEia0lXiFhCL7El
mLav9FosXBm4XRUEVwJjv/XytX/cM4UcyTmv9NlqAx1qRdBCmwpYk0JoIjokRGMonSsUDGft20g3
k1W5FX8IwtU2QuJr59N8MHo7ysuMZTfVSaiwBNufhlMMXVvEYKjnu/26TXIVdkk3092aAzdiVDQN
RMX4VwpJfWp4sWcERWRLXTPgbHIR/C9Rzy25VeuqypHML09Vc5r0YW4XgbS9oyC89BYlnylYMe7B
z6e0GAJQ9Qja8ttgYbB4Ic3z43BtQU54ucm+Bx+gnsjBqAi/zZAkGaCrNc0BMouCn5ArCi7pdw4S
beCV8p3bhMvePSWTNoh5hZm4rApZjulhlLKsKBQFbEBkn4nLfuHXKGWC5OG8GxS1hr8C36Z+xZbW
sgAuPNrNFk8VE4Q+vEyMALGGg02XIu0/W2aYIKHylEjGCfSgJzRKZqTTsYwsqHrFgPTYuN/eLC5C
cXeLJt3AOyGHi0mu+Vx9zyrjmxgo25pwJivoqalrrS0WadZIzqHdjODRJxUcSgF/+4c1x5t00tuS
qTmnJ4WmlmhAkFcRtANkx3PlQUPNVXJfvEFDM3BviboPn6OnU1h02IK/i3/Pe2vNV6NGF/G4rB8j
LNe3DAkqyht1hrFInX3BWbpWcdj+iSNcJgCYrhEdQqTgRQYF262JWyhKGVeyR+BfbKEt44woLA88
+/K0PFQirKfJRjmmnVLv7Q2znwBVyA2MuKXifwaeT33HhbwtglHELDPuszsxBG8rgwu3IXp+dkgb
xEMtUQFms1NRtYPdIKFn+llHbyRhBRLpaokIvD6V20AiGBtUJqzTGZOH/A+0++XCaCwaAxogaf17
E0ZiuPV7t3+eclo5uuIRLfK8jvTbQEH+9kYHpZWEpvgu+ljlXcHG88i/z1mi89nxFCDZHlas95bM
aElXKFdmTRQFIdJ33pPrZWvUidF81IwU/DFChJrTetcv5VZmmKyWxmmPG4jDtYo3kqEoqegNOPd3
5tpjKueFOat+erwWuHZv0eLmYY/Bs4tYqoBFkAFGtFMz3NIE6q98W2ZsVe/Vzz+Mryx3eFZvZkao
c+YxjD7sybld27N9hSE2iFtSPSiJn4mEBW04Gj2C3rZ2NjxuM1LOzn25yXkM5x1BDzKrEtXAgu0p
BzbSPFpk3m2dIp81KLj1fvdyByzQwUhD2mKkveEL72nIa0wooYfK1r1kMEXRNM9toEghnTQhjmyd
6xO+F+egBwpnngMkDQV6IYfBzUVhrzFy4V2JEllEuNcuY832OeztTEzFXfE2ZtBIVDMxncxOmPnf
23Kt+qmc5dGuptjv6WQzBv84frbViGnvIrP9DI9uJcgHQ4FTiDjn6NiA9yDuFfzY93PYyYoXRGfa
GbteCRJKpip5gEBXsU08zw+MOw3fQR85Qj7lqqcBoCROaGxZ79Rmrva40KVHaGpkKp2K77wlC73q
18N6JXpS3NKyb/ey+TC0bJYR8okRsXIaRhlTyfLTwinZicKvlIW5F0GKsXMECdH0gWpQl0z7THNy
8sWeKdsHm32elT6Z3Tm4o0NxxKW0zQR/9MLCYs6F8KZBFgbjnpmQQIAvot6uVh4c4cSogeLgyAIB
l10e02F66eV4BciNVxhSAT6MDcqeMBZIOqQZF2hFvfkZ9mjmDuHfDysQ+mydumzPQDfD6S+H19Do
8aKYO8oOuqkcIRgjSxwZqL0x9abwzvbSQnZKoUA2PxbNnzasyguPwWNFmL4PlZB/pyVX570LYtJO
0SbTSBIGggnu3MeO2UqpoepmveKqEnx+3XZOtn21a2OtctCYqRHEmjzA2M4IKjdxQpsXJzIfpCg+
XaphUeM6KdXhJa/dP82Dr/1bqKj9Fv17A+VU1Mg75BAr+6bzYgdN+FtBo7G1mwaedZcrHb/zPRkS
bNNBdKciJUT/fUBQNlvCJfvhNyxWLl5x/0XnHRx0bksQKTtcPFeHxQ/S8Z1uYFfUCzJKemwtlk2f
8LEEJ6jvAH6CwSPw2xOS++a9Wh1T9cqGY6jDqDmxod/vABCueh1c10qOO/8lJdgV7Pym7LttbxUG
wzpuVpfuOs9kCS7W0bdzeeUK/CvCFnYwamfWix087fOG3NFXGA/BJ/IRE2i4C641eklIC+i8VgJH
Mdd7LOWyqyfdlVwIp4+8OxeuqyOuRp2hPbOQxscRGKGbaApLLwIIrQdNMk33h6Bch+KqNstEBXgK
DcHKMdpF3Eaflx0/T0IiKzghT3db+uO4XpREzeipNHwpPryTqrZUrjxIW1Adze2mgibAatfmDpgH
dHtgEQef3wwfkUAPtCpQ/zC5VuWvZvGccIquKkZNmXwM8xMucDuG6sTPnV2twtJ4n1CFBfNAbrFq
t1XxMuG+jDxehtwxQHDK6bFlmoJ5zpiQw+HX0S/l34wiA7eadYh33jU4V7j8Qoo3vL3RzPtdoWDJ
rz3TFSxBYG140ZBwMtSxiJ4zykfAn8gFBGJCxqpCM9nIBmONf9nil4KQ7gCfghTxDZCoY8ViOyqB
LfG1GJclippuV8nI7ZMsT7km17S3COEnj98B5Sd0PpoqMCCaayWM4rlAPdJbTsS4DO7GLub8I9tw
iur9xE0w0NdXtxQaGdfYf2WVKuPAULdByfb87rKH/OQh+iL8tvvF4/m6tu2h0GcBgPiWIDJ4fd1m
72y6dNS6jy6eqUxw3MeZUHGTdt8RjIdBp1bCKSf7n7RHo9/nD8x4W56YFp8MkdvkYyOPdqbxG+J5
qodkGddhtPzILE4JGpmceaNvWI3hduCRZanpGBocVPJiv7ZnOJ57ibV7U2E0ecappjJCOuwgBEXl
2robT8ZPz+G+u7R1BW/w+4gjTGRNmopcW9USl4Ud8BbLmXOn3kqbVeRyGCDYZfKCqH60s3FK9x5I
7Y+F7J0m5Ut4I/Pdq0aMHXc6EzrUvH7lwmUHbz2Mx3beFO9lATh0Xgsm7WiyEN9O3IWSwzW5iWMC
gGrLI1ManCt+6bCSp9oedVa9fvV/qh2OnnegjPeRfHd406JUzK6MWEt9y3tt6io1bO23pyG3VojV
VkvPuexhHrZINxBIRsXCzLVIE3A6oUnmwjOhssub0Vx5sjme9Sg3C5Pk4QpVJ3Yo/7M7JpXWATZI
E9dALSPjv6OBA9aXcIMnPsz7boI0JVHRB9jfmVh9ODdDI84u+DWNzvkyCFQueenFuZ62m8N5xGmt
45FPYmgwzIteQOwM4MHQx1T03jJvhKrTRd7/r1JzhF6kQnVdHM+H/2j14gzygbpQFnlcVB1uwSNb
AQX5DUClZv7OOc9j5H61FffF3oDa5rApXqpTWkGg87YXu7YHhaWM4ohZV8vM9R2K0GsxkYbd0wZS
K/eA32cxsp/dff2dGZBfAN03r94k7009zOZJFR/2CW09FI8M9R7BSOjXxvirZRBAEJtXDB9ZFyDV
6u3vFfQetYSRvxn7nARJ3bk7HnsC4dIFNqkQDfBghHCtLtO4FFShqRKyxLND1lMor/8Bi1HWYR85
fsaehjSuNh2yxDCj9YHM4BLoxhV6yReItEhlPOn+0QC8WXfAhVAmk5AzI7VmA/AZKj5LrLpMY5Db
f4V/YN0qptiZGfULZXfIzm+yOfPCTWm3PeGFi0iC1tBiikR6zDU8qDi5qkg4/wcf2uW7+usDDfYW
cy1EGIqDXgEEGkvd4m2LpRmNAj/cElBx3o8eH64aMJUh3Bwkjrf4nmkyd2B36wAQf50hizNk8GCa
TmocmfJkxGFxnNC7WLVyIKXV5MKRt0E7O96bHEN88ahnlz68xbg8D2tcLIMrLj4R7P1PSWaBOnL0
EywrpGVttjphG+Vu4O1rUPrnRy7BNYwvr3jSOjCNzVse7xMMX4QkmO47HJPt8ftD6b6oWtEntrH4
NBQ8gwjPVIAwsJKsiQTbA4IgaMgFUPYo9lvLTdiRCnRazDU8AUo/sZvWfPnL2+hMQThbfbw99fqc
2vntCusQYwgGn6j1uYFq12ucazlVNoQ3rZVjv6zPUR6dYx5jAJnOTbSMcL8Pvu41LuBxp3zGjEJr
5WuKVcHt+V4Vvv3sXLxGelGY3w+8uHmbyIA5eyqHibCBJH4VK3JubF/JgIiWdB8zNAJPDyC5ghhU
nKOCF9trNy8X5j6Het2F4jvueGmJ569t2p3CL07v5wnQTUs6ARxVWVDCgHW1EWXMs+FCUJ7rhdFR
b7q2cIn96pdZXG32KQ4iAP1HTOlWaDHl5G2qNRWCy/a6m2g6Zpz8W4E2LcDOaTseIxcdSmaR81F2
Rp4tyCwBXsHVrm+KVjW7fXBV04I87h0ZPepOq+UjoF7VOvKqCUsZUlsUAxqa5CVTBWY9LRDOr3De
3/knLr4sZa+oXDbVFH+S9jKXxdeaSylHGbpFY//dcLUsEn8V0kHu3uN5u4DIEz9G/csDXlqWNRtV
mKfNSIUPVzs8rtIaws961H6SVrfkJKB/74fGX3ZsJdU4CucJzT5QZZM0WLZKv0lhypWc8BemJGKK
eroBdobqWzb7pXRR9ulLGdKpLm2NB+/P8OWsbQWs5S3hRHqbdcPA/5RRa8liwxs/N4Pm4s4Bgty1
l/1Du5o8gww5T6krmXek+iy5aZJn/Ff64QIPOtnjy/wo7F+gIyUx0k8gcH8tLb6zaMGbmYeMNCmE
NtpVAQ2VHIWTbAeDaQghgJmoh5ur4H9bKmhxVSQISGZMMJSD1CSMwEvRKSOkFg4Ob31ip3odaWTV
z60bAQ/verAAiAqckkWDOYTybrxwc+cvHnN5Yg08gS8lEMJZTSrvNClW2Clu9DA6sG3SbrRQhU9R
Ri+PH0pmY+SKEev7fqZRFS4HzM8gcEXo7jY90sh6Xgq14JA52T5n20sMstlkfSO3EYZjRblMz5ic
aGQ+zspwzpcXTnw7Fqy/fGJgyvE2uFkAzF3ubaUD5zngfzhloj6y9u1esf3skNy94w2A2wD/h2vw
5fDXkntutXytEMqRzfRDq+ikr6SowuHJaW2TAyDoFZWa0A50gXIRX3zySmgaAQ/5YBw1AT6MXqYL
aeS3gCZEh9vmt4W+CqBOMO5Hft4SNKUx947vTZuEzz820U0vvq1r3+hCqq4mGuHSfTuMo5rHfCta
54lWG6RYRN/PwxnG5ET0wL9f/4a48w3Ysd6SfBbClu2r+Id3ENxJWZ4xOU5UWG0dG73S0i4aQ4Ia
nvFZYnQ9a+Q5TAEqL5CmGJYlbh0FbwBzQeavV8lLaLa/JliVEyUQ3BmNp+OqAKzwkx7NgqX8CN9d
wHPqzZNyNhpJK5DnZwDPIG6WhrJnDFj0/DjhOsJapiSROdXJK+sC/BKzQk7NdP49bHizOfJ98z5f
nCn0dHswbGUhZ4xCr1toFwwcfv67M34AEkwpGkwtZ/weyxqXPFmJ6MX8uqrn+cG/BMZXG+kyBFqq
Hwgz87TB1DKZFtWOCZswLBCy7tzWueefZAWt8ryTn5kwm21zh5ld76hudKtUqDPDHC2gXhhcDHHG
c5QWM+CzPVdaEYeQSDJanDD63Soo+vtzthdUkTwxxbCy2jG+HQyCHpFmDFGpd2m0B5q4ICjofSyN
OSUrQ2T5VpvaDDlHfEtEua3eXDCy/JnDX/fgqofge7jhoU06CK5/piCTVjAqE6BKdN6rc4tgQxHn
+L4C7zfQjo1ts9nuBXiv9HwY+9NIf9JhKhsE07uoKgVKt6IuVEgQVfbCFpMftsgkH/EKVfHKY1MC
EtuQ5UpNxW+oIa297ItmhvQ6szXUy55s9ODBH6v6oeOiYbu6v/5MzsvMqZYs3mfMrXY8FWnUdk2Y
dvniGejLjTMYkNsPKN8bYL2NMpa+PO7zmbyT6lah/Z/iXRug2Xe/HR48jy/cb3mKWnHaAglNeJrs
TNhNLA5DLHoDprvvVmPELoz/F6DQvslXgn3O/I3zg+9tkU4deSgjZITl0ZAYvEZCz8XHum3HVpWZ
oRuCfubk4mzRyLLAMKSKT549pmOwqLJ+bruQP59ekOOWRDHXYPygS5VBtHcVyMMuobVmsD7UejWf
h1tnfl3zKXdDV2EXh8bW7+Wv0+3VdgsxnwZQBEg9sOl6OP6Q0PoVqzlZsQTHhf+HrmWmFm7knNSZ
yuAriT4n1uXxNBrQwPqrW9jvUeIroRFbfvtkRGcx+r7Cp+hNbbhFhNUvejc29yI9OexXsy+bk6xj
z2HaIW/Lu2aVtTmBU5/neSYHGhtrW1pLlOPr59PXHZTgQ88zkPO8jgDBjYlnbgKpW0cwgYziSsNN
ZvpxFbrZFnot/gs6GtYJenmCs4y1kWML/0ZA+VoOUiW1auOK3qpnDZ0+FGJ5ZRlR9jeU9ap1E4n1
F3L1Uo6qlC20cGuJmKeSBi8zHZYBct5xHQ7BSO0TW+8aiADtXEmJb/E+t8DaymCU4m0lPKR2sEPR
nfFiN9/vCyjLZQX5XNDLVyWH8c5iFnzDKntI5DOqtcP+3Y1WF1irZOAa0A5IWrG+SIvOHUCa8jSt
BbKvqd+HY+nQ9lhKwHysHL6masEKC+YYmAiJA3aet+Dcmf6tT8Xp46yHIpm7hUDlc1uvSMFqHioO
QVSnT70BWoSZStX+4ixBF5TC42tN2rZWFTx32eFnPpfeNvsSLBPiSwTMTspmsw26B0JvTkwICJxh
VAyEh8McJmxw9a3V3q9Im/qsddBaKAHqf5k5nS9BqykVn0nWk+jSkZrQMftFbBkWa14+t8xALt+T
PkhgkjiUQ3BPZGNoju2hSGn4+CLDwPSdvFK1LdUyau3Hp+SWPvwbN9gzL+r4JtyGIPc6o7aP90qA
bt8t4uBIpCJHZbS7cITRXgVb9KhBgxZYGrEG7fvSUzLJWiLqf1oRQo5v5zDfTwSco/eFgyn2eJ14
ygqzab0Bq8NZWgKYMFobUk3QxdEkfsAypHYHHMglR62LSoUj6ALdcrVN3XBIUEQyRf+Q/eIYujpM
ndaiyGa89Kucr89qUVGyGei2w5oLo6o51E09nLS+Lznp2twGOz0Atud86kHiol+03YoyemKV4qvb
IQeKoJhwE6LTgyMWHTehtAmO2Jw/T0vxFLsZCqQLxOyhdl/pz6J5dXr+bL/tcudde7Ha6ANZ3cyc
A6Lzgd4leZk3/H4FYUlUxMZJE/wyMGiVrd1mnYElbTEG153OIBD056KQmO3kArJaDCPcMWLdgY/O
07NscoZiQmbxU2vC60pjDecxQT04ac9jAOcTD7DFziD/p5Sv/FEcKKBqmmNcC+dq45MffrO/A+Xi
bgeMrylicrf6qLoREwc2dDbOh83EPFI8L29CRHgJPp1iMnoz1LCGc1maFSas82K8iS50+xKPHQC/
DpzKPBh/c5FJneiLeuijawxGNX2AMQ2rOpQIiQusJwQZj/5/qY1GFSWwiDa0duYwdDywheJAZ/x9
qdeFXdXqjkiIaEXLSNtenusoB4+5ngU2gChGLCdPd20XjQGv5ONPyrIYy/o9+MqDCmVDCx0X8T6h
Xz0qiJNnw2q/COIquwwf4Qq347s7v9Dii59AYcx7lHaMtBak8Wk6FTQK4trrpRoovDCPe9W9qSy4
tMEAdEk4xIQRhboyovTOOywf8R6jbJmO/ACgZ5rATNOjkgjLsTQlVzLCSsO25sTio8dbqlp6QZsE
NvwPwZnVwjlNujL+ZEyjG2lMSsfJZZa9TtJzLRj8GiiVxmJDQ1Vsa/qKTRoghce0TFgSXIlt1Ib0
DvQ0yvuEwjheq0WopK7CAQHoScqgO14I4XzD0LhLodKP34dPrDI2wtoqVi37/h550zq73dVPkF+F
61HuyyQB27ctYdM/QjcnHRtambB+sWSfF285oTax9LA5I1ukm6MyXwnctI5KJSqCUb+0q0Xeh8VU
xVvhRdYfUkVt/tjaAJ2kH5c9swoAnyHCufddhFJEht4YN9PYMumPOTqYNYX1nTRA8JOvhA0YY8lQ
Ye1/r8yvhIx0Y03SGwWef8LfJPelQcFjzGAeOIb+5eNe9vlj+mkhcf6ZAafm3TQxqK9p2AKyAhey
M3bJ4ahXNR9BvC+jxNfxfJZPcf25cET3JuRRwwbLjqQ8DrnHdl6ES9vdBDrVt3CICFjDfNpcPqBv
qsBTE04udZfZnad8LFRMJkGDSzXzRN7vAuIGPkA1xOdCVE6W0DCYcVwLy4ughMatpwfvZOEL1hle
GMrq0UqDymH5ibyj4eLzME4HrJvw/oQNrDzRSbI7/6LdsA10kyVTMGrLZBJAcMeE4ejtDDDa2mPG
baDeQk8ao7tJ3w4HXaWMw7Q8isuoyn0wNPDCmG8j93sE9zitdAKBHWenrfSIQOurXY0xFrT8sWu/
lLZdyPN1+fm4W6+3r6Uddt4TWEUL8Lhq7cfCrAbRPyUUFhdKaEDwB6z6/TdEtTpsZSRSgsYFjMyu
ukVgN4mWNI+2KVUJ7ayeCIJydSJQsUrv9ImtY2dew3rk/GmUImC8lSYNhNQ+Hzh9Wh+8rwtunnHr
Mg1c9jxVCQ2YUllBIRjLJVQkoyZdIzURY8MnJN63iHrLnKc4KKQoBBJsANLZs4rdhgl3M678ky/O
LqFEjLwqLtaZsuTGB0RfZd7Ba++AwxLtz+Hh6XL/xRM3lEKluupByBCQd43zILxdeN4l0LMy1PDC
mC4J25XKi+Uja5KgTcgCGjxoVRyz7a/HObA7/3xdQJr4vBBAMmGzno3lQM8Uozo1RW1+nU2IF1WX
1iJ0Ck3zHkUamFNZltnruXL3ocfuk+niJgZnt6buAOW/I93xgenRBOTJZOx/fJIvneKbNvidHR53
W+qYOiGHRc9qTwNMJ70HWvOV6YabJhC17FvYP3mkUYWpOndVlPdIIGgvGRIYOCsvEheNVhPxjHJS
hlYBFUkU1c5o3UCb0LA2BLrthRRVkqYpkJjnW+crafY4h+6tJPEnd7I++rUng9rAej2BGKMIaG8w
x177PpQNCu+QzeU15dTH1ND4U9K0GpcatDN+1y6tOTk0wJROMhGIok5AHXOAwXW/Tb08hJx8kUZa
cqwDQag82xU+dSkdM9jx9+pXjowZI7yMZHv+UxEKuQZJJGuTrjWtof6JPp6J8IX9VKnZpJ2FZEcf
22S+Qln2j5cRGn2FUYtrL5z/1CI+iuwQVF24wg0T4eP7VtV1k49lS/QuAq5IfOVoppgzx29Xx9vf
+shnfFfxg/3Q6AcFB8Ba3ArNf3sCLqT0P67YcGHO+CvowWn72R5JzaCPtN4tgPmqRakkTIBWMZK9
5deszsXB8IsXOrnoWZVgMRaMfXFxR1SyJmJjvJ4fuVaa2uVBRW/ccjKxl9MAcVqWmFWLwjKgCCZs
Z3FWvUfgU2DR1Fb3kLNZymmTRGTcVF1cmf9cc1DkIX4utI42RyzI6HZEILv4sy3r3P8KqlYCALX+
IwcqAXSlNvJlqtGA0iPeK9ecui3H+7Dx3LSmYsDUs34s4RR0Wk7Vk19nCJj5vzLzdu/aLTbhC1oH
qGF9op7eLAWb+SjA415iSVKCSQrJ1S/TpTu2OEQzeTQ4UgXUC4C17LTeVY1KBfJcYAvXEHafGhpR
CSp47DqPYDPvjDxk3Y6aLDhvKxJgvZaVzpAMbeR6zkqm7yfmsp4Hb3X6//Kac81z1e4DyJtF/W+s
zPC5RGbEF1Ph/B0UweII5EAXYSznt0R2HP6VyU+WKkIo0ehfsvyyG/LcBLSG6FGxqB3xKt8xGEoh
95foYP8VdshyvOnoifviWI66QvXuMA+TlVtGW5eGZ/n2Vhs3rAvzxMMn/siIre7NPcbuEFC2jRam
G3HtkIiSLIfUxASgJvdf/EZVoBS2TLCV/URIclqs3IkR4XqLP3DAvs9kspFWxDfhYHtLXDFRgJkS
V2pTf6xo6f5jC9bCxIZAXwkLvJsdBTWycAU+dK0fS+m+b0fpcJkipHllG6m5+BDiMHF3cFVy4ILF
Tnr+RZyKO9PXAccPSYl17wafwWyLUGR+c531jAEfD4EeMcZtUOYwjhIQSXS3zvHgfBQQx11iwkkB
w6MotE4g7SSYLoKDBKSaiA/GvVmA89dT/Sir+xQ1JrE+zziT/WQVbDnQvfSCkYZOTHTlm6TEqa79
BFF4hwFexhinIsg7RopGEd3d+ewUjJ4O5apdcdNq5zhU4Bb3CJiU0nmOcDkSBYKOEX27YCxWJlv+
PJlm6yQpP+vq1cLYVxYp2Xu+EC/l948l9C2mGUd+sE6kiC+3PhvHtLKOFJdMllO1mOOxyfRLjx6q
5HLtUWlL9dcZ23UXK/+M4xR7x8WP+GAy8GEIzkcUyRozsBUjalMRZM49vqVwQcdkhOaSraRfewlD
4za9n9Y1oDrWphtmX4t0MsdHqPDpFfRuoojUVq5OWlZev5FWyTvdtlOorMSSwdHQfH4c6qD2HInT
T8SGMyH+hPrRKNyHvLe+dUbX+Px+O2veCnXwT2TriFlHvHznnbtMvEppOsy9K5X/t4K8wXC2q7vl
IIfWaLcgE+nVSBlY4Y+6OCE+NOaW53beNdPyB6xGO7kEhLj84drjlORjRFpmqV7p8EwtjD8ylfQE
BS6neBsWxSTVleuZ4+SaHrg7tf1d7CECIgEQ2TUFyZmAYXXHvLG7QsC9+krSSqW5s5/puMjcQdGH
36E0QHpxhy3Y6bEVtESOuiqCR9Kw5r9ksXO3/XfdkfAP3TA7TgF7yevQLA8uBVNbCBhr/MsLgg2K
BHDoq0K/nOua97ghvMb4WOvUPuTJ1xfmm1/syT2jMIvxerocW/FFCw2FrZpzqbzo0kJOSUY14WyH
z1IRuVgwICIaaI+Vqpe/UHRi/xLcDmgXuiTwM9ylipk3ZkRlYYG34nZa3ssTuchZpJBP0JiTneo7
/k3ezxIDQ1Tz8JeSnNqWNA5v5q6Twwo7YZzCVZ+0HZ+f7oUSc2rPyX3TgZQyZgm5bPVLop8o7Hep
ARQ3eGlyDudvhIkQhHYSfRPlvXa/H0V0gFUppo/tx4FCKbwcXoT/rjLA8cCXgBUYn72FtZPZKHNF
K8pxUcgMDX+o2W18/8uLw4MimBpFVOIEUTiUbuNJjNxjm8J8DBzT7R0F+SKj7Haybq2iHj/WtREf
txwqhYLSWarceV0K2trCvRepVcyXtbSWgWAIzCTcqqalo/6k9+5mWyWJ+Rq1zubFqxVS8HStOhXa
8TDCdoQuTUD3uZotzdLBlYkqlsSY2F3RvGgmLFQ3vDjDoks4Inu2U+1YJ7DP/mNSYFfTmntW6ksg
7OwYxSoXJUS9RI1Br9WCKVN6X7QFK62DwJ4TYmm8DZjPmD87r25O6gknvNR8FmrdkXRBYadnfA/p
/zX3DkR2B5D+/jYJOh25lKHIJQhPzzYFF2z1IS2qzO45y0RS769OQt+COo2PXBBN3NiMyqFQXhAc
7Ds5nIbju5t6VNZv9SsYfOQeqZvvYoN1aO8BSpvIoaQjP+/acKAstJaE8gT/PABCuMvANLhHHrAP
wZ0BNvSvRh/kKIWAvzsFm49hH8tk8/jJVPvcd0tPcDOIjyq3kogfehAl/vsuervHpbi64dihnEb8
XkHv9fOj76EAcsHwYYawjFLnKJOJrEWxZB4I1s2oyMM/JifJYgBtdWoIQDC4LSX4XMjy611GqKsN
HDQloovsF9G0k31YwhOmM7zAwg5dO6T5Y5zvrsAD+Ii8v9/qENoS6GHxOrDodH1VE7OvuROpjQ1f
Im2KMWzR9iwSv5R6MkuMLA5XUsOSoloLzQaxEBXYuegYxdXJb5d28a2ODe6VcOZDu8/89oSwev96
kO1yhQsH1nnsDmh3gOP3+rTmojwErQTvGIXfnFB4u0f4y0beHDAsHSMNnVdY9zipt0fLsHQ6PE+A
RudRe/IzZylBif2/XTGEVs3zEd8oOntQF7f8EiHaLvvr+LV05QQwlU/peW0TJdWXyHZ2X4ID2Jko
s1V99OhH9KlNWes+EebSTpSZbC3QvcKxeXF1Og96gbkvOHomOqI41u1rhUFwFf7QWoY6zcVWHyrd
tC/xN56iQc69f1b3PLgJvUjs6BHUuptDFDNU8pWQOST7dlVByHEvTRVwY1PAld7itwGbkRwpqFuy
yQE3R4wv6B93nerpxtY3SegWDPzGNbD95nhvPxxUEB76NA26QKvkA7USeyo/KZO9k7YEqiGQ5q96
T0jFBoCDlfTSaKYpa6bpJNycanJQGbRa6dwy/+Bk1Ep1zsqXQusV9fajdd+V1lahsFjuA2FiLbek
Ps7fSyvDyiyK9taHwB8HyZxBHvjp5HgWi1FZNsVzAHiB6LUtaHhlu8xCf4LrrW6DX7M9zaDKumtt
HnxMNHyqTqU3vAjnFPXbkHU6yMKJdabSeXFIQ50BgKUN5sfJqE8/7BwrEKGbC8Hz+hohKoi5Oy3M
O/Cv1kp3Lqi2nO/lHn1xQvpOfKjK110bVTssD+uS1LPs5UTDCmIQkagmNRuIR9Pg/mmkqYXZnntb
HUtTjnlSLt4bPHA/r1SY2oVBAkNBabI4ODRavuBZ2VBYSShb/SEgp76ensvijzRyTz9pa7sa27/4
VxQcHz1ovGKNH1UAzhixpVDQngaAy+e1zt58s25aROx10mf0uRGgCgSSYAGn3m7llDKYqS0MPLGT
Icl/1v2I3Pe7O0WEl7wUJecxSs0SnxtXvk2XUHruW3+BybkSFO1moQIyEHczrTBMSk/encvGhG3h
in3DBc5Eth5kJp5iacCxgdQlsfl5h61Yv4JrYZVnj+m9VZL3W+bsTPTEycJV04MdircNxXZmHcBI
hp4tIXCP5hIizKgAaIfBP2FV+XiPrIK1Qy0HT5uwF/M/9ofv7Ft2OcWvOlybTJPDhelyzojCfvFb
+pZjqdRLByCfAOUcxDQICj0BDI3/ksPfnoV1uMSHqpFi2W5tChFiN1MIBFyAuyoFVKoBT38sW0WP
VWx512CZfvOjssCznTeecamInNelm+oIVqqTynWzCslhC1JFM870F3MyJKlA+H1hoOOMLpkc6WTs
w7pmIJLu6qraCEPJlLDAufI1KH+OZwLls/KvF48WUxU2Za3IfG8mM3449n4feblWqBgGDDMbxz/M
/hcdNEUqAsLy+KvejGvGUMNfh3CstMgeSf3NSEx3WkTMO+JToZGJOvqMwpW2t93v5MV67Q10YQat
d6rxvSmItzSE9ck8NXmLLbVoMM46EzIYGtZTBy6Fc3WOTikIvzEHzf7q/Mgb04Fh0mE1nwX7s4a2
ZlKqofa0rCTNOIGJ3x6+Ay+psDLeOGJPY7oRvz5Y4lYi0OvXOEVwuAEXVY8bAjm2b+LF1hpx9R8L
72YFM1XRWnrvvyhT5xGc2s4rnWWwNoTsJFNe8Hhc7A23dC188+RWcfCW/oWAaoIAniLjQg06wCwL
8C08eJESRDbEEkY+S6ilh/u6FhkxZlvO8x37QK3sNCmy0kfnRtbF0fmgqM1nvEuDfRCkfom07L6w
3ho3djrrOxIskjDGRwCesFac4pPicIrwlHVgAmDdV6urFNj7o+xipb/RywF3RanLH+FZpj50vY9w
ghC+lEBjlaY7XRWW56XS0zaBG8ZEmXjEo6TAMy60bdCQ7eisvrDn/lmJZ6DNKaUCDhwG2OZwF2J8
Jz6mR/mHnDbJs+a2Sj/SBwIGiI/ser8R3im5GnmLKj41mBeULjE5hoRcIR+bglWOHhjImUovCBkn
FuhUOcfaf9X+CVYTOrmuZKI88E5gT539kXy2gjtkDR/iuvxW1sV7ArQDONlhQOdMNi1wvDun8Rou
X2b2uig9FZ1Fr7y7Qhu4K4K6BdQbsZIgpFGxHDNsf9E9V7KmMVrL+n2mKfFMdR1tWeO8Y3OYfTax
60wN38RLY4Nm4wrzYEaTPz1kfgaklG+FXMYuorrcCpjywPAmNAb7qUg289pcPzQn3BSKnbPTjnas
lpowTyMjWXp1TGEVUC817gewx7eKPpCeACAap0DkLYXCCEHG95fyRIm9wXP4Ll6VCOsvCYuQq7/x
aeMBTepWYBUtwyg/GA7JN2Vc0I+kFU9D0Q5Y0xlwVUdXqrgE/Espn4frTOYvNnKo+OBvjkozlEdg
ylWRY0ainp6gUncmeoW2tnuRV+24JHhRVAOsguC1xq0YK2MFhxUTZR4KpTf7Z58pafeA/yK36nLI
xGI7oNV6Aui7BVSWZafv5HIhX3RFLN1S/etmPV++9dtFCOkejk8FMptEXWyi6y/nuifjFH1dzVxW
/eKIFE9WY2U8EP3QfkVP0jUqRgsD1g1CIPwm0oMJ/4RJXjqi8ciM+ndma5zvgCZ9hKdH4HzMiKZQ
zbttL0zw9Xvd5I2MdUvr1t2iUw+TCme75lWXUvTBodLtdPbqN4SClV6cNxaABAk/35lC2HJyCh8k
WjXX1zYvOpPoFqmTVUJumwk4LcGrB5OZOmPC9oNl9kk4ob7I9bCYgItuPH1rsUYN645Wvz4fIhvA
BAYiqZrf40t1ZcW8YEV0nQ576t+02YC8MVuVg+Tghp3L9WtKbMMSdwcOTaHw9Gep2QAtbQG+9vV8
GT2ZK/VfeInmMljMx42y5GFQnzNQR7G0WY3XCPgOpKyvkKuhEXA4YAbVDdtdqSvE3aQjEDwekBYj
9ep2z7Nvv0FjHVBSL5+nNrMKzAbLhhUMoeiS1c5B16RmQLQYDXSOFKU65lMpnYGZ7l+zchCwAePt
wlHfr+LLiRucZdT1Qfceer4RFsCpPapO31z+ATQm+mP6q15Mk94xe1FEGKvwUMFxBrEGa1RrMGWc
fWNEdfH4ttBrqB+2VZkaJ3o5eUU6lYmw2iRsivuoQIkEJ0YFozw1ThfolaDP029RucQf6nSh5EEg
735m6/oDbt9EOxMXQAqC3/d7zFiAF97K4GpnaWIAaTpiO/xmMGbqKyFCEHaFK/JPiykUesjpkUOS
j3B5zr2MjGbPvLnQUrth3cbF0ujssGnAY3WLgnzGJFM1yjkgdQPR1sYpSwrccskioxd1pEFO38zz
UAjl/PHfh80pyQ7ry1ChAA6uz1RH1UVJXL20mEWGCKBhcHk12L1QnVigPpAbXZHPKgrfrBkXgEYV
IqV8s00j2AsP41t6EiFYx4izxLSdrmoYqbo+cfRTdx1VV8KF5Ff/eK4juE0Y9SkhU6kdpqdDP2jR
NfJa/R/bnuoJE3YBI3jkVOUfBb/5HN5G+pxihV2yKyw+ocHHrgLtcQw2IY8kUNuXeWrSjDDmBYo3
XmPxDu/QSKIhFRDWjcNQwbFIetgeZTEyASUxpS188uTfj7RG+PuSMi19N+9j3ZIvEvnHX0DwN4RR
WeaSckzME/+s2F/QwPTeksY/cmKJ+/2FRAgGREnnFOxYQIU3DSAwUaEaFH5mPPK9i0n/JusDqgng
wDeG6qHq57PWH4c6xR85hM7FY9yawYhBpRF0Wq8a1uoSfmxGqsa365hWaQz0itet00M9yTVkEEm/
u1ZmW6skk6/x9b53FXIyVSvkzAv8bnurkGBCOnuvxKMWJYQfDSsc2XMMv/WPAeSWG2Z6CMtsntZ5
T1D1US8siX/ygUSufcy1snIYPewJkQWeuzwjIwClu8GaBFouAq5bW4wWulur1wIdzpE7hIi/9h4e
Jl6Dhlhhhi8LBvaohTksWiRL68Qrz+6jMLSTXDAnZb+W+JMgrfkCxrpYv2KNoRJLfcq25hqXSiMD
rsxYyRR1PxfFFDkktAyuFGBFjZFMZ/mlsSBWZj+M6xL1t2VTfyQl8AJbZVxLiyAJhWPOtrlu4QzO
i21YX7GSNQjF3tUviP7/UA5ZCqmScv1qF3QGWS3buGIDpgMCSBCCtiD/o3GxRpfIwKFYpm+qaE8H
32zCcDFF/I2mDqgZqvwubZHXud6IGvBzmrPUGamuPfXMJ3+cCfxVMiQrvsFNxk4t1WlXppPGnMm0
b/AcRfxgZmt+C+jkdLkX0xjYJMJr47Ay3oU+C7CvW0GXem66vArHA2IJbt8DUibURAShFkfzId0l
xclMcRJjMbg57jtD+E2YM5itaoSw3Ao/ROHev3QMe3j0qrMCpsUQG2OzPzoT+ke7PKwrATaeKlmO
8DM1PzH0JvoqqirIs6s6DPDtXcLqyOBNHRTkIwtq6nLNH3r0LpAbaOaTmiMwxVGTdX2Xl/gV+uTk
huvlD+OhwELYvCUAvIPn5s11Dpzxb4k+sS8i/SkslxiuYxTVgL6hqSF07zh1y/a3mf3w3AHl/ZLx
vImOLQAejmdulyJkpKaWDBfjr9v/KvBpkNiWrunV4AU96yg42UksgAjzf+Ec3Wz7gUoKsFunsLkz
wBOfoZjiOJAb5VcbTbEMp0cdTmLHUGOaD86TMW2ycBdxJeaUGMiFxdEZTcr3+77TT7YoHW8KG5py
Xonku7q9ZlNokAFUdpD6q3oz4ssC+Qt8bBdEaOIqWqlcV8/HoFR2F4RSAIhpQQ2EZ8KuGcxfl03H
S6rFngSVMxGTYZDnMP/15W3QWO09tgnt61k+7K27vjBbFfqqx7NNtvDy6eLkAPu2Bvdak52Xm4sq
49id1NLXIle+A09/giG3hYlfl/1ZgS/zP07jX0j91Uc5+q+9V1x2cVh/a7E4/w2YFBPni0LtW4yB
ZoiniJAACbW0l73f9GsAadbzShLKzwZcI2/CXd19mcFuXEmBYRwx6ZQEwjMuNFuet6RmNXU7y2EM
iWU05szV5YPPs7HdgxmD8RT5vEhmNmO+DsKvECd9Liu08r6D2pNYHa/GFB18K6mypM8BN2NANfNl
YyATdYG7wrbSWbSMVfdsSf1WH2/JE7XG2kEYAy+QX18ZGbHYrsdmybMDKc4MVtLnS2/waBGIIUI6
4BMuMDT5h/w1c9Zaj4V+tP7VI7KojQDOwd9hHG7ZUQnc6h8DkwDJ3hgxkp6+/SCidCUqNBy/0y1Y
arOwGnGoGkwMcPF9zYJS50XllPTmMhYece8UPlvpdHA3o9rDoCKKjr0JNPwugp+qNSV+eT3PLngz
LlyMz4nT+2i/hp0mSFK4ts50iBUbhqZ8pmsBUPFVU0OKq4SekiwvnNl6Nb3sTU6b7lv6iIg9vtM2
NPUw2toe2g1iC4TiWk8Q5QdKiI3uVBqaiXWOOusUtKH4sVA0XTf9jpJWi6WCl5myVGvyy5U1lX0s
1yw87ZKyv/QR2DCZTy4eKxnqRUPa52KfklKVbi5Y/FWL1du6QXIb7cG0AAxZsiaS8QIUwMutTrKq
UYej6pWQZ5DMXPiuMrv5efBXmZ88cG2Zp/hE0zpcuKqUpvFqtRN6tRpUAaBs5R59o4kYBXJR1JMx
Z1L1JqjyczCi+RJwVteKsMfriY3Bh9uza9vR57lGHK5kKJMDhyFUyx36e17jPIfwekyuE5EkZkdD
KZjokiPk8z96NSha5GdKGhOeNBJuaRs2GgHSLh7SPP8AfIpv856rca/8RZ/039Vu+wn2/mp6h41U
tARrDGXU1sQn+Z2kvXDtH21GPqoNEhf2XPha5wG746bxEG15y3sZphFxr8NZb1wb9nArVOg3LtL9
1ddjbOlxpwnc/e/FSMoY3wqIduE6ZUPKwSJ6Yp+mQqsoixro4SwcLU0pin3GXHo5RoCbA19wAFL/
4DEZBi5qAASUEZSsDzhGDkepsKMV9+c2TzE4s7mSEMIpvXF3R3R6BxIVjUqKg6VDjL4jS8s3y3Fp
X2MR8rdaYKI3W7kuW7zlbDJBO+Okv6UMk6+dPVkAF7yBrZBzQ74gOTj/nd7BD9tYiuL+MK24sqnA
moZTIrHxf3vRZyvd7INA5lkF+hN3RWLaN7WAu+UZkqFoulLuimwJnSuLqsK78BwUdaLIxXBHicPz
7U4ErmYcOxLpe1cffZQbeG+ZG5rDatD83rVfKBEpfwjXDyT1I1AyG1mPCuJZ7VTpEhGzfGGr7Mqn
T0/qqVqy7O97dPgK7xJvX2JqZCoAfRUrs20nXtNpA67+ZtJoP4pWZQQPEkHUngMSGTl9F1xB3qD8
Y+zFYKmKQ5hl39x+ti0Pywt5kYkh5E68c41WUmaqEUEkqkqmvN8kwtYuMVgvNGaMrHwBsWmZDaUE
OBTwEUUOjCoYE4AcTQFV+GZ+gxaURo24Ey3iOuklFsz9bKpH1QfbdQmIB8f0/KhaYW1o/W3S8WUZ
4VoQFi1Yqr17hZN7w1KQYX5QhB5w9ZRoVui7HmNZIn3oBAZ3AtO8N+boOpmJL2DOAoYiHDI3BJt5
4dmAVNi5kj5VsibzX/DkKBzEu9Yiz6EVnePSVMg+MH+fc5xfIg4K99JKTcFtJRBbIw4C6CTFSdQt
+QOLak3mdNQk6LGSeU9RlGIH8XZ5rAyv4nERculSAvu+5Qx2AMzMwXwGVEXo5rSi6lslms1BD+by
gk+Zv6pWxIntsH7XJPp1F5KspPGHOagfdQy11Ckc6VMgQHhUWeQ0mcc3JQUfcsTtHuru3dzYBc//
qCGXrdPWE3cj2Fs5iJeSYRBYUsUx5vYOf5t/uJNLaMjxmbx75x66CFTNjpk6JxIbvgGjekCfZ2qB
YsgrK+rtJRRX6i5A0JDmK3ZWKgNPDU8PR5gMdcNelEwjOCKzVSgmKh0bbgJoceBlJNeIxSdZjwh/
Del2Es80MkaT5IBQKaAWPTD81wP96kEffIykZR4WNJcrOEY5Hy/cLjE373ww+HVUC3xAO87clHOl
bEVogEhoR7qIVertsIB564O1kIC3llabXeGUxHZoDCkuF6HNXTRZtCYKgvXMkBv2r9UScyxDDrq2
0CoGyFblpicRh7IbRzq6VxwEP8ycNauGqvI7Vm3pLLNcgYS4i1aKRvjkCghKkP1axZnuYFF79JK8
PRQ1Hl+WobHkSDgbMpNQT8b3Xw0hnj2pajt4P+T9ViC6Pwj/rH1KqIB3G955+/HFMBcl5A4H7fkB
tfEK0AT8PiLS/VTXY3yTcCSE6LgtB3C9n5rYdTjKpKq8x+AS1e9AW2sMFc5tyfoRUXGBPDgj1fAv
ajfHFD1E5ha95nKB89GHbqcgZJXjVVClUfHa2tOgKGZGLSTrFnHt5IhxOBOwk9gNN5lcKkQIv/TK
DZE0V9ibkjDCdhT6EFDXGVMsGp7RZ0YWUF8l7vPWc4gViXO98yOABkDfGNgNbo2qV4l/BR5YigyY
eK07ENi3Ozw/hSVCjDtg2dk1wFYbgfzMz0MZHKGbRLrK1w6HsR5K3uadsVc1pYpHzviPjcLNPWP2
qsLGGnoKUpzjei2upzQgfD8U3RB8rz4ucX615s1hRZ2VFf3nh+mWqkx5VYSMfPhIkEn15FULZKQH
rd1RHnYnzqWT74SuaP5iGuNI2IKR2fO9RgG04JlEjQ9s5c98T0p45mgipuHpJmiVpZmZ4uxs0C5S
7EfxRrk6FCP1kH/5QwSvjmzsEnGWARDbA52gjJJHy37woYtpmnTlbNomyItFPqJx2iLaLjQaUbfD
9pOAYRhMH6WxI3BFq4xsRNtWPOHERK6t68NS5xg4eXd/MZJuXSEG6akJXiAQ7u3fH6Swykvo79NU
pqLyKdur9zrRKelwriEp6/u93C8VxWnG9qSeZdxigPaphBn36DWpgGg8bZ0S1qOAufLtf0JK3kUd
S4x3rg47HMbhilkTO6f6p/rsiHsO5j0/GJ6eOtxXI6ctwwZwNepLwQyFfqKCB6vdQ6sVbN7pxb9T
TXYTCQ6nccMydNtGSeteo+ufrPC/EkkhqtHUM004gDmS946pQnZ6MPF8XprxcvV2u6EMkuCc9py/
TpvZ+/Prwu9ErY+y+eqlE+9N6pHyielswyPZ2JDIyCvLWmb0ZH3CkXRs+yHdpcIfdcrQ9rK5L9iC
7RwCjSKEUk7HaPq1hyYc9wSDBePb47yF3SXf5a6NiPMl3RQl9mBRf9CzOWewSobmaabMIyseGcYG
NPUCAuOY7I5LNqyU1PD1ssuFVWnbeqTg+N82CKpUYEnqkmIXNTrAKUl1ci5kQ5Q3pY2RFWq7i8ZD
lCN743ESfi7gC8heVybb7UAJjrXpWKMUo3WToVc4WDBn0N+3U9j56UZfi6mhxCdN6m2uJF+g6FZR
BuN/O5mKBSVB4fC/Pp9BVaQJ4JFVsOvUJDKZN6K/HWfvdQFOFjNQvRuyhBx2U7hVfdT5xFThZkiY
Daq3bRT9H23gqYWRlgiyrtuFuFUpy8Rpw0aUBQ/hxLZbRi5QDquEU3RYH3JiWMiznOtUODxSNbWO
z9sQsWkCB2Gt5pe5hMeDV3oqCNlLIcG5/AWzzP9zfDzlh/bHHcwyQy96Damz2PTuwUGstW8Fw/d0
b5/RRniMZSrufgdfi2cS9ZLqZCMkPCGryGgYtO8f3JT9FV5/KFfUFUclLvKSI2UKLBZKimQeZUkU
RUxYtMEd4TnKnCuxTKv/UwC8uHzK+E1PnXh2eC0bycHe1YXS0U2y/KgKx6hvBoFvcfNmS0o7+EZH
KRB/iSLxAaW8WSmAghHDBVxdWA42MnHJ3TQGmQyI0BsvCedafv2QRHc0je8+kLDTRutzsh37LuC/
RYd3ckM1Yxjjh+uJA44g0W0283U6826JsuioTDUzpqZqNqlqVSnxNdBryRZ3Xv6QoqfqtVNnAkRj
DlTPhoVIO7iG8pIdUHHQAlMP1+LZ/SrRtfBP6ikAJ9WDesQdDTtaesjB7VRZ7lKup6P5hk/MJSKm
VES1WE0lOwBB3P4f4Viuv4mceAhajWblOrvXBTccClbJPZIRODHfLP1uGKI0sQuJ8TIyiiYuPMAW
ItKXeNiJ5HDvDVmrT5Om79FO/Ap5lxENJtSZV2XxYW3d/eywndpesEyopBAi7X2z0BMSgkm4aoxX
d9N/DRXJF/H+/iGKSCfuOlQWMcSb2WRU4Pw357Yj1iwi9+R+htJuCYnvcWE822sOkFZKNkySLvzP
JhEnJ6MgFUwSUh88qTo0p+UGbsFVNaoKowz+7SnX6UfRdwPhyFXhHR++VRiDFzkqDme6SmB7u52X
g4NzMCvXVcdh46P6tOVSAqmoOVjK0896MOPhKOYqkKev1QA07lAr/F2yBH24GG6kde7vE4hWRXOn
NSYp13LW4qTmRqtHsHZyB81I6ePRnSOiNBxPzzpkGN94j4+0K8WkU3iWmzyCLF7I0DGy4sh6PPED
zNxeM9uMsEkAvDN/5VXKffU9Ucx2QqVnHhtIzvLdxSc0fDb7F+g47KQAvjcO0Ve5ozz6iHlpVGg4
G9JzCrWAf+oG0u72gom6d/3SH5OwuFOYbGQl42gnRGuJ/IsLc5OMFJCQH4TEd7zHnbj8OZMARBG2
w4kxNSk8mwJ0FLU1J6DHtHdp/KcaQtmAJemAm5YIyNPv3VonU4cuIjYGBbxJE92Fub5g4XlFsW4g
0pikTrDDd/9huQ0wGUsy7vXmB6sFihhHeCLnNDx/RM/MBciVqxxc3Nl5+eJ/Ncar5y2WIBNZlTPV
wRd5lroYyPq93yiflKwX2mvhxB6c6gbmWH2gTBCX1iOwo4oiAt49vnc9+LDy2xwdldy2aEMxRcse
dLCMa47oqMFiBpYjf0D1Uz0tXj/wi/Tw1WpyoIQOXg9Wis7bqmWjC5ugGsWDyUB5nqxrrE3aOutH
dFOgXB2B1uIV6snIIvSzahZo7dAv8bSBO33rF2j5KRWln1tqA7almKN6GG7LZF4KKOfzPM6V/DoG
zWNUQCaMtUotIZ0FHysROg66SxfVBYb5r4VIkiAQRJ/gINnbG6Wfwj1DD7sy6tzZP2xZJ37YKb0Y
gwaw3Spwiz70MalWEc1BoEpky2B0z4CtT/aWIx5DOEvalXYFwQGTSMm+mWaE8VX5jRjefll6w+k1
dEHeGu09Z/THbfAl9K2EFuX6IpvHHpQDQqmtL6xCiif+D8gCoc+TCLTYZk/UjLv+wSranRkvZ+lC
iUDBHU0tKMeH1MXZ7nPFYQHwiDGPyxZAXbfdifr4tMIkJZPGzswZcCuSSvPkyBOdZrbqFlMvaIlZ
KNpvPt4LPX/J3vhgDFyA3ie5v4+f0jl6L6J3QBWEfRU2llOcbMUdHi7+FxIBClVqbvDEf8hOJjbf
8tRD9LzHLZN3GFFP8iIKA7gLemu+vit3WmLv2lH00SwoLGAYdQgEIFsCnUEIz8t8lTF16vf3DIr8
AxtxEDSQZSHtF65yS6lPH9UfWQwgtvcmTvX6JYOCSdUemtUdD8CP0QLnQ86W5yxIjbzE6Qza6Fz6
9V/FOhsuOZuX17pMo+kkFdbtdvm7Cf5xKfp2Y2oC7naCQKFMeu/LUNnZMr9gSXfHms500ZOIdcbJ
fPYcQvfjmHBlITXt/akdXIxQeHObPO6VDWB0vMvkfUfZumBn12Q4Cfcb9NT3YG7k3E+QbQA5lB6d
f4ZwxVVXT7M0yzCHmIq/hvpBkkCpsdRBggAzPIONUw6EoBUl/0z8TePZ4gCd2zLQMSTAe0Jn8SuK
CDcDKHBaOiZzi5EjOdyNJ+AOYna+oC6kGKtpAcs/ZahPuGhZ7ITj3GNowy4TaEiM09wRRbOJZFMr
MIt3y4tgBJBU2EhpniCziSNb3s9d8hDP/pD2dlMa8u9qMSHrTP5zBT+JIfv7cxE94bDSsYXazQA2
0HncgGZNYNEsruJ5Ced/b8cX/yZJXphmvevX6UmUc5Un2sKCfsjmWtB6DPPTbuBXsZsG2OrbQgso
bS/yoLbCjCEvTCLv9KvmDrVwjXcpdEza4q0s52tXD+knRyXatSKXkEfIT87RDtzcMuJ8s5al9xx0
5eFJ2HrrC5jtSgzxeoupWP7XQBE5tT/QoZIw9QXz1BE+BptR9wUgT9w6jz1TXuxi9WD3iaGp9wfP
qs3A5MgQ7ItDxlwkQxqQ+00CO0qgKro54/tyGS55KYj1hqxkpSEJPR0ULiCK7Y5tjEeIDrEu7S4d
SjqjsRCaxNaJ7U/CXGZL3zuLL+WtutbQMZOHho+y35NICnzyrt+CdgKec1mWVlsDY+d9CGOM7TnS
mAhy1oyvUbOw7cZF0wmm4NI5/UFXVarcIOe/grVH6QidpLP0ZTdcZVlDdyuGuIwRc67SZf8RU5Zu
ELVsV4izrp3Tz3kQ0GEYrmu7qqM6ElAJS6Zad1Wv0U4B44X99lIfzIgItmFvKtifa/GwoqCRpLeO
HGgvNqvOPc5ZLxp7OS6fWgxmhajIFb1Q9gRsYgm8SkLWOeBvvIqe1fdqpa9Ra+qgT4+nGbrm1Tee
Te6GXhSxGY8gn/ljxeNYrF5+fX1AmBDS+u7/9C+m2MAU0Wq4hcu7T/I3b9UKMrmfGJBhvQrVzXX5
J0/joYR858BbSKXt6+2VqWf3wRyj1Hx4oFAZOaWgpX6uVnJR9jXGMqInCJzNxhmZvxDkqSUGZc93
AeN8Buy815licWH1Ko0oh7PpGxhD3Qiqlt8rsbxxLF87yCCpVAs0Ja6pzWTG5vt5U6VlTEa6Z+dw
raEI4q6qcibM1DlxvyPgUZfwOID7Jif1dGYhTCS/HGOZ7jETsunXFcvhCaujvNTJxN4ub/TRI6Oe
xPydoAKdiaFbMzdm4Cv2pyxphffe7pH0VkwaQjVDxE/44bUzuzwwPh9+rCszPrlkhKG1/0NxoyuE
K8w1urgVgwSdbEzVPZUknQMamXNPVNvbQXOO1+LDyK6z5fkumjGYsnnBn4XXpukU2FmZdb3NpfuY
FrlYoSlEJ5o33QgGGSv0uvUTA3YCNLHaWQsfUrOe5/f5xNEJNnjTjWbCAtf74XSgjbF8M02+0eym
56iY7aFQQxMw6ahLsygfjuUg9q9RAPe4DXE22vFxMeJuaTMBb2Q/rg+cPZeg1JVhEcNHHi1GFSqU
f/iW4fDiXCsDIdWyV5jr+XPvWI8sm7yZmpBrxzRyRSnwt86TGMA743L9SQf0itn/QCEBS+I+Wc0a
JLDKVZt/pxzgPtLthzIEmLojP9wK/MvjEq8G8d6i6ZOID/ZhGegbGPQe90w1UypUj3uqW9FxNGPC
h0mnoY9u3oRznPIb3Ww+lP6itH8a5FmDIqfaur5JO6C/8YEDq09HJ9JLzyA4h/C+svuNLbu42ANg
4U5jqk6PSz4tsa1kZ0aAI5d4a/N+pNwxRB0/mi9gDPMpa8uk4JaoJ0Ali11LUS6Zk8r0R8/5PWrt
FGsemOq1lAxu8cmErZTo/zQiCsenNchwMXBDpmINtgvqIklj4DfCJYPOMm7EZHUZAsBuTyQ3V1u8
vsfiZg0rsAdCzAZ2AcTJl5kHRK0p8k4fRxQ4tCekSamEmJFw7x+XVUlE5c9cfKA2Bx1F+me672/M
24kAZaheY/m3AWmJuGYbxYAdj3zC3osmQIdhERK3Jqe3yWVPKG3Vf10xwSXkicozdPM+Ntwpbw9O
ApLGMePolLp4RazwSfFEFrTA1sTXFprNYiuWJ3aQJuctR5dHqrr37nx03wLe58YyVp0iUbf0EjYM
axKj+PeGqRkMRb66JncbNdBjNuNzYene1YBFblIwpfoD/3A+ySw4kYxsSGrWCLm6HsM6hPBuIHwY
uzPMlBeaILdMHCcoOITJ7BVTjBQni13NhacRK1ppbrP1ZPfzBq8MXw7g7t9NFz0LIUiyJs7ATaeD
RviMiupYw3auOmdN3TRIsnezGc4rMx8k0dyMSfJ44jStwnyU1V31jbndaAcOnMGuBPgMiUMHgNNT
nmCU7qEah/C0sBPkWhPXBT1zmvQTJoaLQcFFugpM28Vy8BK0VM0VR4PJhUtKL9C6dGAyIppEgDnz
1UmhYJaYVijZynv+Iq1V5TdxpBirnNO/xGun7Sxq1UsyIYXNjkFft4qcd1KqbbKxXG5nd8i9v0na
QKz+90NGmCJ6pLrXWfWWR5k/dF46oF4hkeD50gPj7XPOX+tVmIjDZxOwAV1+yMwcyLOgqfhRs1WU
dMwD3Qocnof8oHsBa/uXbMZIfbuZzx1Ov5VjU5NLKeLZKAWK/G/4Lg9AXjxebSjwdUvGjMtuTpjL
wSdvLoSlofG0IXN4F8HGpVAvR7vXXqszw0Veuw8SvxKP2Ltft+IXOnWD2+834bK6IevjTqYt4Je4
y4yDRdXquNpC1G2hRl4ARYCllMZF6v/kWT0OMkr7DbXb71zbGaiduV8ztNv6iiBGOLGfLm4aIInm
t7tBvAiOWEy6eYdspLQtD+XYT66dGn44YLwDCddaCU87q1xY6JNx4PF86J1DxZlRG0qQEoetj7l7
JjG1EHxSasxvC3hmNaOnvs4odS0kleJLjnAz9/O7whDmjKxkVICqa3K4/uQRG3ulst3TAFFadJj3
pRzBZqVjy4uRJ3l4hXUvDQxppQxdalzTfpwvEMZ13FkAPRxT7pDkrqOJRh+OK27ndMQWeY0yzyvk
UpzbTlFOQBtXDC+YJUJh5peg5tNeZcNOzqFTORru9eLiWQw+F1miwlOakcZA2sgAAKT0Wt/oyf/2
YGGnNwH80B8V0slbBkw1jPtJ4PDoflEtTOVVE6sJTdoOpOePHdjuqwvCkvK4YX9nCmJSuWjpgqrm
lD/oEAvpZ/xPD1aW9ekHRhLlQkUJ6g9hpEwzQ7r/HQbJBv2JuJmt1HT6bO5VPEz7yZcxJ27hoRpN
+iov76cx5z+h7vBc5SCKA57jwgDnRvzDeoczST1NeZTmeNt+OSmfC3fwfR2OJ8Rxd3s7Dy8WB3qA
rRpMiDhaIMomUT/TciBoSzQmFWsBHfISUkIHGvV3vpbZhX56xgsX9M/PoEpfl00oZrOQ9XXO01rp
JFrBueQcETjm69xOq9n5BWM4E2Yt+NPQ1kOQgHYQovtMbLI/KL2nsxqPtdPxUhIjgFTcblDwmpBT
OmtLXTXn9NBE7ugeUItOz9RbmSrXkzsbU5s96G6+VpPrzuoJpFBCYKFBvJIX4crC56FrqgAdz/EF
2gMVgvbhU5Zrbv5V6Ks56fqufGIpRPzh7NLlQhB6EW+TZSbloigZgFbuWCFB2tk5LysColzX838j
LQmkHzIWrf3FOjXWOBAJ+i1NNTma4Y88kfvaYpllzyi0XL4KijVWtjgcesIsMBcvDxEISAIpK1hO
SskRhs9bspAmpIsm/076NtJrL9BYPNo5FgqGhuReselfGR+i9sch9iGMjI01qgNVFHxEuPP2mHqL
NdqxwupzWWH2Atdt6PsRYA1nxLjCx0Mq6BaxxULmmfH2D0PiGsB1F19AUDqR/tImiOhgCtkdAgo7
oahd7UE9dz4DFdc2D/YK7HloitwzlJ5zTd2HlIm4w8o757IHY38FtHTUdzcpf4+SVzhxU2I8CHSv
kxvLBO6DoXw33KQjli/4rF5vYsPkbXKFrWMg9S/2Ygplg8WPAluHpQ4CMkCDzjxRzo1DWcD6mUDn
D/a6sgNWfULUGcBNOZj4cn96hOu4Gjdin1DNBk1gzQqSlNapOdRWzAGyQel+vuauB1LymSSGCzvF
jD1yAJ0YeNCWCSHatPbakk2eAHQbGn3+KQlKmhWvkycY7W86o+68chAnLxZvxYUbkRuZSHdaHeNI
EwtpRhTmrH1ebKv+xksl7fiFKonkplBqGuM22pAi5CcnUpcbmh8JkU8DU4gihcR918xjB+wxBs7k
gOJredg6k9LlcZPNr5IMrbynlWbzpHRDX0brclsOC9XVA4HfB9s676p7zsytRLfxxZeyMCdAEoO8
TtH5yStFoa1IS2N375RLa+SUEDp9lUMpIYUrOKsfyXtcpu9KwFPozdoznGnCxpxsn+TFAyBYZ0w6
5glmalhl7zaP0LuJ0rONgc7uB60Tl3FLlSTbRprJQ6hf6etbOTSwVxK6rZmOZw1Rq6eXhS4GDtUx
VfR4U90u5cYyNhyQehS+kKQI1aWM7JE7Lg735eNfkkuoF2BbP+u+Nyw6cg1rWXCNdjHvt9fXtO3q
lp7KqhUYrVr2sbdUdVn5LRlpzLvra7qBTG2iV/LmtmOG6vUKSY+v0y3cw3RAHNfjfA7hpTLY+qIu
xNwGamOS2FYTF091ZxPpiwLi3uhmcZzIQljcudkWbgUBUH80ErF2gctCEuBVJBkQKIactLvc3Daj
pnCqJNEf+f2zgDz9I4ogGVbJzijXf+hEoh12HEcWNDwNPsLxYRVrvWqVM3psZJqviSP3sKAVn+u4
v+BXRDbIBG9Q7u4vudYzIo8/qaKkqSdxjDZLTHfFGD2dAif9mPEG2fIiy9iMb2wY6NpdMQiNSUST
6DuPgjJ3VUEwrCGZuCCRXzKKsh83BBcurxpk9jESOxYx6hqb2qerxj/rk5sxdLXGE+Trtl49TJuG
EfeUvXLE4RIRJyq2xJIQXjJYLbltbCYBtZC7FAiBDV8UTUEjPAQiIBM8d401DriqCsq42wSmZBeP
f+sM5Nyak6dPIFnVq0Q1D5DcCjRqldzQwNiSMWi9bcfLYKo/4iuGSCLCdk2rUiMXSerTHMZz5ju6
5PpM4Vks4xR6UCWmtVC1l4Tmsq29F/YSVz/a+PR90aw13GJHajkL7SrZqDy/6Zj+QWQQS9CLQP2i
DC7IvZ1G9eS9kFRy4UeQ7Yxj/qwFvwzO6wEvGjE+qFV3qQMUoREGvx1GtCNQKHg6fK0D0Qis6ITg
rENcqDL4Hbx8y9n7TMILjVgUGqs49FJDp+dZnflZKkcC5NZYjVl8Ut1j5iiNiD56HlX3qJcdcnML
WsVj6M4K+sCcggYOP9uHW78yvQAMnsFA3/BkBEEtIk1vB5z9Qq9Bkz8mwkj9/P8RvZq62izZppvr
IRJ0GjnGRl9igddgsVxCeVfouGF1C9ADeJ0821DxXy2/qGsOofjea0HrdsmiETFlArgjXAT+K88d
tE+U/Q9mzh8WHzJf2/AWsx1ZwXZrPAzNKd5vRK3/3QniNKZ14D1BWAWc54agtP7+DH9YZFr/bspd
mOLH8ARkqNFhQ252kTOJ/XiAMKTOChaC/O/yOKV7sz5XBScKEkbRqQFTkirqmbyuJYl3bBYm0VMo
//aPnJgK8UlX7s29619YXjBL16kBlSzHcGoo83v7zYkQ7ZTubCBhjyxiODIK91qGN0H6k9XnjbC+
0x5RHC/L1teV0viYXVLTGLdGbhRkGFT8mga438rdNUq54M/mUa1HJ93vRMIprAElfsB/tuENH5RO
fk4S+uuKYwVPKnwpn6YaAdRVSXLt64XebxVd+TabXf6Jy28aM3NEtqDcwXaHLOy/WErLDkUO+lCe
WYSl3VNtIglMq55XI4V3wDjKk4pAkdVwQmifBK8KQy006Vvktj4ped2coM2vfDdmPGmXw+o2aYj3
UvirL+zX4yb1QpXhIBEz3tyCjeUNgCDjvbTbtHefrj7N7BwLzg4eTsES095SmEWAYYPv2ByI5xqP
P2vDetwmfDi6CF+kAmmIBa9hd/HD+XuxTWBpTDkdBhukzD/GpOl8t0jZFDnD5Vf8/XYoYI2Nuej7
rnQjpp2WdtZUirgt63440GvGe8bokXMrAdKtx9NXPrP5W7l+2N2bLwYigP2VOKTosRRcLYpJlc1u
JGAmT4TKalYrfAX6CCojXWgxzDhpLn8P4GJBQ/M8l3gfRF0xInDtqtknOBGH9d0HYLJPuBltqIKq
rrZ1Z4YEfmhSGzLgmfARb0axv/IPe0l5/6OBXutwbZlmYrTgnbXo4nI20jhXmuPkkIMH8qfNg66i
9lxJ5K0iM36Lv1ZO+MMh1GRAVY74SKx7daNvPpz7ryETPQw7cmht66ApahBLK1S83ikvTzzOE33d
cICpJPNgWLC2+Hhl5k8SqmtJvFoxtppujEHgerSwgkha0tO6kJPXJaDIUl05r1vBE6bVRqSFl76r
9E73TB7Aj4s4/CyKHM/7TbHOb/EptuzzJuojmVbcnCGhHfiIULaSPj7DWvF+CKPsgi3oCp0hxkAo
Y8RdzbwsNkUyOCJXZrextBAkWhaEh0GuRX+nWzAwMym5Zr5jK4gWUPCMX1JPYHRciWd+Qr4P1TBd
8lGEogp6lXlLfEmZY/OhGPPqvmIQVUwQitvqbTRJwwnVDbnDMZlB9H6DiKEt7axmrd0haiJLAoDN
fbCmFXaLPImjQtDEhU6The6Zp5OdyBw7uqiCwYyLp2auZt46C7tMluk53Ypgr5sqFEI04IAlqqQ6
OVXDmKx2cqSHpd/HUPgczz6iqaNArT3y+blrQhzoFdOG2sT0i9dUrHUmiwTBX2X7Lf4omFAudS3K
S3XQF3n3+JBlMF69vOtxicTu2MtdfRWayxf++xpP/rO9o88NdXgm2Gkd8M0WY7JSJlEiAA783VG/
uwHkdImTaFW6N1DPdtXPzB1bZ9qS/yUvFADJGcEYD+f7Z+3Nz2SGyFS1zF9TA4MctOY8d5MrLNjF
LPrmOpqRQu/i4hPV2S1EAGFHN8ThBPztD+d3ej4uhbGQVdmWfmtmhog5ExSymV+/frXm6ALnNQ6Y
sM5xeYhc/un3y2ASWndNb3UJGzbMfrYmZ2xJaW7NRdqga7AhAyjDD4OgBDeUqpyYFiPpQoiWyoOR
WjnoMQJ9yoXUsbJ48KtOW5tVgBXdY+fZW/XwDQ3erTHu8N+86HYPdtTS4f8UyuTzSSsitR3Dn9pE
EFRy+R6AJVrkAzA77DN52jfCbmoj4VIX97N6drhZ9DqKjFkx5kTmuNccFxWg2/QTR4SdOtkNudwe
twJVv9EFq3IODbCNCHb8Rn0RG6vLr4wd716IU4VARFwOWSF8aKQ1NC4ktvdtz3iHWYOFbuEpD7w7
KlpPgntZQoFSnYpN50Hvdrog3yYaqjNxAp9KWQq3ffGQkUvSeena4LQx8Jb2bPMtTwvOibqNPXbi
yu7NXXpJ4ywPaxEzm+gjOASQP8/qnu91uozo9/KmM7kSkij5JyxQuPcYjj3AVXr/lhcSsmKQSZMH
QLOiDbcDyHrsc+ELkiFeqRBNrEibjn/mruCJ7BGICNz7w4vJqgnnE41VDcZYfwHA3zU1E+oGDFLm
wV6yvag29jO5D9BjGVRAkZZQRqQBg5fU/2SU4KFn/mC9YZH8H3VMZSfnF8GVdLBudBWxOhp3Ca8/
UzheZf5KCsqDpPlcguSsPL/VNuXWMaaNiRfhs55k4fIhM1aoOUlKGurWIlS4XnWD7400pbmouZaR
lOxunat2hrpmUcAsstJYdaCmHq0ynpEVAYsUmAoweI12sIKPiBbCoNi4YdKShsVK4wum6eqXHH36
9lKhTlWTn0G8J8JGXB9PDEGRl0Njxd6kanTYvFR0b88W8FfEc6UJPSmdpffRx0RXaXjm1qXkTJ3e
sFSHG81c26vhAVYfv+uftpYs1RszPy2vRjo3tdDn3w6gDOeliCwE1W2QtOnHYHH70QRG3i2fR0+H
kTWaSDxdJEYXUmlw1yUmlemghUyHKeYqHyzUyukDZI+cM9MRW8ihXkSZKkucEnPfyyWcIeOUg7Wo
hA7Js7T/YcDk9Yy0jiETX5JA/3FcI40xiTpxTVQODr8VITTMqc5d97G5zZL1Mde0Vqzw5pf4G9w0
76pT+WRIoiDPYTwwHA/2XaQ/8vL7K+0AsHTjxsRg5T+Q+z0flsRmpC9kAjpm6x1U2eNWDBPB5Iay
SuJfNv/YsmDCudvee2G76PcObGg1Hcu/KzbXnLm+oWsT6uKnw4nq3BPqY2dhqfbu6ujMbFHNtEUi
UlDOhocWug/GuLCqiZ+SjBGS6nsD5+aNkm0gYrq+HooYkotWgYNUDvaXJJNZJUtfYixrs1PRa2n2
oq2Es3ra3TSmi70qcg8EQd8/eaEdAJoHiBp1CRP5xmQLwKMdk0LqGTU7jqvZLg1hF0BWjQfzM0Te
vh9Q3+E9s3bHRCNX8QE1QUGFDJdSjfWutPIEtZb/7l6wssorI7FfsI7oYP564sB+krkWbzfgiLaN
6CKImA9XLoyE7q7PRssNoFDJnubMxwsow3LoUhguxo5IxzrySYpkqeo+sbBTireoee6pond8GVXU
aPQDVZa+qQ/cP7jY//OTatqKbTrqox5Xs5/5ETvHbdIoglm2QHf+ksPXIgAk+Bx6MJwrRtB5hp3R
SRjB1izvOJgMfsAg9AXs9lz0+JMeui8T9y1t6/GvZ/C7+KGeNfa9y79m8aDqBxyvd3aZS3Vh63Ty
KhiGkauHlLNAsVN5kO4uag+swdEB5CqhAyYOVHlxMLOEwdib42CJiH2rRD+uZ3NHVzv8/UqMKBYC
JChQm/hwNkAhbraJ4N2xb9oFBc6LvGTHdWJ+/a06GzCBZe3HKr6DS0NKTFfxRpbkiJIIgIwj4bzE
qjTLzh8jp4kyZLUkVu2b5IF4nL3udx01XpdlejOahDGi2y3vJkxHe9DG6WfRr76J3vL/cLm85Iw1
EVXwOz/QFAKOPuUz8f0tRIDZiygvulsp5CQwuuq5NbwPYxowM0DSVY5KT8/bL0RamQkwmZ1SibWA
SHW5XCMcPAsETJQegSD9s0je31xqWccUorzLQmb+aKL7uMhLGov/+XUMEkyklJbF+RBUXroU1jQN
1//G4dkw4EOFVCtHLmRv9X9A6ILS5m8OKM7wRO5aib7XR7s8Ic4Ron4Sq03qnUXrR6SLu/zJQ0F0
VIGXb8qe79f+jY/clnAXD753I7zlF7mouo1KKw6S2q8oJm5Atp+44lY1iq+WMnP/y4KOHOIXAxeE
km0rooOkHIfI4XAWZA39KxJ9Zvo6H9rSkwW8e80zpeVqJAwA13Y5+9UkqrYuutnTpHJJwF67DwtE
Oww0Vw1p1NuxkgkJpZLeUQJgnHPVqjFTH28lWN8fQzMnjHLR0oxdLGe5P4qIsGpoVfpxJ7x1onVp
Sm3uvooPjpSCzdXtLhwYyLv710fzON+H1PCVPq6rdAbhdKR1uSrDByyMNyHj6aH1PmcljnX7jiQw
YRxOyR78brTuyVEhgc5ORCEdbWR5OZNaoJEWbngJriQ7K7fNjAaqW0Bwxjc7TB9cHaIcphAPS9dv
4gGKz7n2yzNZ3/JRCtW7bDOeS7K0djBLz/lF/y/ZcwbrGGVq704d41eSitOlrCZvqX6XdL3ytaxa
mVQ+zJNWrGRCiW43oB8MtWeY5t+9tihp6eHktHb4QCWARUtiN2xoAwCv2AYwUBN8WBzb51vnQEnd
rO/zTJE3pHONZsKzXFYsnTwY597kSzge0+K88DqcFAw7H5VWrQVvC1DwtGMyYazrchQZgJkU7fya
zWLMhWHgi/3ym6yeExlODMzrL4T8KP4BZI46Pb7FP8GuAINizrw8jcZ3UZb+55R2pPKfSvNXwv9+
WvLIjKh1YSkl6pTvKOZ+mCt+v4p72J0CWRfehlsYHngajvHtpmC3MhWuc0NvIVkMSuXcwtON6t0n
QhFx1wULoI1agSZN32lt/VeUDk743nBhpMarlnjXlhuR2yUdN6XdXAHVH0we2Ohk3qf+FMP7ThVk
sSSkyalvdkGTKHRRP+NG5weIGQgTU9bOhxCfNkkijIAaB05zT3/KrMcUpJcjdw1os6BOxjLDuYud
nWv2C+BxFxJx1ZTWIZAxpX6pJ2zmSh95LWXExnJsLG2H++InZTR9JpDjsTLA6Wvnc/YxNYAZId41
RP0SiCrDO40UpdLVLnqpPM8VBzcsOq6aY85Dx2xmjn+SRzZOjvr+dQJmfK3jSPTrJ9TdixK7W3uz
i/yZaBqjH+/qukVAVVnM7jQPFMY6uAi6YOZexMO2Vy7hp83sn3lqY0XxM3kfw+LZkvwp6eWzJ0tP
5VsDLqL1pcoybdJQPYRa04DlU0w+/fOBAU6IIMCwwdzXGuPQHjtn8WZjsOSaAb401OdPEzzYVXdr
BcXUs3tCC1v3pMLsbvrwWW/c/dP2u5AEC6Y+X6Jj2W5JlLpr2/9x9ZmOlznDn6bYl/d0TIaqqQ3w
0bISKkX2M5ZelDMlWjHoftOin1OUtFpKfFLeEBPSWmaLYFzYOIM8rpKqskorWulfR8Qj1hMd6edb
zHJhxbmDMCa2fkKf7xKjn0Rrab8U1eRwVxMCSVbgZJ7SQ/COjalWDPTpma58ZmjK02+niSn0Rvy6
RBzXIrIVGNDgxaiElTgpiciepgjDuo0q4w8elIwtLykf0CBFk7/4f3+STYXxlZIUHslG/HlSpYLv
04KDzkSAO9Q7BjxOKZdQXEx5IiEFedcSudJFYi8lanUIQoTvSh6g3N6mSLSI+3N7tqmr92rv3sLL
NAn/9HPRyCifqoPYqV+Vxgfb6ZhW/cBfLDWQGGOEuGMIDiEMNc0NVTkzBhbGZcT/f32lbBVwTsVl
3o3Q+xukWqDJmDJj0WfNstViWbFGXVuKH0eMxJWvdrSDuCuc6K5dgN+yv2jMiCzlYyRcN5EQNwCQ
VOayq86NErxirmNzsf6BxJNk+JDjZyTlqJM04n4PNiA3HLi2yoDKb6We9aT5NSU8ZxrZOfNm83sY
Wys6OjIxI10bNPxC7ET8XGvORM6ydSjxo7kdKZBOY2RBHP3KIYDqOQbcFpq8QKLuel+KyJ+LJ45g
syPZGf81C2umoCs744hBmlJS46znPPI6/03r/X67lguiW8boeDln51UA/U7qRcXjjUs3APsAATfk
KZeXHt6u7XLr3HM/pMVLxSUeRDIOvYTf7HJ+pCjSZaoJMcz5hK1enurIn+dfjEVUh/z4OReVl3PZ
3uJeM+/eEuc1MsjfkPs/SueTXNUyjXR2ijNs7BlaKQ5/M+Ekp5fIOzpHnXO7mue2BmhMh8kKvr3C
sgMA8iAq8rEQIk6So4gzq8Zp+hAYvDdRYocO5NCio+BqGOo6eLuFiAtu93S1b4ionDb0C++sK5gC
ft+9K1HKLo2kXJ1+l5K1yAjBZwytADd9hiWoYPqrNS2DgL/OBqQi5gL3tDEn9RyDzijWOnncdBjZ
nLNVAPbUQexOVB1KgFJA2KXMYK52aulwITIWO5yA2eePqAgP9t19vUB8KRbB2a3qk54v7TVnoDPy
FcGOlLImYpBRZ9cUto9opzfPnxKxr9o4OP1Y1G4gsXz3VLaY5QptjMPsxdhekXKFEvSKs2DVz5HM
qqJfJvYZsJnZzAF1nh5jrZHGn03opgbZ9FsqtHcGl73CkQgkJ/SvNAzn0Af+hEf+0mN6swz8c7Ac
KtV++InjsQwCjvNPRb1bzTdhqn3oyDBI6pKWArrjOhWRCxctRD2A0PBOMOp2z2jMkJIoVc5IKmup
6ocAQstgwyonjRg/41EErf/FgUQ81Ko0XdrTIkun+sd53ukc6vqOI1qSA140aF0Li9MfoVU2R1V0
ekKqNPw9ygV7RC83eqs6cSKEMNifcolt0Yh/SdnGnUXlmo+aziJCA4uo2NQBg+SD7bXpsKaf3huJ
aFVejV4VAOPnlsY27sz/LiDK15nlGzFdzgkR0ib3Zw3Xzw7pGZT2wAIvrs+5B3cU3LatiRpj5QF4
kSMV+dA5f7ywhKt1AnTIj0HsBIJjmf3Ug4HT6H3RtCFq2+db7uM43wlq19lmsndoDUe2oEcCJXrc
+WSxwso6yD06DobmZkz1V/hlixFeQSKPhbpljsLiEhfXeyG2Mz2WEGUaUV3NXvmNQokynaAetlyb
BqAGnUJnDyMiC9hXPIim7zxILEncc/18wuPfu3XBqLcvWjsDkMGCqkxuGShapU5TDVO9rhEfdckw
VXTSfurfn1/3ljAX9og95aff6m+TDb52MhLAedfuYOlzVtYT/m3D5Jb5IJcxW9eFIByAIW7SF85V
6lKbLHU/ex0ny8DQdNfRV49s9PRl5zQQoUTfsHphRYKYML+thktyVxDMkmf+tcdS6VQTlwIi9MU4
3WT38URuGOKeyy7CrFsW+lJHnN0131LlPdTSPTcdLpXm2htYeGgYW2sz2vTYPJN+bU7Y2fz490sW
HuOeAk4YlQ2j7gGrGq1NIaHKFh9RwC2ONp1SqPuyQdodq9avSmj7IZ89IvqYvoyIuHsGgAL5gvOj
FLLX7KUMhs8o1PN2SPzcd4nf8d1HpWcDgo4ZzMxZd5I5oBtbgge4hMYByMUirSlYxxN1KdzVtrAu
EtQSKYgEk5cCv9FhK6SQ1Hh9dx7+SV1bPg/sQX02Ni8ZjOh6y7qFpk0rer1mXz73zxDIBpVT8Jk+
hlSAkyAcvQkaW5Ts2VOE6HuaAn7eUs8VkWXJqhfLcpH2r4C2XDdkZdlGfAyRK0aLH/ql3Dlxy6xN
XU8uhex4ljaQw/mFpcQn9hAPP37wJ4boa5Nwu2izmZhyDwmxs8WJFshP8Psny/P4crnPQkXJtOA2
IAqb6L98g/Q0L222t4HMb2yMS7xJIluEji2nPSsxhCcMPOy9ulS2eistiDRELICLctJq2pfqoQWd
P2ZHWYv28lTJnDUx+XBVnHFTKEGb/313+RCqskFAj6qU6Zb+Z4bo6ZXZ//6aLhVx11OjEuVwlr3k
lPwzPRMMcIa1K2Swahx55WX/0Bs5wKhl+sZGkqq5/EYoq+eIDCHn25BddL/rzsarmc3CnTxh5uuq
c1hTd4llOs4D0GREBRPlJR+U/sj1H9Felc73n2+KU7W3Y955ddGxuNmrcyh6TtxH7Ej+4M/hKmhO
IQKlPt+qMMac68Cys40weFjRa1IRlwwFCpYPETE0jRbOVXMqsvQi0jtp/R5AedbS9osl8fTmD+zr
y3gH+O6ZDEkeJ1f+7EdrxgYLHmEm3c7IYbIIc7cC+E5lxNOXEkLLDTyXtnM8mUSgssXZovpRyPEM
3l1FStZ/fOtCK+iWrw/c/EqFYciFSpksmIc9KuHqkkq+mfMRe33oN5r9jhTpvNQ+74gxn3JWq5s6
CHPXVhTcG+9cVfJRAsyYyDyE5zQeFPB9DL8qyONqc1m6Xl1nAUw3vgw8OQzZ2Qr8zftmEOIMeCtr
hAILNJogc+HjnH3wcwIT5i8H7XQJZ5s0yYj7jCyYbNinYOJapHCKiBxHFoVLpRH+twUuBy2S5Of4
UuTJhkyHOw5TD20Uiwn0S2j4IZq3BA8jXjtIAK+sxFP+pX7OANsEWfeG96i+IdnuyA7jLZU/MW3z
FuntR6H4CePUk+5NxsXbao8RQmUyZQsUD9ZNbdjzlqD8qeJbNU2nP6Hh50H442OsD/o4NFNiJN7C
0pU9QxINxF9mMmrupyf7rcEDb7N0+RHixgqA1IhzbOiaSmiFKTw/FP3s99p5axQdnSsZIOsZtNWC
qH6SikIZXZKRYUP/GDGcY/vODQ4FQgtFo93U+j1yCCHY2RueXzyBULLQ4f4HOhyg6z2zXamACLvG
Sa/WU2D0Tmw5uYIhAEte5gyu9eussfPlaJDedjaGfdlkoYHV8zjr0lWPY2AcjN5uear9lfqjwoZk
egvpMMfnc8r3wK7Qvczv0Kj/nk9rcbzZlZHnQAhdYKAM88S/2asfu8nNJL2fdQDZ+r+AA64P8iA/
CeOMnfQm27k9SRRvjSbStpqwlnq0XG5f0EEM1zXupH3WUXKmuxW+CzzosjGAfdy4EySgoaJoyVle
glrDNw7W2aYlQUhOAzTtZYeQup1cPGTHnnAlTAylfjqk5Oy4Z9ozPNGnWsSJwpxkQaV9/3ecku4I
bRvLNc6C/447Pf0U0U16eFINKYEazm4+dN+9cWRWF49sJdtuSBQPUEjqdcQfCE6WctflPSc29bW6
uit+JUH3qOXeHuu0KL9KPKvtI+TCfiZcof7rKkkPJ8SDgQ92RB+QDDqNLFzo7/1i8rv2rJleyRV2
EAaLkwXsvspbr/Mw7sGULmR8VX8nv8PhBlmMs7E/k/3qAH3LehXi7APnBOwl11Ef4qaUb2okxk6z
UVi4+fRyMyF1G+gochb9yC++gXE1yoOaBEWvbMYmvszYiIN00WG8Jd6axHuHOaPt9poTKTMLIV3g
CdXGALbT64YAHbsJt07G9+TfK21ZPRSb/6VVYEJ/lT/7C3qLoXWZUe0x/qPg6lTXqJHBncCIKO5A
AQ6z854xZIx0HmXOOUp2k80Kx7pJF9wo0KmNRYrROaW//MZr7P8vm3RFul+n8J1HzMK1q+YCjXwR
DD0KQCKOslc0FSJHyxLzEVP8dGNgBwESdfuPaWHR/H+W9dQ3NmQWtoDBW22E5ENng0e1cvTztLJI
vCfzv2qUxIJcnkmP8441hObaJxFThnSk0icixa9BBAxmVZ2g0efTgguwEV6HVbnP6MhxuZc2IssE
MN8m4Tzj+O6oaGm01MInHBO//Ozghx0gUBzxGs9CfGEIGhWQVlnYI78J6WTNfwPG17XtyHi9pA83
3JBbHoTTZgVzrzZDOvtzy4FeihiAqeBT3y28zNHXwSfCuR7MWhj0i4YF5L/5emttYuXNAnh8qdNY
NVgYIo2Y3/AVEF3vMUGnC9Jh43oMgYjaZO40gLf+tporzvF6HYIUQ59BfNZ0Ij3VbTULeVKsZ6Vc
Pi7fWpUFxmncAC78mJlRONjdnd9S60eTlzaRwFEWipUFKrucZK6sdtXgWNNzGFNh8hxJWpGtZmc1
p8fmYmpE5Xt/5pCGepY4K2SY4CrZLUcUBa9o+DV65G80A+dKiqrYi7Ec3LNS0LqZcT2jDwSd1MTx
jMeyVS3sPNmTCpR3NXE1CEtiDRlJ/nDSffCxy5tbYEvXMkRhe7Lqgbjb44yRhysHpQm/f/OTeuqn
NFnGhfBrJrXXIznKT8mwwwunzfBbB+iCWRrggI9PUCThjg08ERErRWqHl3Oyo1jrtjY2Glc0lIRe
1NhFboM9PG/qspc3RwNJUhpnOjWQ9U6ZJDwPAMm4xHC7DLcTIccnGd70icVsUHeXc/7+BDkAb71r
Y0qrmxGKv3TX734gtffvgeYuoNOILx9QufT/KXRg17w0pTjLFARYTIOi1ObXzmDBWg1DBTI5r3yW
kLOgOxUinOZlRR70TRsMiJKEj0rFjhGEPk8dWMeqXPT1b/Vz1etK8h/ejEkpiG9lTONOqHJc0rhP
94qkhm47mapxQ11zuAKP5ESfl/pP5GgDChjfS8vRbCUEpSoCT14OUxaBvwn9sh712jIyEo8mAVGo
hn5rmnOFe123W5oPk7UkOgsgrcoD7Hv949+GFbBoDgUsk7SMHkZk2V1tQo3ZD9pgXS+K6Y6Drvl+
lwqrw3eXG7oNA/mu6xEs6HMdES/DwqfosWxtRu7zfFZAU8Qh4lHxxKTmHSdofL2NsNNJLmKDVKtN
E4f/uasBGhrNHMY4BOVYZVKi9MfFSE8pcrogs1wRsdmCYZ0+EhjWNLWg56rMIQrxhaYg9zghPBU2
8ALfH3vZ4p8pOivxaZ6zac3pb89tNjjTu3tGgFT9JH4gehEq7aDV04gBr27rXxL0GkSZ46pkgzPY
YANGwpACL1dfddzZ9m1vsF5DE1uNtKbZ8IdEFHP0h040yPlCY/dH3tOZG9Qon+SGl7dm/Cv68mg3
ua0qlP9cqO0z4zY9Q2DsRA2R4K7lK1I1pWPMk/Bn/nGzZ88Oh4cqsyMbzGEc6Z+VeP/23vBeoH9s
n9oNMTZfejFGF5X8xoTwMzZICk2Aji0RbVh4qu6y8slEnxzrQFYY948ArKJVexNC16ZkxDPDrlaA
YOs7xqhosFWf8Jj2KdXqLZzUYNuFJQrDQ3kARGQXykEFgNPsX9uG2X/acCpZ7GPwJcOcu/xTzoFY
6qa5IXr2VG4RxaJe33LHxTy/ZKBX8q6IAPG6EW8JlbE8Gz2twYl/8bKrFPUsL7891uIogIvLe8af
wgbdBRtFBjWe07D5/Wr6/EiN/BAn6E6C73hf1rkPZdkIk4f4V5Gjc5N3J5dVMpT7n9WTW2r7aHFc
vT/3sKhgEPJx6HanYr9YyMgK09slVrBlkhg/otW4Fp2TyKc7oB+IkjXZf/hC+4oqVfZ+ZrnZ1STD
oMQk/vGxYbnujczTFAgS9ch88CUTZnwKhl7tq0t9v9NQ3MO+O16rRA+tSTch5k/TZKu449UQgBFv
AZEXVdoAkH3e8XmHsCe7E1L7nlnpqgroYxLOzC+DQqL+gT2GNe2CstGRzbhS810Zx1O6bqmnG8V2
hC6Nuj+RnueGDtWKrzR6LN9aLxNZIXcVDU7Vnreh7hlHth9e62gl9k+TQImiKur3iWgg1Vm16DJE
b6+8QJKXPW7sW2Z5C6aD6eQtWL7lm5AXDKx9Rn1lEYeZRfZIOtay6Sesn49Rr2CCRmEUsBczmALW
KrlLFU9+un/baJvDjabrZ8CsHaT2pVvoNv75G3mpCGIb6LmCRaIJoqwyto+rUuSqvuZwx7s2E8CW
IXBJsZ8NR5R0JbfDNO/31W6hNd0Blhm0LpZsNgZg+FLZdlYYwSWKHJy4aFlDUqQvy/aybnMtLGyY
2tJhtYCrUHnoqKhcVCneIImluecrjTXqTMz8S4QwcRDfWSnCUocbM15gaTl/w5XgLoc+Bx/uGF7n
GqPHmp8eT4RY2CqD+zTyBBI0+8+66kqYWHKsaq1bIgmJfT1N2tO2AvdM1Fpf/1kLmQzgJqo0imWk
Uadm1p6l78LQCPKJ8DQGI5FYaja8xpaDKtQqHS9N5pCzs2h7IYyKYjZS5UF75wPOnDpvvmwNtS3t
eqJoiLJ9N/ROqJk2DFOru74tTJi3akNAPGnChQLEbcB256TEWk2IIxvq6DEPK0uWJ3gl/Wzdptn+
mCEC/Q3JqbcThdLE+//RcXMF/4Z2akjGaEtOxack1YPYenNGD8XvX7E5EzQyq4Gqi776xEUJxO7E
3F1U7DbM2HTYBD/ctBMVKaYHhOKgxmMZawX/xUOjijJM/3B5hgJEJ+/y8FedNl1Ua2POjPAsy4PD
lcrI8LWLhsHPb6ihQu/AonThjL9HY6XffxjRYz6bmhZEJs7G6dL9tS81cfcguBuwRBgFwlIsLZ0M
pUVcTqEngnYfJNqQTj7rfcyA/2mK+CeYEITbDB258elnulC0fz0Rtod/dfH3UeNo0AbEu2HZ1B3x
7M6TIBCmxPlolLmrZ9tFSlUTZ96p/m4OI9GK8Kwk3dxmKIxtF+aogpmgJnhuLBV0BOPu0bqUAJyl
XatrLdR87OBEATvZxuH/ojyZisFnP4CM+leErxIOcIyncg85DifqcEawVe+k4W+niqsUTIJaEKeg
z9c5fGJs5/yuszNAAGAm2Ia9VpUqgwL7XRIaE2gBvydt6p4zlzwhq5x0XZwUKTlXH/HRs7jpiSvo
6GlOIdP4QfjKHa3LOKAdzV+y5QqW81Ayt6rxCb8g7ZfNi3CnHhkOx8ibZenIIraSWX4yYC8qI7W+
xrJq6ALFiptSjCTs8vdNZlfUW988D56ASRLiCBp3wFaroXBs7kQp0ZAQ2wgouguWkTyHZNlR21PM
XtPFXtwsQUZ7Gh2nCgnkuUA3458njRLqkbmvlBmqvzrFXDZLUdGoae0VQrMoGhAProPP1fOVc176
hlYQIxIDMuIj2J5gBA99kh3TtAN74hYtaZZotaCNGpJcqE+gzXIXZ5G7dBpj/VrQtnNcRLkkhPQu
eGaMilTD7dxNM1cxz5d5EmRkig/bXMoj6RXMPdIsjjNvzBsDaYHwr8FK5KCbuVKycrCeJrN86rVp
8OqxtM4SWfAwoGGEI+EyDfpI50t6wxy59NTJSsRfqi8s5FCd5wW2iGKxnbFvUcQ4xgexzIzoHyls
0Yr3iAHWdgEX3Z4RYWoTphRGl7XCGBCIloR6/y8zgbB30nTQXi5pGaAzVaR2b9xNlZ8joAGiKKKt
yfUz/Byjgui9EENm/3lJ/jCclEq15zqa6Nc7uZyGHl1BMJzHj4F04TrQj6DkWPE9jgYzLpe4QppL
myMr5+RIU29CB+TR72kIKub0hgTOnMdVIb74QSQLvU63oPdQ487Vvg66FAyxtx8jt/I0X6rC7HQj
PaB/4bpJTDHhs6LmYxKKWjDg1uAYjyK+MgQFVBBXUzXJkUwWlMecSB3DEpWyv/6S8A2ngn5yFUji
lDzJrvm3SWwpNs3cnkTFJc6dRuZCIOf1w0H77A19u/ueQBimvDLdK/R7Vm9M12yVAIZp5iF2du7q
rfK2dM3A0kLCx009cFmhbJioZY3ZhiYXAyZ88Ml+2QMTcQVJKiOfUZ2AS3qKtmmSCexENh7H1v8H
Gi6fxOdwCvp/YPPxVxB1EuHS7rseghMQphbr4YlyaNRsiV3rUZ0JaKT4JgdDyzyG9RZDcoBGN5qo
IDTzAzzbOPChrYlQ9vCjms1QUwYM8TNWZsBY5yGGwJ08Y+Lf9QLSlRQY+QDTu6jWX75d6TqApyxS
GdH0whvsH9h+/2Fp/nPixlnZUEkMe4KmNIOh8SPy6G3ozUmiYAEk/Y0JW8XUmpRHQyTetVTqby6d
Rr8azV1lE1cCy1fZqzG/KuUWGD2RxQywDP8qkD7RtqlijavIXc818dQ96DjjtMRkIhLgf971M2Iw
I+9aq2gcTd5fQrkG7qR8gNwEisPTZszqdn1aviYQSN/iiXhaQh6xa5MZ/45vtXelkE7kAgHjk/fE
6fvseC0gMHVZKy+y79gxazBrnNyhjXLGyg/2if1cLwGYMFQRBCKFwsLpeJbcnEy5NUwyaQEap+Ic
gJGw5ZwmdOwNCn6+dodzLPDV8kiZYHdl9gPHHtiJlnEj9j+8lriJq3omtRr288ekBwPtKmRK+mUN
KaUgcku5+ohOC6CpOACUyaII6OS6jYCKSlnkMkVNa9AAPYM9uVfdYXhOMljPu8UDDvMGCvPmGWs/
cLJbOq0QANs9dpwb02M/jLgKnsYp4JT3zDQ/r1+zUItann8BeDQXh1rwaEbF93czhYJuaCdS+uJe
t6Sya1NTtYhEiUfmrh6XTPirPACE50QDEPV4ZTGEE8HDrBr8tPU4ox3wnDCege/ng7lvP/37jR1H
23DwuPhg0VzMtbm8PtY7U1f8UrPdrmrMzs6yH4zrK0rM03VQzVEKsWLKMtopyIV/LBn5MNoQrz4A
LWl3wtwsUfM8Lkdx+CwmGCdKX5B6dmH55LIKCbJlD3/jHZuIAcrHseonTIERnozyZhcVhIgZE+7N
hdb8Wo1igSGwEa5OPXrtqvsOPHNnDcaRaRMtG3+rJpV0RIeFA1Lo4s5EFVrGDRi9tO8L5oo6RT3L
EIGGn6JQBwt/ofh/oEzBfp9XNzhgEq3Nn7IQPyxwatinFm2kX5unqgSAVz+lpJl7duVqaYwNlZCs
YZi25OzY05PPc/ZBC28AShQiOSd6q9xusj6n9YUbVkyimVxbfet8xIDVc4bZzruc2eXAoCC3HEDH
uChyVafa6xU880Isjw9TOgqVR0xCuL6qfz1QmkdnSo+8JRGwzCU35Id4mGJEKAxEngjrBNBeF07L
eEa3brsRVy/qv6mpoGZlf7qSIAzQWOQt8yauu9wcxQme20w+ZeXA+0aNZw1R1WEWqgQHV46TNvEw
jKuE0D1juAVTOFx0IViznAL4lAy4tNiRXydk+nIj4bdqh48USaejKwiOZ2fuMo5U74uejNdu9KWD
qrWuAwdBzfJfH0AcIdPnRnHIO9shK0kkZhlvuZEnBLNSdxVwET+R9kQ7EaXLdDPR26KoFCh+KE7V
psMonPnLmbsijFH3bS1lAuHN027n04zJ/AQeNHQTqPt058qyP7a3MUMZsxsQdiam612lOYaYBSof
/DOnQkC9qrOElOxqHEUKoIyxp4FsCP9tHu7lfGXOlQOZaPbOdGtjOLdUzeRMZ46cpALalRtAbRmD
w+oEcO2FYPkRXUrc6eyMLBlEyMaV7xBkE65JD/HoCMGl7h9LdIfMUylAVQ6O3Ghfi9AzzH1KpMS6
b3aXETGNY2C8EhDxW9miWLTJpV8moH6lNOLI3yYdrxLxLPWSxXx1Q1YXaLprUq9TtSGJI9RoYzdP
+RmjP+CCFBbG7v96b9Z1ZmF29ZwcCkoXeKOrtwQqmRj0Qv7zu5vee5yFI92tc93R7ZZKAknrfuCn
prexqskz4/cGxLbuFqSz4eav10/5eOPXm4Oe8WcdZrl8ZpTKBu+JwIlN6hLtQ9AH/25DD6z9mLNZ
XmDpnrNk2AK35sIAOL48UuUyUWoTLowjOPlL2IjlOGizEeAVUmz9iGvEjZeUKmoLkDaBWN5rHulz
U5IfJKSHiCrH8kO/hJHbgRKn7v4CzL4sJkg3p814oCnPtl2Z47yblLyY9mEdAk5A7WVy/qLxVote
wzHkYStlxkJklW2jc5Qm8UvjIriCoay91V6FAjMYL2uiHUE5L6W6uR0kwCuDpW9YVvUjcG8kv3Az
yFyR6RybynaknJhF0nSx9a/nCORwYbB/CjmjodCn4WHYac2t558qScqug5x/VxnUWhFMBrvYuX12
6V2i7OKzE+E8IFK+Pu7NhuW/QR6ho2SnIk//00vk1wR+J2retMw4AmJ3iurOAQPn8P3ssVRu+HzQ
SrWP50Qusp0WzdJZKMnTQSdxEQn/lRvWWiA0ZjQr/fdKucL4EO4nr5CQi9Q7B8lvbVZ09cdWLYcW
jQ7ZiFMgEINVxQ+b6iUnDzxssRT0iWWYa/ybUD9oEwVT8Y244AegIeDwUVHjduhUF8+0axGkehbv
l4jPv6kgHVVn0JwU6cvlLRh6LIdhfFzbXujxJ89uto4joikBNj0DB1iAZoVFjzk2WhcgS2CDhut7
G92soBSIo3BjKJRUmO3K7bkf02ENnJ5fD4N/uX+IohqWJjC+fTsYC+Ms1vbDjKuXeuj5o8JwPBv1
JZhwS+TeHzLZAhcaelWL6X6TEKrY6IOmWzV8jJoTNxcBYWtYgabQv8X++B5f1Y3ZqO3Fm/duqowO
tJCZQojUC4qVnh21cwAHvKXyveJc8UrjtDy7KC4dWfT8N7SHMjYsCgj7zlymhlLBQlmo7P4oRxVR
xw4ZkXMsliQDZmFH4LxLWx/oMW4WYk7zk/n23u8FyIOnGqkCWgW2cfCUM0O5zZKxSrb3A5SAQFX4
Fij2huHLUSbDLxR50aDbbP/lDeOABBZijRsJ9gGtXxh02x7Wq9FWOMRltvsxtLV2rdkl+fry3N6f
8+OF1bcITClZSF/aR5EQuLTflspQE7JjfzYBbd7NVaIdruFgcUbBRtg/AxgphKgoBAQk2ksTOnLp
MQ4Lhn6K9vFu4HzBV+y8FvKH7nTdXVPH6r1HWzeIFTXIRIaUgLoKK0dMxoA8BUj7VKP2Y7+TFsZX
eSeJAQ2Z9xEC9SIX8tObfVDuKI/9YKt+htzd/D7HVpKQhFBO08QgpUpcLF911B/8b0pOY6E3wzwa
0I31TLm3I91mzkbOOWbN5qPWaPJxuYH0rBWrI+4DjbhNC9gYJ54ylgq54VvQgdP27mXuPX7TjlUH
j/nNt98WkHTOqUyMNWk/XdLC08iiD+461EL+i8jquGAjzc3QsBoYgFNYw6d3YFuhVXCDlXTasiLM
mbU34EMx8bqjheYXtw5w8o8QkQJjwk2rTAbPMai/IWphBhaBhyXRvGv74Vtq/jOyAbL9nYhYso7J
SJmo/+KX2MJDrh53FnP1eiWWXhS9h66aYPzR3NZ60pWlXX5Jt77TYUUJAzTyIcZyaLGJXrLKDHpo
O3hZwgsMCGP8YJ9FJdiueENLDTs4nF4EodhUq7zTr7sJ0Mr4TUWEsoJwl0i7k4vswXludiGNhdIF
081jP5vguw69IiMnP3rM2+0+uefUy2zcUovdJhzl8pwjSZn7z+k18X3ySN+YoJeEv6Je7m170Cbl
AZcKaJJMv/YPUqF+XeRhQf1Kl58RknCBiZodpPAjLvfxdzmQ/KSOoGEmEb5DSA0ZvSTqw9biy4q8
KlBoXKt5uajOlYy6RwdxNUbljZWGAc2I3TAt4L2VHJS3AyCxz09h3RudXoyE1YfeUCaH5odHSvEp
YL6gTkx70Fy1pW/x+4+F/sS9Ywi2Tc0bxlM52ZNPzdITS+NUnZgLRTTz9os4TjchM8kNnEiIHzzb
DQPM6ESi5Owphpojcwiny7dKQV0sGzoIu4q/lFoQiz1z1+qz5b5yfMP0J7bIyoUjl2prHpUrfQCX
/qdsejZXO69FkV1sQCoxur/jgNT40IPRWT4lrjuI81ibxj+TdJ7/Uw/xsYebfMrLk1Adouo1Ejj0
lMN6ApH9IG5LzkXdPJl/jSwzrp1sZBgp9H03rWss5Cb7VFVcGKPBHpkXDQtyqYTkfGE6q1OOJ741
ZuhXcIcEI80CdR9aytOAYJWcWs2A7AMjsuIub/eHM3+JFxKRrpCWF5+t7XGtUlgfhLyLTjVipu6o
g3UGGesmXbreJA859xfvmhzZ6HNZVNb1/pPSl1Y4A0GBXNqX9BdiFcxuvTVVI7GHbcDwFOo3pxny
9O0vt6uyEGoLiG3lw33YAUR05m7sexsS7f+NHsiA9qnBDqY7fbPkbuA5doBhSNH9IPHRYlMyjqf0
uQ5KBLfqjC7ZWWrSuhPnQfqa6/jOKoqy1kBlDXTI1v0t3Pxx6cwUULQP7ckW5gOz8aHomlGX4Nff
Klh27dFPARPw+M+OjI40jK/EPSZfe1yYWH5hjUjD66uRIOCI2gC6FOcr9ad+Y7RXf6qTjXfZwdJH
he2bh47Eu97wu+8kNJIWBr8fC57GHirzabV6mu357eJcw2kphRym2egX15BVzYSUP+kaTrnYTij5
xwlwjXTaWMv5wSLnJp7Bv9rTZRBN2iBIX8gJlVIpgQW02i/HWrcwmHlI5/hCa+5SxeHtKwa3PggZ
dR3vVzOlp+8TWglvRakVwIyZpD8UApKWNlBoC7f2ogK2AfC7YBUtj0rQbuBHwmtoQbS42LpgFKYv
l+FkBWgIgmHIrIPlee0S55ME2uDJgsKVMFiLk3QpsapHKqw5As7mG8YUXb41St8mmf0gZ7QPK6uI
tglnbwffw4IHen9aSbmgkoJ+AEBJrRCRbDYHlu5ZtHQtr9QPmM7KPi6vKgqL8dSXHh+YGhMAXdJi
vOIijGBNSc6lvcrXMG8Xf3z+nru0tV0j2ci5WMxgVSoeCuq8obqEWX7z7q1GSzrUGDrnAkpnTVCq
PIql7mwTAL39GeGK6YXIIa0hKoFClR1E2la0sYM+1sVMcevbXRyOzC4oOaCLQm+mJvPub1AMUiws
8i2LGeVLbGPH4iaUsIv2+/HVW4IjiQeej2f9QbWec8ZwegQ8fBfQw/UOEVPF5N6gY5cyyA2K327A
Y3Xv3Po16UBooevRCO0GEc4y0YYUIrrGDI8mvSy/kygEshyntKXG8rVLPSm0UfZ+UvMGkCUX2DJl
LdxPNXcHv/1pFQqA2qoVadTBHAOLVKXvDFRteO/tuFxNlOb6Oytl2FrCw+zHWPLag8uGdrRmgUTA
dLJqKLgFOcZs1qexrAZvKJ3kJfVbErj+8/KF/PonaJZXHbHrki9p6tVeBL5BsG00BGXeC9yFm9o5
tv3P8QPakuhk8HnPUsWTU7roCYc3CRle6Jnsf88DFjxzF91WdCsAsfcGIl+SNYXWzxkVkModJ2V5
Ib1dhifHh2lvgA6/mXUcX3ByAndS8+8/FODcBHsRqXyLVeF0Psi21fLawvMhWG/4b363F3VTGf5x
UHZ8CbKDQLD+wZEOf+VntmQocbsD0m5gb+ZfT+CPlEv0t61e3MTY3yi9Aug3i6xrhrKXY5jv17/n
vkExrZBNnVA4LjOdzdT+wJEbHGi+iHCZrOYPbnK1uewzJJr3b2b0M9qcZ9DgDcdoDGFBh4C075hT
0OgL71+xEXgf9sYO4QuaHQ02THmRjgvPhupw4600CbmbYO/H2l/UVGC4Xm8jojSf5bj68/F127+K
iglBdLfPwXaBRwC0PtRB/F8r22pP9vPVjEMHQrR87YfhOmVZlGDMK9bTn0MfJPW/aMXpXdHOgt+w
ZLVdXDHl9xL1omNbYyFqkqJnuLDdK4sQYR0cBnHqZexJwzO+Y07l074x/o9Rz4RuxqGg3d/eNQ7w
61srLRfNPaelzDeW0L6WcpWtaNCABEQY2/6j8nuPAA/Y0mUcWpIbmSUCULcqJBfJP9EO8io3Rf3V
ASTII9J7MEY6ZBwliUREl1Vq6WfdyR/qyxOu0ff5V5wbnx6zCDzha0e1+sjhEFrfYRfXI40XU89L
KVad7fsmgvPPnpKsgtvZ8f000w7I1KXFL3V5UjnpgE9YP8M6wQzolXi/VfBBUOl2OTs7ujp8wkhr
yR1owa+DcuMbqXSa8Gbe6igNlBUKmawBs4dwzJ9uHJCWilBCtjWIjEbBjkiZNpXeu+DFm3U9Ugvy
p9nId9UC7barMRlreDV/5WT5X9gE4LwL4Srmd1Nj85oqehE0hCnemmExbAiqPJVTxhzqsV5bBwhz
MQitTW1xR2YiGRzwJjNhin72CfGpak5+iBCFW5KIBFR3ZL+CJOAIoiAfbAmvWd+K9zTMj51j4yRU
pMGduNnXDgVfCnHUTjNYjnkUdN7KaGdeAtMmyMOEQQQI2v53digZs1yuD9xHEY8RgVSks6sFyqTi
otKANlBea0phnorzVeutU4y931b646lJzEiSQ05hVUHgDkoRu9RZ3dY28HypPb0xo8O+OdDHGC7A
b8GNta4M5AA0vunWJaRCUobEJ8dFpS1rMF5i8f5YAKWr8EVaIdbs4iRow4y5nK6/E8a6pSQp5QfK
cUrSr/ZelUyMKA/oqV8chd+HPeolFWyT9moJ9y7FML8fLh8QeimvyeKfdWxNy6vxPau/yDl8oZux
NqUMEVVRJ1UOEoGdEupJrZcDaKWHizv+7LRsS5SM4vMFaaPhhhaGryFGtdblIgfH9UB2fqYod5Pa
uIwsN20TGwbQJg7rrxl8u6J7jy6+vbk8iA+8DMoBxxY0B9cdLrThBHDmDHsoh1pu1Pt7t6ZACOtz
bZtZa/4/NqHy/Ej4kiYCYAZ8b+3jqgk0yxueNq0yNDoVxwTLx3qZH8PYfAgM4K++zC4NjYAQtAPJ
QRAzJBTXP6ocqQf66vaILFIzAiiXWvtf9FP+Jn0F0N7IvF+bxQ3vNzHwXdYhKhhKPSwL/gYB34IC
gf+ZZWbsCSrQJYs3r0yAvqRKaZCzRgjkoBGZhEaxixVWsxoPGj6HlvPGbH/dqm0T14+mzs1y7neS
/UZCxihhaOiWm2fMWttg96x4+9xcwG8Nc2U7Fj0uu2bhqm82I3X8cvAhRvgX0j6YGl0XyPEVM1yw
ejhxuGvnCSySwAyhru07e/JxuXpYn1/T7hTXayFQYjPTgAhSPCAEPsEdw7ZibI6n4TAvFUM2rcE+
cLz+JfWZwOLusIIK6Ue/J8ORJ5fYlNtBq/8HE4RLV7OFmr33uvGrfsvGO6kgee/iYxYyNGBExzmQ
vIBFOCxvWHfUB//d5SMSxxuCToG1N2JPPRmMQb9Y8DXoR5CRHy3Rr7N/7UG5Ag4BARR67cJ/b2gd
xbg8swDIFw5L4hxetc0e0Mwzt3GlbvCW1gziqtxUKaSiH1XHZckYrVbxbca6MAES58GM8aDAK1Nh
V25yR8VibojekSgYJONr502Lj2xcpSIVFaJpQHdH3eiB34/BUBa6KgJo4eXyrTJ/ERNGBtHY8j/t
Aosyveulx0FvfYOR9VM4/VcwvfEzSJaSDKHllv6pg7oblvaktumKMhkKrDARKYEHR9UpIdeuGpsc
gdOqv8TDQFoIBP8Sq9llIvW5hGMXQ5H66VFMptGbkIpuk/ajUrzbjhv3UCZXOV35FeVTPcqeGTyQ
zJS6KqsoG9WVmd6KUrds7UlQ+7+Ud4mRbf1MZ/iJnim+MsVVBhqrlmbbdrpBSwTGtY9D4dgPTiKS
Jneg4140J7xQuccbSg4FUGHOjXmvxdM9sR9zxPIoPBeFI+IpbFDY/Dc7wH/XZ8LPy8mgYNVf28tP
DgTNtAcR2+cW6xkczWpfjvVnT44Lfz2vGnljxF6/Oh8+lvonQBycBgX8x7CwOKAjvJGjr1ThC1KW
LHN/3GzflySb3lCSgyn5N9ldCduhwvDYcm0RuVT0geIVnmM+6AbVHni91L3xI8OUYg5yBuo6oz1z
xbfHvOuRrffJuEiuZuvhkpG1WwRqdqJKQoJc9vqMZ3fe3UyMxjfPg6SDumLnRKM9BULee6Cua3ps
JX2HhORxl/rDogFJzJRbuQQcaabiKrI1vKZE0ZsRyMsUH/Zxulcj8K3FGxFsziMn4JfC2xol4/MQ
0FvwzUqvMe1A4d3g6hLfp6qpIkFUR2ewOPoT9C7Vbpi1MxugavLSPgEupfSuZ4EVZV048mbG5fbb
5tyq0lPibopUzlKj/E2Jd3XcxZovEOeRCtyxDJsewnI5c+74L3sqoaZYn13BVPV9Igyw7jf+e3q9
9+3GXfgevfPA/fqXQ6S1hMlUarMLash1Wir29l6tieSexZYt9Z3r+54jZjjf3TNu3w0b0i53M7t9
+fqmuDMZCqDHKR13mPmt9HRIuBqiEHm9LU+jLt7ZdpMh8k3hI+zufobNNjQp7MDScRAuzPmjMtAu
ZbyeqVHWrZ4EKc0OOMGRQgLa0klUGgjfLAjUBTqQaMHJusAJgp57mRRwwuXu6HB2xh1jR/IlNg5u
CAao9vYLBq5AuKz1EAxWVxTsiex/is+0jZfsLzvLH+y2W2okISon8NXV970z2Pe+EBo7HZVChXsk
lmjy/eQvOtY9e8DAN8JoiNxVOoRmfUPdBKgYsS1aoKlfh34NaTqjL4fZn8dRW8GToJS2IrFsMtEF
DEwAtKNUZn/mWSEqnVTYtdNQPEmotc+2H9pVdrWWCWJhJ8S2HQfc/CmdFmTLvqJ5OOOQ55rEOwtV
8BTBCNKGwJ066zE+2FhVWdx3dEE9Ys3IQnRER9rK5hY0JRnXaSAGqCz2cMMp3ABCvTrqQ+Q7tu38
mcFOlRTHaj8QGbG9pHbeQ4PvRORUuM5XhTYaQUf7VB5AVtPQ7dM02OanOJ5uIm0/yuI0SMrXSz03
dYamdtEp9MNmY0YdM/PmbTjSIIjjrklJ0yzf4/DQKckkzsEgivJjRnVHKZh49UI1JfaSuno8s7yg
TH85BquhEMNC7Zyb+ed0jdUdxN2FXj+MtEIUzUCcfMjfEUYyg8Lbr7N4ph/uzfCStG4+bdMO10N1
e0pQS0tjR1jyZJ2BgUfPKGPqKMUwWc8CIQi8geb7mLlEtbFHQ6BDhB5T46YCEdDQuBmWB3E8/kYo
kt2nL82mt/Mb5cjf0x3qmOB42cEmP7bV8xl7i7Ww+iMTfDIvQu1fqhwHMOp064zI+2eFOVcaazk0
pgZnE7GeEw+DXZNfcmZx+M9zENTM1mf2ITGf3r7uhX8P/lT8kvA3pCFVohWggWZWNZJSLqWY1akZ
SKT6EyxKPJvqgFRLHjCN2fo7P67aWkQFodI1NyesHXqsvruXlFfha+qj0OEsmcrPWYrD0V+begZF
MqnAiA0mDBj/x9S40FV/izqxC9PqF776vGUkP/TSIzguaCXCXqSejIVzAy1j7o6KaMo34xykVXfo
ihS5eAwDMVBdAPgFM95qZQ5a/MLUvR/IVNQ3dF1AqJes5oDTrc7YX2ry6s+iFrcFx+ARxQGH3Hb2
ErrDdh4hkdVzcCxMFHN4kPPNYaLBDLx9wnXYhcXaFj6OVjQfAVAxuw+r6OZ5k702825jJCPTWiRx
/FYCRa997JzWMW8V9bxF0Q/eYdvOyUiRI6eyS+ocuhxLYzTQpPIYfPHJGmcc2FThQhcW5bWKr611
gAQeJd6H43D9M0LnUMyeD3k030vESAfmbH2P6b1D37r/IwqFw4s7/x/kpXoIQZ6RoQze717159Aj
jlvzcA/WAq7YIufcAcO+sAz/GJdLSuHZ6srNd09owIZw1+UixhUYCuj+9QVlgMEnUP8WUvaxsAqY
ecHZTfVao+mwIfE+1NdoIfCVfSP+j1cu+qA4hpg2fy86r6cy1utFu3o6y1CPderPYeHeCTct/f1a
afbeVRa221S7fwzVLO+4CWTq+l8pcdMN19QOHSRAiBU1f40znMq7NYvlILmnAi3GhqazMiT/uus7
/e7jVzneKOHA2gRGfCIwcOJBJV0pLYQqYIkEMfOgOh3yWoy9AnkM4V47NJG2Em3W6LtWqke1MUL3
9G19r+txUMkqJxF4F4d3TP8jYx2JW9EkDJhaQJ2WR1OJY0wha8aU1I7tOGlmV7E5lxvM0s/+Obtj
oQQ8y6IKeJJBP5m2HXCafgnt2NZR5Sbc423Lpv99Pp87LAZd1HFrvKztGVaaygyRKzooNcKdvHpc
yHCyFa8CMnh62VS+92jQbALuicSEH82MZkw1tFXrRZ2+8rghmNqx4Km+E0hGmP1JNhDwHVIYKQg3
1AZI5fwTRGTXo5964tVlq0aW5kTT8Y6UQCYiuiDQkdCbBj+j978bWil69GJexN+/vZEIP+OpiIil
xj+Fr6s8JIAL1PIeZUQyZxlN5RuQrJwuj551Z0kPYTBXJpD4Pjuxs65PtcxyHyVTRDZeHFmxBKBo
hTRpqMenr7wHBi/nDvjDDH5OsANDnRJOqgRwCH0jTbs3fcOa/lG2nwhUPPaDbK1NYW7zUxJxPS6a
PLP45QygO7EC28CXHDzLynkjGUJfvM+7fuJzQsPgj1eZG8kqx9k2e7B6mXetavUYXkdIrpARvyO8
WmxVvmDTqoyBP4jez+VIl27wEZrPecEWSmwVPYNjEb1vCrX60XcyfDK5aGJHm1u8RzVTtIh7Mbst
7usvM9chQ0RdZwBbbZW9gdHTCGzNJFe7y/x5R/REZxiYmz8DwyRpIb7LWNSXGARVdUIXUICqj7R6
v2dkP0ttX3xWVL7FIQybiUWVSow4AbU17s6AduDSnNpbcNjmqeqzU3nmWzhvPU5yM4p+LUjmARsB
oMiDAjisSwRGzjoDxnDqXmB/PhbFWJm948YSjafCHWH/wrH4JNQYooNoBrHRDN8B+w4PG/4z3ckh
a3cCo9XZQYwPQgKChl+2QlnPIMtaasX0HST3ymDZ8X9XqKiTJyqjOrDKoxgmQU/vCtCYexZRMzwD
Xc/hQ05oqIqbjjXbxscNuYYsiAgUznr8yoQl22cBRgPaOCzsb02qz96BrB3af9RX9d/ZfygKT2zY
xuZceVHyCJmVgDu4DgOOdf34VyBwWB19MCIxqTfNxUEvzVD/mvRaKzJYzNfYisp0bVeJuE9G75xo
p64asPEJucsGE7d/F/2jciEVg7ncHvGjeUpPmvw77wb325PR/xnl248nfy1/qkXT9I0jZzI6n/f9
lHXYqSn/vZPZRgg8gdfDIYBIRh2NKjXRfdZnphaRIzuOEi9n7fURgpqVOvc/3VljcFq0/amdYwJW
chlo1ELkYp1QgsZR6Im7KE+/sGG04y74lEo2HAbj0AKo42cU30XwagkK/xbOv2VvdwlKeiIeBKLn
4pDqnaIeXFTfbPOksNGAphb7bnD92nm7fhMWZX/aVUSGtxhZYOaYcobUK2BB/IOkRB0MnbzyFgCz
Jt61X2Sv6jebVQLhUiTBqJZ1NL/5m+e/y1/n/VKoeWFqq2BicyriOb47n3ux3jLS3qjWu0wKZgxC
XLtVQWvdgdFKsNnXjCa8heYaBrq9iB1abmHl8xnfKPHIElCMZqbGxhohSZCK00Qr59i/xnntU/kc
SVcFZ98yCUQfJnMtEOwM8RxUUbYS482kUKrgp5BYn9vYO0UaRIkrzK9vqSbYKfkuW9AnUBaA2R04
w0bsRFDxWLLUIviRs/E66mWSBkW6T+eh/hHPLezhH2x5IIVZXUZSLADRLA6robB3KneuATbIsn+U
oO9hO0Ueb9ucolK9uMciYoNQMiR/WdoyJGWXqhq04CEhHDaOGFMlihSGzI0XKfpbgoud3QAUxPYA
4qqw7gaJrwwAndrInBUjih8fd0fRMtvDJ7xMgpyBXiBLiCbLsKFSVAUuC3nDfQu4yWEqdf0/QYYp
MVrtYxWvtamuny86KoD8M1/vJgQlo+n3YEzyJsTIRDj6R89hkI3dfC5Qbnxey1hx7Pyq188i0qSb
Ji5MdClHkGmTjng07R2b/U9kMRBaKsn583HRDNvkiVxs5mJa8vhN/iNIe27suKCfvr4PAHWYn4iO
Y1ZOTGUslA9i0gdMZqO2qAn5o9TiZf2M9dca2smo4l1Vns3sP3mGuObEu7wLDz9On4pt/3TFxohZ
DJi32YIFrGfrpmWSdmHQUwKmenfW65GEtqCGKaDWmunY6qPbEuTkHfaXNXZS1hnrCcbKj/VCcI2C
j97PnhB4YQEtpN+/ZvK57Zo6mIZFWjwjCzMOxAfvMIYerAx4h8r/aZkEqiNRj6NP8VKzhJEmIc6L
Hs5z6jg5XzKykyPCmLMVQY5x06K65NAief32amZP6GXiHcbYk9FOdQJIN4BnbXLuxqQGkrA8nGtu
7nfTrGu5/1aYVQLumLomK4FinzswP+B6l6IlQJ+ptFK9JRt9UP5RSRt4AYgzmycUP1hknByxXij9
XACLe75bUTQyi5hEWrRgs+SxJoCqn11Os46rD2/8N8mSwZjbOqSDe1y6+rGVNoFYA2yuwuD4rL6K
qGY+tep0zsTI/FBJw4A//U5OJkVc7M3LA0aqNZY7zw2LYy74VncdyDln9Fuz5KtZoRT4q83g0CiC
D74DFoc2J8yy27Kf3Y2fMhtY8zCtZKwjLa+GxPaRRFr44cULgMoQK4xsbnzIZpSYJA+zUAicCFLP
K1jfadgla/1Tx7818IECpFDfrIHSyhd/1iXFNpGFqPgnkeBgTGip+Q53McGJOq/91Ew65XARi1Dx
gq8y9Nj/4+G+YvRcAOrZ6rnFmC3IDzOZJtUy8fmgGeCGTI+DNrM2mU7XV5X5O6Vp4UastVGZ7V74
qQQOkviBrzjhd6OE6o1r8oYi2tbl7ZcgUNBLvUvUsrqy5fJwaZvY7W5DD+OC4fRvlr6E6ASV4T56
IHnapqthlsZn+arD06i1G/GOLaqUZFFTOjT/MwyBCpyJLs1DDZI5bf3KUziYIKOFkuYPuumYzbRc
U00q/9AS89FFhE97MRfeh08KX3UOnEq1gp6oHbAHkbRPLLi7U1SPGr9kbrSkSDkjW1PW0Zacd0e8
KYA+69H8yyoYy3jNjRh8M0qPaM0LB91d2pjmHCBYw3voliaUsVqrnv6R3rhMFf/gDrwCg+nSX+Uk
2FAmviGFnbOVtSgGx5a0Sq0f9FGbVVUrtChyoRvpNjx7HEOyvkesEFS6Cn0MSF6ou7YP5KjY8wlt
4EN84ckMBoCQlVJwMWT4u7OX97arAdywKW6/2yADnYaBdh3KGmYQheeNQ2i+YcpzDoNMcj6GBppx
72Wk+/eAlOLF5RyOF/lOsVTusU9zY/Aczb8cFn0Qb6c1dyFRcL0YKGRLmGDZQwjP7YSq0d7q8Qc1
23TPGlAtKNvz4xRD2BLJQdZqtxzpHxBzgQ1NgXsssB4wRoocsW3FPllWuhANB2cGPKJthRVZ1Lm7
xvXvW1nB7Z/8wPc87Q52WXkUmu6QeAe/GuKzIA1ukG/OOmgeQrTiBKFDTgcSZSewowkfBg87SoO0
A8CyfRNjs6NNk2ndMzTbEAxISLQ/ek7zx6W+jXcdtX2dEGFkB57xoNStlB6hDRadTlyCpD6fNjoX
Cin96Ii6rCIsnb3MWD+UJr0ozxB3c0KEtQ7OK68ZzogqxO6OoUVHnGouMgMCp0JFx7dRvta3aflc
ypztm/mlw8FoG9BF3/669KHqYe9UwxDUoX1URdUJZW7v8GRx0NgLZIMNaiRyAeV4lo2uCypmHlRr
IO16DBjyfYbg/2OJW6/0r9PD0XNyLwnaMsVDeEKXoUms0gonfEuQxHRDSgYW4vbdMPw2MVnwJ8kV
XMZjkuu8a1Ub/aD+Hdq206nfF7hueOMDOAb63qaUhRJcUYEiJSyHgJ7oCJkKHBN4TCBb/tBz8SKd
EqP8atzkvvBb+HYCHPwZl6VuJK+KloGtOqacm1ytBJb40rFORDxGzoNjnUxez99lgJRUKWKQUPvN
rnceJBD0SoXp320bo8F82sQEWQlv2sfiitX1ppuBXkHS+CXgEvMRpHtmhzwr6pVEViQaf+DXLH88
mAme2z4+P7F5xFh45rXZtt9/+flhfnVSfHar1bgGnZvPKoGZryqCgnTGv+p8iINT3SyF6bAGOHmH
llBiT5k4rMX//8KsFXOAGfvBpzk/pC3QrrsxcWZeqvIgGP5hxNSVCZ2ckJ7cMEw5PHtGzDx9TImZ
OtWXtz2qZRyp1ICI5f5fqm6hjFU1nfF7AZAS/4Rgl15s9/dxG/K422BK/jW4i+sTjGIDL2GEKz7U
XFy59VsNtzRVcOZGMhN6jH/Rg3n/LOfKRWLsQYGwCRK+qCNW53lzIWS31Xc5bshsKraMbsgRSAJF
t6FaSUpEeWAzsuj8P0BrB/bd1m5j4LZ37QxgAuIAnvas+ncjOXRHrnRzYWq1FOqQLu6Zk/lRmYxK
/wPMSho81OSS+6Bd5auraDuugqsH2rKulnt61F9ob+cJ7ki+R8MSJ1vEnteQQjS2s9Nc5ABICh3J
56Yp9Y4F+JPKvv4+ghspb8r8py2BJW4CXVzgtMcuMRb2vXcA/c7EFhMTXGjCprPg25f78MHpHYdK
pEmJcRlBCMuPIqrsYvPgjAXD7/H1qKnwWLsJMyJDwONntatsY57+E2tQV/+hUBWA9vxKK7/NDflT
sEeOvVBN5auWUKXhA3PdYltuQS2dsG1+ME5cVbc5u9Hn9dfOfT0PeMNZO8FKjYihhitgyBHtkqlK
GtJ30FTz7L3WSuHnijD1MyqXkwcknExmIZLeNuswDdHVGcI48jmcgJq3ZZ2m6Thk8MGr3wTMkenW
rmdxAMPC7b7Atf7aRiF0TZecWQkTOKmIltZHjJvOqUGaQrKTUWwjX+JpNcT1OfROGSUpOICZEzRO
KiyqR4VAVU/oSj/R2acjANJJGKl4FLqeLlvXnA4RjyrKUw7HgWW7O1X4HbDld70c3/4SocmRGpTZ
3o33CTD1fnGLQb0SPSscNRvUqKkRcp2Ydlx+89a8ROH9eS+2DNJirjXpENVddj33CnvmnhXbZ3lE
ccPcMDQXLYg+dgkTPp7g+9RFFmpYA3nFEuD4uhTB3Ja2n6jOxUmtTkTc+2hxWV+suT65v86Nb51i
Amt7Pv2lDP1Qv480HXEyMTlOyuwfqCDvx4QB0sWLxYw7vqWd+gQLaaDyRxcNN9ic/mZIQJTctRr+
6Nolxv6PXxe+PNFIaf5n+SibpaCG7kaLFwpZwVX/Qv0AsMCpPMR/wQ1FpWx60Pf4UVSyznsbjtX0
4/VL0rcgx2tlPaAVyGmE159XMeVogRAOuXHyuMwmQScQ+ThI+GJfLhZwgP9lnFgPxUuMtPVfp0Cn
ATgHnIqCzJIWeXxZ+mhZLvLnIV7FD5tz4WRNtlKzG8X8CVTsFag+XLjZSalCyy8kYJLsnVTgtixI
96RK5NR9ncenJlD5mBopkIzN+cv6HQ9tBisU6aCnhqyL3CMg/bwh1OApZlpW9jrQTGkkJNTJhaC7
6z+GNEnH6PmFtRz11akIg0iWTB6kbb9Bl7Pwf9U7M1Sd/qQSgex1ZZBqxNpIJzn//X6ePheKgoWc
M6SyVcb9RiYnuMHywq1g2OF+7Gi7KVleQyFgxRIA7JFMUfZTLIRRjvzF7j7myImBPGXIA3OMX0sB
AEEZZQw/W7Tk33ee1BdTEwQ2Ohj0SbgK/HHmSGXoSj3qIVTTokX3o5GKPyM8QkeSoJkEdqKn+cEz
SCsZdg1xE96VJIWXBMMqNknwFGYKaJTOmdNqhPwh/0ctHsC6Zx7/J9hc292jsiSfnHkASoT72iWS
5HlQf3Ham6MDEdApxkcOZ1Br2IepexcUy40jfE+FHqy9G018KFWf2vvfm7Sx7s0kx1d3knjOvDl5
OsjlIxNz81aV4AbT0jOov2wsluuEDkqxj5E3jwqMLYMhOwEgqU136zdb3EX7r7voPl06UyV6djqP
7Laa7RZ7Z8sFUhpG/96LjKGraoSH/+ZsOIM9QdPSKG3ZspuxbRyz1Yj4YtrLfKVre58ECVXhKKjs
DbN6144f7GkicN1VCe+3td5Ki9nHoq9RGos//dm0QkcM04bJuXtPrzLXTwon8Pi7srKxkBUAKrti
KMybr4tGiygzocI198SOsyZAg9MNXixVmHkV4IwFC0BHdIDl0PEY7lJa/hnAp8uwrV2d2xD/qXat
lUBMNZ6yu1P0jBRD52QqwU90Dde5FjbFQN86CwGYBkSFE9r4pNhk7+gnIzHGZkDiAoQ9PzXBOXL2
hB+/Q/3PXpglJGz5z0EcQf787A0/KuxO7dAt9m9m9NCuwqzdSlxVjpj/9Z39eiDhqHfmJd65MQoW
WXEbBSDsYNoszg/9FQy8x8TMa2lYVMtIa9rSFgAKTXUZ1tFBLLxWeGfD1XCUD15lB4Q1xaW45VPC
Je2bhVuUV505AMVKV1HGw6eOY5K+8sD327o0pRQIJGYmH8HoGeJ6cQKuvjnTRr8pHvnrCeqmTCeJ
xEXNtv6vNeGkQNNsY+GWNWA7k4BhzbJwtfhS3YMz2SdEeMw9ccdzRfH6lKmpihSDqm8uiZVz4Rk8
MBETQHXqqBf0BntdCiQSmW0N7uvCBNwVopdPZ9mR9NZ6bLQaf0vtA0l1+c1YwsB3JQCd0uzpMCTC
WdH70bBz6Ku+WH4OyTQx4IMN/NxEivJ5SLFNyGHkfyKn0D8EqYd9HDWtxFwsQguVdbHAVsty/v+M
tFoF7NtjyCZ4HYt5CZirlnRLAKcZc5tcU4sbE2f3SF+OAwACx4IyxSiJGT8HcYoWznFyZUvLtfjr
aVVmv/Bwnyv8xc3dcmaX00TZB8N63T6aXaOzKPHvRl2+BZYdiDsK1XKQ3JEmIKYdzaPD7G9NRC/M
gqEpqtaN9yR5HxJ7VcLLfsQzS8o7NWqkhAOAqbgnKKIvMuMg5aT5X1yrV2rUmNLwNTUt1PwEd1Ur
UBkQlzVBxKuUZvAYrt0pKIcOaHoZ1jf7U+yla5fIFeE/k1sBbzZQC8NA3blP06IWM4Oeqbj9iv3W
U4T7um3F/unAJzswh6P+JYxfL+TMXF/alExR9+k86PgQLqgzLoAQxepRVkGsWiPk86LTinvc+qCN
fhYLHE0zJKDJma+7G/mAhgc1Zzyl8NWC2r43Wb1hewWUPfM8gRq9XGAyUGsN6gJYnJKhRwboqOrt
vuYpsByPOwHginj15rQfptzTZQoqO+l7R8NXcjNHV0VxDSxwkqwlnJJz1DV4I/toP5I44gbwNVdw
KsVnRmumpmZmy3zCT/M4miWlxNH+IWFNlrcOzWxWZRr0IHx9shH6LBVF+Xb/5AZbSuLtsUpHVOup
nEASy16x+bJ0RMAFWgS+5MaEdZ7jIcD6NXPe4Mi+8RbLmUpp/pxXnTNeq5jzLw+yoiy3HEDL+KR9
K96zsJ6bt6iAXpQ8P26/nSh20Ucv8QEBweQaroCjyKt//xU1nCB7g3aZsaQZgjNRqY+vlrExS7Ie
vKf5aPMPUf1sKaVEn7XDu56+QQnOTsOEdFdxV5l5jay3qz4FClIEgW5QwOvfAL+1tYWdK4QmK2cP
hVEuwlk/mzz5cuMOiVkKb8IictOLFOVWVyG4Pb3YB4FYOwRgGzgTiGlpSPEtnD7hBJTjl/o7DXk2
S6TwCqM2kFwvOwyIv5p6Xm0XJY2paJgJeHD1kvtUDm6STRYGoUp/tbc3inj5pVyfBPZFIzAP5eRJ
tkdDEX5wrhUm1KS8ypFCCzWlgvjDq04BfduSqQkcgndlDDhgWMIi0Z6P/o58ik5zRGZ9k5mQwE3n
HSl2FU3gcoK00W2OOdntqRBFEdlIKqUWPP4ty8vhMLbVhLij5Cj8qCSHPXYk5C3hruNO0FzBOfrO
kEH7kkTM+ZqSvzHvaOycv+6IBXU4w6fTeCrHS+mPHPBR/9/mUYSHMyohvPv2sbGa2WqRxZNdlalk
kxdxl/V1YjRl/rMW6L2/2F0l3c9Cn3kHOeGjyX+tl9K5S+pCwk33FnPZ9h/YTf4GKaoHVzZGstXe
mYP30bJnwXVkl6Aa03Kav31beRBLIW2OQVwtNiBUk7AMzCk81DkRkho3nzmpkRAeL4sxSwuvzlb9
GUrbfAk7ydC285iWvPWRKUW1XaEgT/5/z8mc6YxAMCvz64/22+lK/l/wY0SSlJaA/8ICNOrRCkhn
AcCbqj9rdHXpYyQC06p/ovvZYkyScY/wvbbNUJovaDzEXKb5JmS507PkMMTaNd5Wc18QywewDaLc
yV8MaybJ6ypd1WQ2MKNVFcacmVI0uiGnXtgxaktwzXh2IVvx3lQukoBd5gFbWxzB5jssNxZscHDF
XeacskLVM147fOnB5dkXVh0uWCVH2MntwXnsJUIeUBF+H0/t4ulWienBcUBa425vrFHYDOsb0b3T
MBCgya8O55i6fQjCxvfFjTUcjefyEOGW76Cg2gFsuRHUp1CXSNFUW2PI2xV8+qn7qu2MCFBIkthZ
n1Jz5J08lDSXeyVi1laAQdtgIewJH57C+B7hP4b/jC37yQY7/w0DeLaQVbWc9/YvwZOywNIMoNSU
Cq86fBhmxfIyI9kQhGuvWKCHBN3Ki/qGsxezgAnuY2kIgie1EJ1JyBjF9yyC46OPKta41eNSJ2Q5
qgiAsvYdV7Ya9fpxO4mJrZ4Pc++PAPeS58sAxUVNQ+JxNHw90GSO0W011aM2loe/GFGmPwnrmR8l
uIHwa210H323+Ukydwazm+gVPUXrdt+ZgXTITzIKLdo8CBdqLYeOIQgHC8kyraYZZkEf2MDogXZ/
juaEIX8iDKMMyo+SlNBZk1iO0qbINNgh91oh915Invsf5bNOghXWFQgiNjct2DW2ib7LN7Q5sTP4
ggrUMi79ZVlKxv7+779zun6ppVkU4bPIwyR8P5/h8j30rgXHDqTq5K3VGcIC0QoQGBixHEBouTcB
w9baANuIGSpkMDukQJhZDq56x82JvrkWbBlNUl7DpeMPNB9wUns1+5GhYVR7HDlHBQtfijTn1hUn
TKaCU1WAWmVcUCCmKDnv8RERpI4IrSXFFxQgOxx/YPFE+cRNF0oWFzAGNQ0g6tSJA9Vz2Ld8ZLfY
/A06Myf00UjphI94w0YExGix/xfqeobKguOH2Mn08GjVwYc7XRaY7m8L1AsdAimVJcXK1yPZuFdk
qGPIX/uOk+WyKesvPYLangQZr20DjdN5OOueGWFzjkWKVxatM9czCrBmMfJl6qKVouHx5cro8MET
nqmlTGZHcA1tCgu+Lo1Zs94m2sVya7n2qXG19U/Xv5TI067JEi2TvXRNuq+sIsaMnTsCAP8Hcf6H
OyaDvSnQLap9zFwZEBz/rGsOnLl2P2o2Gol9UObVkjow5Ho3FBJ1mDkmuQueUHamonakN6YJ4uMU
W8UB7fagZTkUAYNH3BYuE/sw+XyapvigewnqgaSh3tuYd3IwhQbguuz2r1moBbtXpRYcq2luLEj/
uujOA8qIpOHk2u1Ne5vsvQto+VVVqGNHjoZS0+8xHYGSe0fSL5LKlRyfeWg7JGuqfie6YRz+xc2A
6wIKkduZ/22giQ/EaVpYeXM0tuRKzlOpNC0LnoDMBmPkSXoGGJEcSq9S3qrnolrzYeb7/ElG/MKk
udQ3jriZ0Xbd/q2oJyoEjykwmOIcy1XjlesTbNSuZpo9tTOmTaM9FW+bQZTounnpPvClezVLJ04M
TcAU7taViNELCBUEcgj4aQFSK9LRPgDRnMOD7pk93rIOF2EXe/jR1i3u9uzkKj83hY+KzcxM7oMF
9faiMqw/QNo5+b4ciJfyyKH3iLm2l69GCiVoULYnG+EcS7ZB/SbuLcE7jDu/JeocJwnVOkhGaBUe
nMyJ0EGtZNT7QmuY1UZokEO+6hlKDFJ7oSW6+Kn4W6vIBmZezMAnu+6d07xst6GifDP9gs5muBln
/vIP76S4fAqTKi86Epu5UelKfZ0hd3O7Fkdf6519VgZSD9DEBL0PCvodyIgwJOKD5b8vFclua1nE
Nd7bbZ1Dh3bYzDT2gHAvsODm/XS9UzB4b7n/nz4NTlImVpB/+6GHoK8EZ5YMcD5RUf0mK7h49xKH
Gz59azYt3f3w4yMpMgiRaHATY/+I5FBYSFQ8Z1L4e9GvcIIGVN6X9btLoEYqx+7czIeFj+smchdA
a5hQ/F4mOOQ5hSQcnq4heeOjSqAcEvFZUeLfQJy64dGsOSjrUOKCicOyT7gLk4d0BhCuR5AQZF+L
AzuTXj/XXaVbNe+8MbwGPWJhtfvmN/LySSvgpUZvU3lg9XQn8kJYdU59iJlzIWDWFp+p1O2qehvz
0juJtmtusPlE8zXPUjhKqSZwV4RXq8NPArTvICFKaoywcMY02MAQyXYql5gbs8d22b+slp1l1Zyz
Liyp3dfIasHQB1e/WGVCnuDAZ8bFBCBcfNnu/HrnJeZedwhtPqvmHTE/bfGIwu+Lr6HwvroyPbNW
7n/HMAAH/1cHF+gpmW0zVLaGfH9am4ZPyH+zjDyUYdj4siYQ/22cOPbow0hN7shWetet5CuOzCBd
0UwTb4GOQbPmTEXM/k6x91VosT3ok645B9LYNE6TscZMaEqYQqk8amUjD2Nt6VNIK4bY3yawbcrT
jC6232lHc7+6t9Pmor8J3uopEe1fgNPDIRCCM5f/crhIoU7ztz7ZClyJxDmoqou42TVtVrQy1Jxn
8MGXmihHdIAw0glT/dn2+LrQrGyrXfSf2UxDXTJMy0+s0cDt0k7eLDj3PcNnhAAtrlgNghOWdLrO
YSMytPsIYuGpKoiidnygeMyzEu5zS+faycNMFBvnsK/YbIzVU9ar/+rH/T5mW9uheLo6/mmQ+7Ta
oILg2thlhR6dWKCoWqcS+t5HdC9XSXtjPMKcaxsPBqNYsmDaxcz+5dZdeKMOEqSWMEJcks6VEz5T
30E55tLPCN1uYa+KmXu+y3qyq573y1o+H3P9wDxNzzoPakWCMFL7GoQSFbelUw85JCmmTPc07Kmx
3Nya/CMTNTcTl67E9eTEw/ulCJJo7640Aund9v+SnNdKEITB/Uv8+AchDD6GzR3QoJo2Z6POGw+/
wHSG8NI6DEi2nwdJkZGDKUcVOlBa7byZKVeaUE4EgyjcWWEAO2ysJgDvsttciUv268n0AKvDFzOI
27FT6SNoo2qKlZxzRoTRY1tkm2FYM2M0sjQmeIGvEh1Ybo3N6C6mY1C8SlvCpmbj79M2OWQKaOUZ
BECQtGmn/0VxKHzEEAKgUne8bP/SZTyx9YKK7RM97ho/izw3C/Hzc3yfWIzzzPIjNCR2o1Fi/J/W
/v67TVM1SYMqEzQjN0BK2oTTlOeMZa25KDzgjikLv19207ajo+hp4TbT7arwl0DTuEAqOXdoB3P1
F0VYec9JpLFys/q7cIJE77bo4Y1SapkOAHh7ANUHN72ysfreO93jsEvZHANcTAA1DvYQiO1sG4LB
nQQWpbz+pIy39rZJ4cZhwFVumV9Zcq7Xut9A1YyEWSCCsRFA+7ZsIWFPusAiUNRnEQaWd0AcxX2C
Lj+4U5HmKe1MEGtWbNwN3UAA7WCvl/Iq0+4I17S4WVvdeWS8k0JtHZlbYRosQKwIFZC3zi3QOf7H
m2QU0tFZRG89AlgDZ8m3CiIoWnKZXiUF5OuVsrRBYsozNQqaukJk53Y+LWmAHHmPCn8DXMyeGtcd
Wyodb50yy2SBFu6YuLKsH60pLQVwwjZUlALZI4po0ejYpqn9TOzDPoKyn8cQco8Ka5CGe7AnNueE
Zof1RfnI1OYhY/wAXlBAnknYtagIQFHpX+uX9lhhApzexOzLWa+02v445culUTEyE74O7uSjsRHq
X4H7lxMFf9sIUW/E43NkP7QPQabTPESgq68qawHsjBgLJh0LmfhJ8Twpdm6EKPwwV9f66jlG8G27
FvaBXsDpS4lNyxW/7LpoepuEfv4OyESkD5Oa1QYM+azM1DnradcK+5zdqIoxHjnWWGwmb9e5kwSs
MTrsY83uu8FjLdTRWo6zhHCcQlzTpddglMC85VH5fAj4fzdh2BAL0j8AfsHvj+371dP/+wSGu4nX
kjWw5mC/abuIa6TL0ku48gw8U+193Zx1tGOHGMZVfEoUXMOSAHliCArGZS19mZzDEJjBBmj4tDGg
WDrEOA14jH/eQT08UnuUOOTpwExzmryL5wIxpY/hd3vOG4F45n0bozqQY+0ZI+EX6gOwmDtMZwax
JjtVvjOWvBWQFzL+EiyU++rgyKho42KmfaJC3rAAJpqyiRGd90pDxVDdBk5OBYzCypZbP0cuCxx9
WEBA5p1k7ykYRGfioK1YXPt9Gmg5/DBml4k9uDqjoa7vLDcly4f7GSUQHQAPjt7ScHaXzV0EKAnC
gDH5I1NJF25JEpPFPppUp0+Tr6rIWNQaSK8vIaUZsekJb0j8XqgUXvR4hXrpbmRT6BNMjfVHRAFc
WmTolG1/CJLx5GN2MaSWt8gRsEGbsyA/Ubp2Q0L7WEq2xIjaSS00hbXUgdrpF6Pbo0xZDcrHCDK7
cU0eN7lRG8bqLev8sKeRVArMNnG3DovWVQyNLxKVnOP4lC3HKRoT3IOd9Mzz5ryAK419DZYXKcjD
8CBDyFpncig+wKGaUN2uFx+h2omemrOXxbIJ2DKrfJbOvGH2gy39kKRZQ1CmH0oky4/4zEKEKdD3
9XmeKkPWLgslY3QCxZNg7/ysfOQmqFeTrmFunc/5BtrfRhApy6eeoJJRH4m5Rf0t8JJ7mEtY4X0j
OiIl4YcztRNWQme8Fb8SOrYz+ygdr7p/iB4XREoe7vmmpf8jBVv/JRRzf0rPzn+fuwms8gsytji7
sA1jWtmjTSfelIV48stYfZu01e9RjDXaIIZXmxdKrWdEGXLSJT4n5mrgMBRcRRgmuXQe4PkuUfG4
SBVIqY4TkuLUdWzYT5SMNRJ4atDBBAURv3F/nemTDXqkHfLb/rAqbXVNyGLr9P35CH5jSiAfm+oQ
S+svJtSSJGKlC0TdDmkFow12ONQqeQ4eH58D0AHRB0947kM5gZA70hKodinZLJ5ItdWywB/BHk+e
vh526OUcBW5pHUu2A6f/ZUXKt+6dhHz581ZTR361Ek5ND3VPZ57tmSu122b2G2eh2qauwywY0Lq7
dyKpBh1/Es5PjJQO38u7M5RhV8BmfVA4cY7no9aFCUpT/KZL5cCP80Aslx+Ur84VA28y+cUV1Rhi
EaJSee0y6HSVXKeYU7MDKeEl7gG+HNMf/kuav3YI1x3aTsUsZiqQGO79l7C44Nn1dcLRXsfHEqUd
xE9eEGZxQH7BRRC+iNi+dV+7rJAn0ee1niQylCqAPCjVWj0W52+/faGCDZnnyp379sYJs34zzTKV
/ANwVcSstzfHR4RR1zHOpBo6PpGGNfayYB0a1bg84R8WiqQFFuGhxI3orHzzDAvloFLASQ62bAm+
WeeFxDqopRaZ3pFIsxW9lbRJspalAhuwmPSpU6Ye3EnUAsk6AlVHQ84lyFEZdfLS6D+ftruRx0+m
qQ/gz8PXy6WLNYqhhXHKr6QYe9U+K+qnYxaCdYJQN/HVvZz/wCFY+VQDFuduEwChnPx0g6fhmkQ2
CpTa7s+CBgyFozqivxaORAOEGn8tZlLhUeQsOQ+yR56AUnVCzC53EuuyHBAP+GRkgO0/b7urr8YX
ECDmTXkXxXsGBVPCM/sI7VNe0AHLaQH9k8YgYRhWr9DuZ4xrka3JRsUWzHNX1WunOIA2MdmrjpKl
oXd393bwdkfdkeEL2h4LTgvjUFDPC7GHh/yjujHmIbdov0bqzqnsDzEM/V5iT8rzrW3SNciXRzyF
mshfVzEwTzPQeY3W0zowtM7x5SR5Ow1xWL7VM54nzSDSPNr3Ob0W3Hkmcd0RoHCEeuwu8rnO045o
DuB+bgWefyY0HJ5UGVDq0Pgp6SFb4sms8pIFwgyBFdjsTntYduFAyRAzrVQhcL3rjeoThCSJwCqB
TQATA5gVrSo8nOIyoW3oli3Hr3y4LETyZSAucXxgtXLG9nehCU1y16qVQt5aFIwfwdi08jtumhKz
dBq0qK7wTWTl5mOEuUYvx1YvEG7PH2ISy3UFCx416Ya+B4Kh62yXf61+uP1jDUAg/lPS72OYeXch
kTewCQakSj4sprnH8HWhTIi87SVKu6lKb9AI3eJdlhOhDiQjNXWS8Dujp5iGzq8gL5u6/g+RLSac
KpQ1wGOBinhwFHHq0JpbG8ZZNggbJJG1IvLVMEpIrBO+5STplF/C49zUHNKlTNil/Y2BzgOvd/JB
3vWDm0Xi/gVbMPv/lmntcbRulI0Va8Z4R+2EB2yeQq+KXL82GtPZGSlAKvDPS6D2Ei9olh5u7z4K
kadcZV/VYIs+fngEzON5uLdFZKNFh4uJ+Tl7RfPMRlfrZHllwsMnwt+RutfubNFrY4kpzE32T8+f
CdQKp359Sm2h1yoU1fN9uOtbwllxW+NKG2v7M+4BukBhvdiWcRORIKVMHrUADfc9RJUgjzBdFhli
ODB9tUCLwDSRhDwCzHitZBGyPt+rDxOtxoHG5FGHi/0OOYa6qIPB6YDeA6H4eAWzB2DatHuo0Ind
DxAuUF1VlCW2vJDY57QK6JKj20itZUL29+wqafA0B4IqLYgIpHHH3nzfaMBmJj6nVWiDjO+kQnwP
9/1RAUxIAGqvRg3JG72XpGGeUrwhObMP6U77X0JU6JdcFMW9ZKsz3Xf+e+mOoClj5EO7iQ5OfMZ9
cpQN9UfKfp5iZVuSqYmc/E5bm+10nz95vCVg+8HW4dxzxhi0iQ3PN6tiZ4PuVRVQzSyOZxO7TA9G
QDe2cnmm1fGh+BVpejIBE23OW8XHlWDaPiTrhbX03QHEOKA7dKMqHh94cnB2XXXWG7jMRIQBQ9wI
+m+a3YV9nAV+Tbh2/t9zZ59iTWbwYWQtR+HDt+M+6bGPBJbqzyCfvsB+2pzybKzL5moLImiYK4iw
VD1FVB1ans2wgXcYOcnOWnRWZJ4v45Sbe4W19P85fBTnassHbYzeMQ8/CNR2RVCMAsLLJGC7xuuq
mo3XzHvS1mhv3Mog+rxHT/1dqlt2unX3YUkC4aleYjxO0byUgEF1Z8DCTC68KZeQE7X22GeSdar6
T6oCzzWz1MrSvu24ohLMAl/bGYeFpY5qqvra6moVfvXW9MKVvvL21uNDiC4WzP+0S1BXJqijr9D8
FL705yC4EKLnKuuKx2dY7DDO4m9Te8AI5RFlxD1oHMsICLLX/4ICWUzeZdIATvVlFHwSs+OlYwiG
0nkbp8ioTse1IG7+jbiaFRzrhiRLi/8JWvZSc+H14NLCpOmxJXzYryfJryGMLAoTR9mlQuFLIwHl
sted9kzSSLW3EcTxgFD6YVeA5khS+Oc0tLvfBY7O/h//shvl7K7fu/LLel1Bi2QFeE+0jxr+jx4b
3Su+dY3IoVIHFRV2Kkiaz1B1KBg+qrG7bP2zfQv78A7gTdsENVJ5HCR69ZP+BoGp3wizgyS9i0j6
3R6sAhLzRiMfOdoZQg7QAs4fVhtjdv2B3PeacEX7OHhEdn6VdgD3NMAa612ZgAZJjZMUkRGblGKn
2r/qRRd+8tD9JgYa2sBft+X3MfXOzti0NHhAYGsaCPcp2CF2clVZ6/deIbZuZNFk1urhxXDSR1Vg
9VBbSVUzSHdj6+SuWtAwoOd53e+o3EsdqKDwJgMQHELeDcmyLxPqQFJnbU/QWeUu1HBxlGayqUir
FJwJWAB3w3n3Z0Wd8StD02QoQukK7GryFpl9KnoxgoKGMZuBBj/iaJRh/HG1NYjRuy/9b7ZfPaxm
r+7E1aO6x/lKV6cTRiEc5PRd4qYmq98kBuIpFjIgTw/yaEfUe9gKY3O0Zjd597GPKJ/6EsF8WTJ0
IPu4KvgpKAeiIM3YX71pVQbBi58K3BDAjO3UaJFOLE2aSMk8WB8XhRjcROKtbPRZTcBAGELj3uXD
XNsG8gBI5xWUJLXtlNKZxD3ljlUctO39UGnjy2IreNx1eKRI+bFyNyPGBZVrwlI1PI5rCa1i1ejy
UdKkEkvvMsKAY/Sqmf0WbiIuL+695+a35w6DAs8po0i/cdF9OXN6RdP+dge8YBG17RlNH+OTeUrk
mThEPjtC4sybeKziFLJB9KLGvdUMtseCOwaYPiQ5hoLiPnuFeEExSZvloJXqj0hzPjW6xCjzwDKT
EUPB9xugz8RzJ8sJYw81CuNWNHGSZnzI6YfvMUQGLHIWKNYq5d73rEw7rjIKKbRT7WfcfRtFPvxW
BCvjsEx7KuG7zkU2IsTUqaRVSV742lLJf9x9e0rfwCb7jFvjm6mwx7lmKBtM+pDFBmt7ZRr18PWn
ltLYLRfNbRkWH8CXrESXMQerpK8UHZUx03uz7xhc0/F8ewSJTrrlg+BQXrly+7dEjij77kyCGOu7
RongnIATNhF0ZZsyNTyR+0cWAYxNgUcvKKyJ3EhKdB2CAGY9wO1HqVATYHyjK76QYOoaAUTW16Fm
NerzucEBHSNOEBBYacEPMWb3h25ZyyIkqficJ6KqUWhjoMqgnXKb0JhCm6mqWKX0L/JAxeS31rCh
/SOooUhODmqQUXXCNvRcnZrKDD18mYKkMTKS5LqQ2ae2pHgLQIfIjA9EXpUooAB6T9IeDYk3JflS
XVtG8XdqAu8goASEnwYlNULuk+1um36l08HwxluBzezdoq99VyiEmpOs7pdOCFI2dBavs/zW79dM
OA7DVr/B6rEMBYhIh8Vj3dAgj793a/vueL8PrJV3/o19keBfHTjXzcybt8ztZEgLtEGmwv46rncm
AzMMk78LdFbB7LhQoVoE0k12rIDZmwjRYuGnDA0Ake8D77+oV7gFSogbCUhRIatCdhsza7fL/Q42
69PTUKlU0jH1+lup4TYmMUSsZBD5/R6/9oB8/5l7PbxNeSjAd3REhDadXm1XrBkbTu2X3N9N4qsi
FC1uQgxweV0EbwRORhU6qbUM/i/4T1K6820LHXX8xsBHlnyqYvBJeObxImJ89PbWh7aDG7xhuspS
AEm36YyB4NuhW9D8e6mwYy3Usa+enfUc6dTdZWMWPtJI5l5En4y1Ghi9MDijj4UdCQqOACgzxRIi
Wu+bRrbKdQLo5Eo3H2W1m6hiJNn+dR22Ju36TAQQqqRy/RIDj0Fmz8LOQAU89dYYQ5tXiFybjgAA
LjxLhYAhbACxpTDTC8+HLes9NP5U1lo4IZ/Jg2xUPyAUhHHNk5VqKOFnqsBeMD5QyzKkblF/uPZv
MHgxhGszjdHNt1vYu4wVl7qhoCXmX5ayG/67eK9vBFF3Mgp98OtpyOGObXmfZT65CZuvDMa54FKS
eRSbS7aox6WEFxApIVljunRAroXODxuvvn5PqM+Ax6u6rlLDS9rsXJqlialxpIKLqY0tpw3PtOHL
WtFAQGMcOvsZbFA49DXKvHwHUSgqebJcSAiF6qEU+67FyTI8f64NryMNlusyEOB+O2HhFZ421aIw
1MmX+RGp0ap2F4D1PGRtl+Bk0ctnOorBxA/ln9XjyCumXo2/wL9V5/6Lfoe0q/OZ95F0729S+9Dv
oJyW8UDue1hzQDi/f67AX5IHVVOmSl1ATKzVbNsoZGmSDU1Vml+QzggGgjlwIXtKgMt4CwjHf/fJ
cknMyZ0qiA2ZxwP+zZ5t4mWipkXco3hkJ6UVtIAh5ivgG81k6Z9cV/ajimse8Uxhd+YB0ar/kGwu
AyAxZ9rogVVou+3nMyhZXUHN8OrKWt/JCf/edgw+Qk2xAZnCrFXKyUUX7mR4zzJoKfYeYS53uE62
wPYfDe/+c38WTAMO60mfytoen8oVBY6UU+oy5wxEehpZJk1FGL7HhhqcvaTxYMBpaD0wynr4ydqg
w74nE5leOVlAlwJnU1vhSTrphy3yl/pwOO15GvJz8oRivBWMB+CLM6Kw9+gL8JAK91KCgGJdyh62
3d8boY8PvvKaI+CHU1GHbG7VCbJDv8Z/Big6BsUgeucwWHgcCH7t7zLoYDduzI5qCRZjy7LqJeAN
dThGqrwWOaDIS+ygHln6ekaYW4p3idLYkwcZYCW2JzaVyL8z8IwOXfQUeAxWq2w90TkBnUb80mL3
cPc84c5hgNoxeoa22hI151Q3sCjKiiKopIVAHOy1gJnJPw2tFPvu4m4RPSmFA7jYbe7RzZok8eIY
yT6SumPoVnXmysYG9wHgLj54DbXBmSZRDerO7F2TOBaDz+lMybfIgZdc2HsVQrCebfXeUr+bu542
/jhuRG0KAHHP61lmWB1T5Aw5o3HdLtrPUj4a8HJTAA+Ws2/I4JvZ5Cri8MBf4Xp0L+o+GEQ7J49X
wgWqN3wfqXOyOMPudvzZ/7Weio1Y30TDSZqPrVc6OFMvaV2Mx/AJZykLwT51iqtRlIBIC9CN+QxB
bGjDvNlZJnWR5EDHa2wGXC64FttULW8hiApkUgJjyJWmR3chm0F+C64sOl5IcRH17z+MVdB1xd8c
v4JcDy30OxbVAxmdl7l1NzZCYnQkDyw5bmwA1rPbqmCSzFdUgE5CxvO5/+a3yICdY3+nXL38SZk1
BkxqdH9zLuViGWyxulZjDaRKaPEZ0cegmBsh+a9lI2DwkMCHUB4TMNVT/yWO0o5tqi6PG0OMkhfE
Zj/2wEDLbcEhqpKjrrLb7uIYa0yPkevwnjOQV1fewP8Tw4hP2UD0Xukei9xk3Ov3XceryvwUyMRD
VCEUq/ERzoOBWwZCoGyPBxVTZmtF7g8e91GfNRnTXcf2ZUCC8Tt2XIq0WKvNlcYubR4EcJxcUEfr
Al5Q1Lr4bByrEERZ2rkee6bAeCjEGIVNxRBm2hMZbNWqTomkY29DjRN877eXvHi6Md3zBjz/F6T2
pylsfoC8V+k4gM/9/wkPRoLgPKakelkCHTQ54UVRydlgs0d9DtX5i571XobnOd+670HTNec05f90
ELBAxSXgzOnhizFms83CF5U2MtJiJ03v5Ivct5i55T7/AsQ2F5Pm/Q2lM9NIXgYtaDMMtTdtZRZw
xb27N7uLgTpfZzT9HVbnYxIfHb+M+B6G9HJPKQMWxFziAq+iCxOGsRi6E9fsrVINB+VbjgE5ClHH
WLhSyVhb3NAeDycbqbGkkp/cRStB42Cde2ScBc7Y1AQQxAYwkK5QY8KUj8BzULXfu7pfNgm/xCLr
YoLqyQVJC4AhMnG1qkQm/z6agqA2O+YO2FuVLzXyxQv8BK2fXtQRSl8nGLvH+kJIxT7MfeedaXch
M950yhsRlpWtU55bTXEG8hbcDfIOTfx6hUUwgxSp/kYgtmZqvfoZ+uKiEpLUAshlblgW9Lby1AE1
rWroSsuIyi/h64vgKolAyF26IQi1hHu8+yLqRLKjtfhi+GJNcWEQLfdNj4bI/H43TofdZGHdFgiT
ynX5Z/ccH70khXMvrBtDhksPNq9dYpP9qq+eOvAHPCmM/aygRaPyCrKfma2ZyNpHpX0G00puJkEH
q6faFJSGQZYQrFXzFa6m/wcvL8cc+pSgxFX9jqO3FbECI1k8ErDYk8ekIztiAJSwU6ryuM4E9irt
+XLXXbfZvhbZrhmlqh6bVNqSR53heAGpo1SLPHBwnpWrjBf6u/U2yewQM8jXGc6MHR1OKlj4aENH
p4WUUOxLYXqGXyXd/rdpt0U+VPd0q3cvAc83dOW2939/qA4fcynnYV5eUmDjwR06+4CofrxnBJzJ
k9yyeTTaDDIKIhDwlM4K6XbW3rmVAEkAhkmA4pVlZR6B8279vecDKrD7xlCYgMItjCglBvfmJBZq
yYjIZexqTCN+E51SoJ11ltMIAecdgwbaz9DrVVgidy0L7uXFBRGPGA0qc6lZ5WS7v7ZQj6kagWbi
Eg37IXSHYbewFHRJkAlvGZoqqzyT+P3SE0eK0NxKzYxFt8FsqSzpeShk0KCmlrATQDh/QveJCVtJ
StVYmdh+N0MpbLwMF4NBLNQPjxyclbdv9bPP4YSOavbk/xnrwfaeXH5DTjSbZdZCnrych/jKrXAF
3uWqpgSQw04Vz54QyK9xxEHZBrBL5861tcQk6ik/RMOEvvXf5YVpQtbmdfVIpybewCKKMarMPk0F
sUFP8dAKDq+1z8Yk9ODfHyfA/onCh8Qw9s8s+I3EbB4Hpf6dhaAjBkAg7brVLtCLc0FMhuRcPB7h
NeposEBwVelhSjfjxJ6SWx8O3IOVEuG6x9MPe9AKHAdXOQGnJe+XyF2dv493t7LC59XrlWklxnP2
6N25IE1CrfAbZZNXTLhzKXanw0fXV3bC/c/KFm969BhiGqjMv8a9WKBr1g6q8YJBorxbB0goOhYb
lEPJSwpYUsnrOXoo5boxaBstIj/9j7cMpZHHh/PUCXUFUrhdbrfarZlol/ifshoGK0w9oycVC6IW
9mJ+HNi6H1cMTEnU51rzgsb/MoPJ37go0hXE8oien4UOl2izw4Nzszn+WH8p30rtduIxwK8dcC1G
tddY8MzElqVmjsaWrNcC0Z5oVmSbEMiU7PT4yfOBDLcjSnjATC4Ob36DxpqWt1M4MdwfkZxhEz6a
9XMmWoqEfvgRTxcRMWG3EVN9Vk/6UJE8paZJ7IVL6AKw8vhriQV8boI6cWBu6YMkq/mG0lEDiwBg
xF/wjMD78O0K/4UO7Kgj7+UJPUfZru8kgKS0fBdhtnlTqGuNC/cyAIQu8XGIn+OC5uk4LizXSP35
JKOaEfASMBT7u18UdFpRH0Ze6gB6tgm7S1SAg+b+FjQf1b6pDiisfVrs6I1hozbGeljXEd1GcsVj
bLqq7BL4FiJ3aP4scfQjYUSa2jmQLqHjWBbePr38OohSxcNHXrLbFM8a0w/OISTeIRDNudiypgtG
P6DMRL3+sdLjDIwfvnvr2dEStAT5KvZ69aEmLIt9zgJrLrKPXgISl0k4rNT/cpMk+tvFK2sAv+nT
sHCh0Ir0hxXJtbztT+8rNgYCw3wHNMRP8GZ7DEqJDGu/CUc3fTabxElXAsFZvWGXo67hXO1Pv7eM
fEUGPwai1A2TnKyYE2EjuKVg9L958g7nbxUVdLQ6Ro8Konh1953CsmWrA3624bI6qGXzcwkytFFv
3r/lBOLa5vPDc9rK0TiOq938Lk3SxjjfFGury+rJfs7ucwcUOSwvUE3ACPD2uO857cu3CmznArn/
5OeKAoIJOMK2hUVI3g/HgJGD955UegCu3Ob81Fq/QL4V5XumEeZn6kjGzAuObsMAbucwHe0rbiNK
Ov55XuCeWdZ0MDnWkkNbz1TZFEhT+H27QpGv11WpEQnMTWWIvHexkZ5E7IsuqFwM+ics8HCd7cNF
QktmLxsjihXu2prg/ruJzu60VnUgRuc9G6sQlZ2QrpXjjtDIdeTVYrqYeB2GIwY++HbultgE3WvP
2gkKE+UImpkQBI3M6A+oOar+A2MFNNsF8RUeea+KNsk0hy1iVMDJVazxEZqK83IIa7YJ+uN8gL+P
y3zw75rHxYNNQEugH9ojxBcBQ/lqRq4Co2phUxw9K/jvNTdupIDJNuUh6QsgEo1AlbCHUR4sE1id
GtEIwqrJJ9Q//8/4T9cHjdaOGu7GzXsX6y5hXAMKh6gYs3H45enbdGWSWO2zEOwNKt4ZrLJATU+0
SPmUJ9zFEAEiLwVSeNjPND7CFSYFegXKJVJDEx6RrbyPQTDxKYjy8zGY2fBjTbEUKiTpHA/QRG7b
uYUqYfxru4JTMP/XKWNATEHqoQbaA1pfxugxmgnWuCLTxwkX4raHxOCpewc5fQ/luRgMM/aj3eZo
21wpQlURsN2OEVubUrcu8ju/6TGsfpTUaUVXAPEBCVfjqP+s5WAW8GPvStZaLZk1j8CjFzReX0nB
vFjPxUU1SQqJXVOyiN98GK5WbWrOxqmuvahXox0yaJSGIhA3w5owZqe4QVPXY3MQiq4zIrHP4Nrf
nG4JVba9K8L6pvQyHT7Um+Zpvmq24P2EzKITs8EsiyE8HL1lMc4L9le90TgO/lg2LtrqZKCA352Z
fIx1m+zi2yuDRyPfRyucOw+LDL8CMYjasE7CrrrVu3rpJ6VXbCGsAQFlY92x1vZBxcWrIFLsOCjJ
AFGo1TBusVOtUb44J76LkWNgGfUI17O1cNl8EEb3MCn+ubSG2hhbb3yoM68GdlCHWo+ELktdAXnW
BquKccW1OZFwefkeokNcqwCKMqlYthCBhA6dcu5DspAOGjl8iiXRDdi5XnGnTtrzAzOpbrUz2aYI
E9BlBr4xi7ayFynsAxTkwAUA475RLD91W/aWeV+PLelEsIIGv5dCeaDC+bcEBpOUMz8SgPuHrsKY
chqwZC29xvnn21A9FlsHWxjgiOwdBFo2BXXRDyXST/RNMmkHsFBq8oaC4SwZOQiSEf9XSaCH23/u
YME6XfKoOtn7cChJ+TPs3llaLrgpqosAtv1LNm7nLnkTHq+7MRmCrbqA6W7Kl7C5M34F/V0nO1To
EJvDjTTde9dRiaIoKIc9x+gcBcYUiMdap+3IxHwi9bYnuHvAu1RTW1I/dVcXTm5KQX9fwZWfnUPh
Wx52/WJX8IZUHsUQ1pHU5SgTVWDtdkULjg5L9GjcLZk+SHbDqRBPOu+RimckCRoR+j80QsMBq1kY
fgT6RmmZG9XmUqamGAXQZSoJzj3eakxYSCo2Tc1WptY/qmOJS6GRkLl2lyvNr5Z92lKZLsMx7joO
0cw0Qb7XFc5v7SgZtruOTs6NyAineKB9SqHDDLqUadpdm3pJK2gRR1ALJ4nAOrd1RblYp+6Ra7hq
FHgAONWUwcBuRvRSWZ7lgGU06HVPzA7dW8qio6rOZsiPBP+j3yEhubIKbQpVM8CZwmGIM3Kd4XA6
gpqBZ+InfdlRGqAXy0QKRjS+zS65QRgrfMwxrYWbaV7rvnUVm2Fbpb53Ek/ogKCTK9uxAkABGh35
RlIeGq3iJhdDIK9cadyt8hfOIC3/mH4uQx/VMMqP+1gf4Ik64tkDQQcOcrFmn6nu+bk8bO2z+3dw
3IvIbhkhtf16p4CJrrZuUOaDW+V5HkQVQdJ/tOFwZcSV1IUTFAPpnv3iwKzqHqIYMsLkEfhmBLkf
7c2Xqnv32bD7meaY8tkiOW6ojK6W2IAFMwRntsVfaBsxol6QnHeILC5KbtlsFmGPsZsh56goV7yf
r9da37Q+tulKToigtMkucO9fFL8ZjCYuW+Q0KNSfiu7UClWAGlsKg8Kk8Qw4rVKopHu9zwn0p0OR
jbw2+p6HfLaImDiJ3W6Eiof84RWupJnpPIJy6ShHDIFyFCbmkfosChaqsbGfJDoeKoSOJ0Xabzly
pOOQ7HO2MHANmeUUmhNNMwsk0mR1B6cxLTmXJReYISVI8fLN287z7FmQDNe5k3bigyKdAJGke4eH
Ihe+YJ+TUrj8mlTLudQjMnEEqRQKbwWq9+U1o1owzZ4j5l80yGoX2UC4MN/FPi+Qr8m6JmL5hZvH
/sZILNiang1bpoPexP7Zkv/DLhLOkBO4sngpWNjRw0PzG9gSbcXy04KrLa2XRoToxDo+3l8tZLUI
jFXDK8F97DVLhy2ot9oiE8lXJL8wT+SR/xhTECJ4g6wNkpjcM9SCssFXUUTXYlYGDV4LeJBo+l2n
kAlzzR84ECMXA6daGC8co4cLq5G3QZz7WOx1sDXjY0AR54m0FIC0NCQi7LaoYeBDxM2nyzNCLJiO
DQmQfpMwt8IPgtlYL5qrm9Y8nCQVD8TDw+u1IoqO0UHsz/iKcUR2nqQd93SSmGmlLO3YELRbf9I0
+68XcezkmUqDmGzktQxrzsSLpWkD8eB3vZSD8g7xX9mmKvoIzYxx9lTQDDdIKG9/cAYOjq3kO0S1
Utr9khDQizaZS8EZFWAFvY+Zx+Rf1pa8ZIicEa2Dlb8ktH7U7AKZmLy6E/dGCg8Bi16C83u7Npaz
ALqjTl15c8QYwwigjQDAxqSdrzcKCh0oz6N5kgpYsP+arGzUPNvou59+AL5knYrNZ6n7OWeAVYKD
+A2+xA5TFpd49WedS6oID7TV9qVJfVtDgmxDANoFwvE+88TWHTjuuRUgOsLhfnTBPaO5mKSg/Gxs
RBG/NjkXEMfavT1uUyAfosmgca3nkGQuBgq6NjhS1cKuHtzGg9WPKyekm0lYTaNzb+aaZ9h4M8BC
gf3RwP5yuw7vKTuFrlCNNrm/f1Wl+eZcOxWPdIKFU1Y6KF/OzHU2BOAZp94zV866TW5iwoEw/xY0
RHZ/ajDC8CXsTrakh0KF0sklrX+q2mKKrkVtohUN+5oJy5jVT+Xbwqw5vBbNxP0oyfg2U7U6etIh
G8YyUb0elyDxWPmFf2GUkv6JsNgPqezzg5Gd1t3tfqb8DD/TvERf5IqfeIs+r4Rw6ZTe5PgBAWdN
EAFfMZCJWVfEljcEzXcNv8UM6iHLxgfjYfFeZ1St2LlHdClY4jP37JBw8eJS+3uYaUItkMfcnrPz
ViTqBi+zy7aMka6/FMZ1nmsdyv3T7iuxx2hscwbvxmtG0Uo4RWiaoqyzffcstG17YLbvVQMPgwjt
XwPnF3z+8jPLWS9FjM4IKmPGbIUUiZJ0aGASFIHAhV6zhk6F4f5mTDQGUkPXKPCxQa5UE4fq98y7
D0HlAstARKFj0a4DuBbpXQeh7xh6AkZUtAWCjgX6gfLTNt1aNpWSlgQRbfgJ5ylGwkyBO7FDLFhu
3kc9L/cUDNmOz2BRdYTZ1t9r2eDQ1O1jXHHQpI62UbOTzyCy3CxX33H532HwbxRAIZ9nL3XHSX8Y
V5SKtr+5L3n9TkYvQuPL4WIb6fYzp4nb9FzMQfEerxvQXPLYakqU6L79EcQ++zvSwFsM2AY8T7uu
KO6d2hpvNPPmd5oMDDEdS9wAAgWJNvn/U5Ah0HLeJVJ8adTWM8a8GCQYQkb7+ndjC9aKupnPw38n
53UITJeitar76qCyCTnPzNQ+02wWTM+KHSewW37H2URtu7+nld3gkVPCXXjDBfw60U1fjn8bYCtf
vsbo4A21ryTu4HgcVOc/PLBTOo9GlzeuFnQg9dmdiaGlvCc3fLx/sSeUbbdLB1wWIpiD1iGHri1O
Ba5hMcsb2tSX+n+iJJYMWHlowKtIDT1vqQyd8vn+yyJgG57c/2S+t9lCFbphHmrsOsQTqDTj2SFC
sJaRxW6Y6QrSIKD8zq/m1/oKa6bsP8NK+QfCWjs5ULVintC9dhnYwyVzwd0y0hRWFiOUdpP/Luki
P13FFsMG45VBrcesKlWOFlr93Czl6bEhHYvaLYEXJTDRsjDNwHe3sS974W3fbepZuyh63M7+sjH2
JuE6dy4rdSY0abcMy2VfaUpQO+UNRpdu51orouQNaZ+wKadxTaNzqwQKLR2xP1CGcKAtr9r4jwiy
qoo+u6XTiwPTO0imCpHnx9ppPdisRcFN2DiHFGCFhQnQ7bwDYVCzV9WogelpKXDg/VtI/GJuuUUE
YbDtMWThCEtGDkOKOwFz7A1lcblge9x5cZvdSOSyeadAQCvBFsEy7281uBAiUvK2E2VOsrhuRhWH
sELeGV1idN18gSwzoL+Sm+eb4xuHAW0FyrKhfenQ8MT6tGhk9zVEYCbzSVFF/ieXgA93M8+jZVOy
jZkafRREt+hg3ApSCePsVOtdBtlv6po4uaZhVuDY6/LbHdk0FY4KyVMBjTjnV0UEkYdF7WHIJsNA
IN0IiyENNY7yf47OQTCH6+egaJpibKJrHmGhWhtEn/LOKnzWr6MB8GRtkFr18LLerNcpVdkvahr6
Bt7hT0b42OaNYV0FBQAo1qfKwKyz5m9lktPTjhUmhMtu3w4d0MpMytNpL2lbmz3raGImUUPt4V7G
/ZGqMZ0yawJ9epO9hVOZ+zasOgsOvUzLNjLDgevDcYieVDMG2av8gI7FSmV8dPUjHhFOtwjvedWr
HVgI7AayDt/k414eaL1yrA52z3srmlO6JqniKL7Dm3KXyNzbpUUGP+Kzuk18XQdUoJ5XYosylvyk
c/RbcrFm2VUaDGXhuHsCCE7kjaIYY+pB1bX1u5RV/F0p3MaOZiGixmetHwSZmGRvAiSGNkQnaTWb
EzGWkX2p5HUyp0NiqhoqSzBUhReB4antU20PovqeaTd8ubECc9dOka/Q2Ivv/dqpFqRJ9iRGPqVb
00KZdm6W49KZRgGgQdQ9B91tk+ZF3dWpYAQh1Avn0lfR2tOiUCUykoMRDz5dii8a2LUgUqw66Eu0
y4vr4sP1mSJPfVrnrsI2gNBDgdlbS+5aVfYEMAUh18CxRJFZyD9QqtN9n51g5NSUSWHtTZJHQiOc
T2kI0QNMemkTaoq4SZvq8yfBMAumih2U1L5qWtDf9TRqFvLHAT+2tfvn1t9KdLQmf27A5DCNQ/fN
LFzWPehmsGid0ggq71edAPgtw6SxYKpnM/AD2/yl3VHdILItwGzIXhiK8i+4xocss0tLC3HdeaJp
soTqQeU+TnmRb/0J1dgCV7FAbLWm7n//iP6fnGngXoZF8bG7CoJb09uR/f6myU1Xy3J4C6IyKAxn
6i1JEO8In+SqmgqC5HVBCAbFE5t1kk4ycTZJd2nl9Y5Ynp6DofXXnttQPj7187c+MKs9HfSfr3Fy
RyPqpTLCoipA6dkcZLMXUwnUPmJ+4ICCcmupvFW+tYQxNyeSgI/yBUPeEKRrwzEPoucWUPiQtIym
aGTudRG6OvoSeNnXgMSe2046Gu1BX74bOHjlhmJYP8sBCJmv6nfeZgNATxHReRoFIQ21wt9d7890
Lntdw0rt4VUyagH1+KdnwqMGEzW33KthcrrBwT7SvNH18P60Y4DFurfZfj8qNcY85Ogeoq+2U1JU
zSxpoTX4ZTwi7WrJoXaTN6ucwCHvFggMSVPA40tfBLMllwXQiO/QKoN9cfl4ofPUcZrJMLrzmYeA
+2o+tGjDi8KVhZ+c0VIfSP7PRoCPe6p4kXDkvHshcGL1NVU5kXS46nJXKgKjOVvaOGCIQO10v9jB
qSCFbiTlESGw59+jYer8y9PdDbqQbLVxzruVfmsZb+fq9AoK+UfSK4vftjOZvABWZzWsAC8ppknQ
jO7KpfAgvaDkTtVOiz8q45/sWO0W6pjuSBMXULK4rTcpcRRFtEAIyOBRvz/S1J0qzBgokHHre1WE
X01P95eNmL1UclAW20b695Mz0iDxXu0KUHv3eXhNFGNMRrJvxclfg2FE1t5oKmccp78IoSi6sFe6
LdR/MEnzDBZUHI/p85yn3WQKJ1H49O+izepls0q92GvEZzsWh0baybtDFbEteY0eNuyyEc162ozS
7/gUD7zh/naaUxdqrOHR5YQ+cZA2LucYrVSHumnFzwQ3D83+PHXrFavMRwF7fqM06sL5iI0Xh461
/A2s2RZXzaXYZvnyxDTRferMs/j/pH4EvZb9tVFIIynlRW4dwKkc44qE4hnE6GywEjjWQ6EeLTt4
2HcPhVZIR1sw21b3OV9pXiisVunsidfKwjs0oSmzstgs1wL99ZwGQbsZ4UK+tQqfsfPYhHa8j+E0
jMmQyWSGHa9sShXKiYcm2d4F1CtCVXuMx0mBPbqxFaVL89t5pCcjLNQojG5k//nX1UXZwkwtL6gT
WAHeR0AEUTuFwPTU7ipIoSezN58n36/zjnWP5jDIBNEjj6uTa4WQbiMA9IRd5YfcWckd2GzEDEog
3h3KQUc3gEcUi4CUvLjOLEb/Yk9hwPL9plS0zd3ZLsurwSVYJjlglE2tGo4YUDdgYZCeZbuhOM4c
U98G+HfIvhtCrRYJzDss7ZZ7cS3igbtlUbX9KHqRpRr3Uv5YT3/MUFkF/PEYDx5sPURrM6wTEVuQ
8n97ZCbOBbMg7i5e0P8jxppnnlNeLsw4oDZUF9wAvH4zsNDttFp9LEI4kafcEqMZdNUuRHHunpkm
LSaQyAZSCUB0DhGUdSR0hUversWbmd4+RYYzSmQHjPqJ2FDqnjerQQ77BhY78qk/HHNb5Bn2BE5Y
nPmaJYPi4gIK9oJawiaI2W0IBY+Gsou+OXD1aqSZr00/REgFX1cVxif9FybfaVagwjtygP0HfiQN
KtrBWS8NicftVdcfjLFTgApVUF1IeqzxlfslAx9mC2c51hQn+Uek3CtJsbXphhmWGIbDx2meMxdk
h2suAvo31r28dQdntIOCISLxWr2jXBLezAjb0WAXP9RK+8De0tBIKQLHf0Kssd28P8CSB7APDos5
SFywi2EUNipzyQEjoReGG5bI4fhgU8Kc3QE9F39n+YXz+HgFqHez8xy0dOH2rxEHL1c1Sl17v/mG
YKjeiewbKKcnDJhPsi6JN9orqOr122snTJpMH7nx9AgVOAivu0Ub/Fkk+0IGYms0Y77TC9llvfdQ
EqjR+/Eki6VE+8gkCTscZHSoCIeuOwolG8ek8+XL44o3trrCPAMolNAKzl/yZ3w6zjDtOArshtek
hUVNzFDtq/AK9y+D7ow21+uVNj394C3CEfvevgPSO0vN/39fsVv06LcNf+tTo6moHzm/JgwziLjF
L65Ap2wUSnB0Hxujte7RL5EFRAFiCqy/5Z+1oPAOVUJglcDt7z13DVf13SjyA7u5QZdaH08YnIuG
rVyoLUJnGuBb/4gJdqkMse/poQzm7iyPJbHGyhLPR3QFkMdmNm7UodMSdQVq+otsGuS6Rt30cSRA
dgiousbt6knt1CwQ5BCH12ryMa3cr/INe3+a48Cl+2Y2LLlwTFJXQI/bNKLtnAdR0V1R9p+V/mMK
/FofQlqYPzGdEyO9RfRlyuveNc8Dl6k/KdQcavUbOyMG/D+Xrsv89Xzpk9sHZ+47Bg3uQnIY/mup
4vu7VwiC/yyWvL+32EVa7NJQ92c2jeuHiiI62f3/WE3Avdvd6MgGbjH0J9MwyN3n5O2ODv8ojeQg
ZtOWFCu7Tx635ivbnPPhNqQkSzOb7oV8LEwQXDNqSqIYSxvS9nEhyOI0tsUG7lD3X8oFriYfmvvP
pzY0kbG9SWyT/J8H78oJkzAMfLse9ST893ce1AZBUV1+CcdDq2JUIz8FxrlKqRFxfArulsQiMPfZ
5P5d8TZBXsPOI374k0T8KTOOEIr0pYO/pRZQjjcOa6DL7BChrvBzOGUK4t88Cmk2XZWf2Nk2/TvE
OReUpoScGidmxQavCu5tqPEzPUlaOM9HyC1HX7XIPadjDWTQ0+rGk8HKlw3EzuuSIWcuVL95KeJ+
7U2th0AkvWIsgab0EsvaVWEMSg5EEz+z6XjkBx4O1nI9JK20lUdQ0AI41q2XWrpM7jd9StCRtWHl
2kP3n4jy+urBNdrBBWWYejprvMpwXmQF6QkPc4lmB+5/9ZmiM+p9OQirFkZG3M0YFqAsJVbtPeyb
bkGwLXZhHhQMGu2YDk8Mn4nsnbOnbiifOSGBveEpy5kHh9O/081KFrt+XSWTUiH+pUJvmqL3zndT
b34VZ5OeEg2rVgKRRi24ELE1ZSO5qUd4dikTkrbjds5I9aebxHaBZbYfE0hgw+I/+aK9SD/C/LEX
gtqogTfp3ynSfLW5tR2tr0YGuxNUyFV3FGizP0m4MBDhHkcTfT9UJLUp0G9g8ZTuVY0YB3Z9jvDV
O/gEPGu+HlK5+vVm0sPaRKtIrHKa5qYBn0/7dYDbLNcsOgZl5uiVkhZzo7ZRhBcExJTmmntg0pKt
/m0t27lmG0sl9PhiFAr7ZRQ0IAbMaMgi50Ht5NA1VfUs9gDYTtfDis6PsQMXxWv5Odm01dsNhMvb
AKDlZPCyUqAoecqlff5s14DmIzLLdAjj85ei/QdWQjMaOlFIrUkKI7HOubTQWGt1IH+HXSpXEPt9
REqhCvdgy8UDbn/C8towkkXzRhxkEjhh7pRbAZ+lGSeLYe2FaR8NL9LOYlWg4zCgHXJobAjOn5Ex
DPlGT0G5AGt7wEIz7VzB9vdsp3Qp6d+IH9iCUz1p0bPh9T52/MM6VALE2tTI3iyKnvdks/6pIfZv
rUaJfzK8M9mlKBPtdVvW/JkM5baUzs0l35Ke8o9xwc/zkDjDVXIMUEtDCjYF2B9juxkddYog/VuS
G6X/kuH3w8MqVBI1+DCDcbDkwa8ahrLKTu2jWo+xULaHAzYGPpENkcTbRwuydjSacIDeAVjL36NA
TRIQNtAO6A5Kw14GujB2Ni++pzTGRtsmpqRQjZT2bWAie9VT3+FjagQmhmAdsbp4UiGBkUDQDDtl
3pw65PH8WF7dYhbG/I3khoWwtuxnR5dgtkdmsM60Yk1OH2uNZMkeCQOPkjH4Js+vOldB2t6qvc4t
bxeBq97l/bOHPW3qpvufUk5PMSJggtgmtbjXaQ806wyD5k17vBHLQBcPnjTmNUn9yeddzHttLD9b
qisf/8Geg/3o+dp5QPKi1KyAna6UOu5vwqE0vVOjSCel8yy/xzvG2S7iaHSPZg0y/MkSTac0K/nx
+bT3yjrzz9xYwzpveMc/hCUJ6fGqEsU1n5Wr2ckbZ7FBGRXkJiO7XtXuDYTs0yqcjJiDh4odVEcq
z3nLLXx6Xd4uRcJuGq2HQbaclrfbj+7VFUI9ddcHNiqStGe+H1kEni9V5jXr4oLGqsJb6PPwlBBG
YZMtKNClKNpZNwesAlWI4iyfx6Yh45AtsEuI0OAxs7P9xYq95D+RnqV5M+nZoiB9lhK4OH8LhtRD
FhjBA1CbDNEu0vjMQzl7JttkoEU97P4tKzYlD/5gnkq65Y/kkQC0l5/SsFnltj5C/CIAqZa0kEu1
2g/cbHnYn8+UgrTmJ0Ry0xdH7kzEJz39I0Eiv12Pu/J12IVRymNAB2P+0TstA9GhMBmQUBmw+Yk+
Tg+FGn1yWLDWSju8wfI1000ufduycLMhWIx+svzD0UGFa+gXT9rDhkJG/Hglo33ztTzzU7TCHdVT
sDl1kq1PRuozwV5ecpqEbygInHtr3MgM9sn4INV2/9bXF5TmYhWuDI9k4VIGF2w6vWjQV8954j5V
3+hAJDk7Ykunf1bzAZ1nwUKS5gla8ROqXEbV/AEFDhLmN8Ohu+PMswtMQUiVZsP0B48LG0LttFLB
hPm6Jsh7SlTLJQp1sMYPowIxtf/FKFQQOR+eadNtDJ0GAUBbYTvNXZmIziAtCnM8R/myLFN6W//m
5+CE7QTdNrU4buiQBe2f4hR+v45icH6joBt3zNVWWGE6p8Sz8aNfCNVSVfS7ddQnM85bNPKA7D4m
BqhtwtYy5909xMLFDIC/2JXwHpAGuXTbPbdCpjVvSpIBUgNGLSelDKv7ce/VHjunEcfIYrTRei3w
gpYM4FejHjld7Q6kaR67XOmvy+gIW81TpJzKxAlUHNYdgIihtw9kvoUGfkgpTZrCkFVVz4D5uFY8
/6UFekEyC3Auq9Qa5xTGwZrgVD95hRjPeze92pwtokWGXq8by9N/IgmGaJrcnEK1+BhvOZjS1NRo
g/jS5QntxaFpWLo0CW6hnuLUnEk289d/VjCM1wSzD/dAkwh9RpWy9fqbJ/TbhWRZ23dnJMUOCdFc
nDsNKu+HGVibnU7O94eh3DByFQFdYP/jLlSazS7Pmofxi8NI0x+tdGfqQF4J2SAq/0bXa1jBqjVW
WHzxQluLquJ8BVUYf9EKesm2mcUdG+6vvVZncVakFqJyPys3faRWV5yN9TzbBiZSEBz2X2LD8XSn
La8EW1AYchE425XmdAqd1GV1LH3xIOnZLNqns/8URDtAr1P1MPWiWev6FqyHrgGqnvk4GqKIzJGM
6K6QGz6+Hq9U7jw52DUv9ICJnmagnOPLI32Ws1zMiM+/P0yIWnQ0PxwmhF+k2OxBoNuN0HDx5B//
CVxeCA8kdgAmdT3Uz7VAgraVEe1hNZsOglEcAmnFOt2KzhNscUVEmMmBupLO0yN2mGMo3EJFyxnm
lyI3Gb871XUiJM/HHZYGocsWdUBeA2l16NpNLQZPTIXsTjY6//QtFZqYu6sj0KD1oA6lV9JJGqqg
O/d0hGRrS0mQiqR8QF2ICfmGPhzg7j0BkYoNfIbUnTGVPrML6+UieOD5Q0IU5lPuJXh4vZYUOx9x
W7l4FAq1/9awYwrXsYJ66Y34U06881Iv1GlaCnjsbrp3lsmXCrRoxlQak7JOBapJ+Gl4otTdHHTV
LXOc4rA42ZPj/WnYaZnK1TgyAKcEuwHB9sfAuUvAj6a91kLmdjrP9YFZEoDvgej9PJOnyIofJzoS
A1au62LD0jk95X4ZzJJyGWnzplz/RIC7W+zhcABhA6M59vTVIuY9YLMRNHaQ3HdZFZ8vaLdRwQjY
gDOsJshOPRAToj0yc6UtKyiWFuvNHroKOnBSJm5JbjcnBq0F/icGjvtupds0GvHjM3soKWxqaLqw
4huzGJ8ZPYPDCMoiAWMR6iadkKz5OUWzexA+v3MA5lEH/a5tSTDcAk0cBuaRfbDC7URd48KFgCFR
Q3vgazR6ldrczR6bld+D0zBiKr0JA5dh+iFpT5wvD1DZaGhuIWBY64tPSAHZnI+r77m6w7kkHiT5
grdCIFlL9aC2PsMzuq8wxu4SjT4YL1+QcpNiNKsicu9b/sEE9wpwrx5FM1I9fLLytkh0NN4pYsNm
eCnpgs6X2cME5/xWaOG07RlG6aBc3NNhq6l3u4e214apRbfyn022buGyocfB9TbbROrmZ7JWh132
xGS19Pe2iP+L7iCpQNpUwtnxXrr1b2B3HIuhulccoM5lEcCbUVf4MtmTvFD/4bg0GFAPsdevn5Fo
jcYAb4FH7YGJJ0mRFF9bcDHX2McvKNTx1jz8JRZtS2UpfWhJVaxhJC10ysS1RvSowPE/FdYLJ2IB
3JJp+9wrmQYorNtWro15b+9SPvCu8sqaaZgOeiC215LqcQbO7JE6/ldw3IIeMeWeFPfBXmp3D/35
PwufeP8pTuluHRvplDNIspqV234AsMPv61ZXpdZsKtr3QqMM5cPQxKxtQPOfoogM9wCMj+xdIz8r
lc4Cgdl5N7CkIkKYMVX7FpulJhnijU6/ZPfCQ8WCl4WpLNVR/gVO/D0vX0kcHZLLp5qECpR9kCxh
6sMXXF54Ub7vuE0E+UNyqU3dMWVHy4OBDC+S5QNosREVbPrxAfHu6NUjmaQmS9BAoKBEe48jdnnY
UlwhMchJs9gEF0FT+EOjselfqcWyvNWfjHTcEHNHjaerIYH/7Y8DBl4lwxq1/1Rc9sXywSLo+GCc
4W+coTQRA1QlKPlOlNHZxSRFWUiGthRe+39CVJI/vO2Ls967Gkfj0qVyXccZa+RocxqEo+H6668q
aYwy2ag+fHRA0YDPifu0oReT/inwnyfVHQUOPW5cS/fkbuKIsyB5uXadgiLPEBtn31KkY5O3bU/h
li6OqN1hGQjf34MisoS3PEXvW+8cIfSFlWRYTvbJq76tcas7jC9ODKNBGqEpFPqhCHrKskgY/5m2
EHd1DaXgV4pG9lD6gBTogDBXAaKFFmD1VBBPp0OwOEwuCUk9JO0KIL0wA+Fb5aYG9EhTe7rGzwoF
CNL99y5z5C+2hfkcvc8n0mThu+hGHTJSobAeWrgovjAFo10cfCJ994wMvL6xw4U6d8hWNn5ltte6
EYJ8l39EIkpLZzd59dLkGY0f2n8Trbs8OzthxJlGZbeL6XkxYbNBSkq48tgfzYoiyIGXxxbItYqE
p25XMVvj4fr00dcFvaS5SeTcg09REult8T1mze0yQY3/EY5RKnE/bcV/QlpYK7iVSjyqyidwEmIR
zB1nwYsyz1nu09VhofgEBWUkWR7Cd8KM5ilDt4gGq3dnaqI0xgxq6t7VqmikFgCN90aKDwAXpX5h
t8GlXZCk75q2zujN/KeipOpDz4j1fdiCWFxjxq3LazHtK/FUL7Diofir2Tv61iFT3rOqFBwazAE1
hM1x4r51aLYY7Kd9o+Np6xgvgAQueP1sAQAxK9h92K2HEt/ZPWomdWw5Ds7b2JhyYMH3HOBvl8HS
/rRbyGOLIWVFNa6BrxigH+hyKwtxtOJhK5MJwIlApPx1+g3RTUX72DnH+pg+7HfdHCVkacusPmQE
7cGUWBDfzHyc9PUR0ExC2fSUKNL9DCBKSJie4qiqWxTOfXZ5Wgio4zxJGXrC1cN2DQBzWLcE2WuE
0VBMN4fNvDGcxYZEBWUqnYe59dt67HAtl52wERk1Brre+ElFsbl9XoG6clQbrRbdsssiCimpsfPL
ip0NzTzcZStC8fN2f+pblr9CaKxyVqfiHFar78wZ/oJ3/yGmDWqsc8QJAohHkb6vem07irwjL75M
UllJ0eMh0qWJTexAhQzgcGHhvj69FvB9ibE8nlcNH7JsARPFjo7Gvvq51mx9R0TxCGGi0ECdVnIr
TeRMKRsTudI5B+5Wv+OOTK+75MBvySyVE0Dobg64Sp9ocuVTSgporf2VxtgrnnEQEgjgF8KWHugO
04P3YerIM0tK5n9do+84r0BfmHTbCUeJudHzhwDP53FiXOqRR/1+0Lg09/qQ88d2CypyqR59yeJV
wbdcXRCWMWNpy3ZtvBRVXq3Ysggi7rjN+9iwFKCdMHZYR+/oISjUHbykrJ1/NQU33/TCwBcft73O
btqmHNPs874gL1lnt1zsP0ce4D51qFjHBeh8lN0rKs0C1pVRZvDuacgqRbbKYx8SYhof8R9vCZpV
s/Fz8AWAvMWUlC9QM+M1SCAVZWvESxWu6W8NfEBh4+UguF0Y66MrIT8oNrGnFn6CiCj/LDyoh9Oe
q/uuv5Dr3NKXFVwY2Vvw7ccmvaUR43BG4uq1xfSAmZLXXqRILiBHw7m+vVDYzFoAHbvHmozCXsRt
v+xnVYxe0eC/Jv+8NAUe9fJeu+unQY+BMRpDMGxhUn29IKBTBzpJAWlzHuUHbyzPWu89r7fdvgQG
9wCZs1ecw/Y0Hnj5R2yDFU9ylKZEaU30RLEkKolpuTg+OdjFTrfb4hFrKII8cnmS23jziGfcQtS3
UvqGnT7NPQugYLjJffVKmoa4M7imu291bGlpwwvh+RCpnQGvmvfImaGs2hj6ykJSbU1P6NB1TDA0
/ss3blh6VmebBaV/2CrpZZgt5uY3xlBN7DY2U5mVexIQzMsIkxKycQpD/N67On5PZoqhxkfaoqqX
JFFLFxn0WzGk7QtZno26kTBXAY/Ny+3vmamimGz/Kqfl2ZPpSJ76iFMO8Blr4Typy74QkM9ifFJ7
/L/qmQjrEV/lEzFb/2JiIhmq38ja1UdltACwZyoWv9YfizM56+sKE4i/tlqcK5x0jKwCj2G9Uz6m
WPvTIfo1MzvtK858WRk3a0klYp1pIKFoH+tZGaE+a6jBQbaI3SXbj+F6eE2TmByzcrlSshkPrbz9
0VPF6u5t2wAsMOWuuVyVwQy5cKDN9EXNQflU1QdNWCAK2MVtsITXejUFgwJd1g9wCQ3qjz8S535S
MScl2B9oCe+TbLGAbTJg5863l3Wq8RcSkn7/qbD4TfUW7wkJmUJamWSxkEB8JZyr1yFPv9398b33
twv7r+i1FxdBHXDff7r2JAVfx98NKJRbpjTG9+ELccB67eaOmdcUZkRZEL4zLcUX1gkzT9rQXlWF
Q37OaGWFXtexITxtXV203oaiLJiAAdgcGdtBil6kCL9pqGj5e1dn0MGwQ15s96OhT/ciWdXQCvpC
aUFVWP31aCC5ZOJd90t4lAvW8Recz4VbgnRe4RyhyrDepv5ktY7cj9HYaFTOjqxqk5r7ttAuhV7u
s/RvzyTAFy0VDDtDVs1gRyyC7igsoLa2v9JPD63kL+KJLmbRZ0h7bQ0z3E9ISFlXazdcRjRTkyTu
JF6p0EGeagOE8ctFFqxtXpfvfM/zQNyxu4snRs5gKDxCCDaJtUY9c7EqFaCsrkps8L42t5nbIapb
CqeR6PFueIjioAArNZozHcqZnQ+N8eqBfZ4z7/WyCSfsaYERU5lexCcGwSS9NqXiWxso5zdCrB1b
h65JX/Vcl/bmtI2ziwjlMVZlOXWX9/omNicf/BVLHKtNrEBOZ6BuQoK57h8lmKvx6N3dPmFcQCFG
fAdrBclr2N82WlVFrzBtCuZSnPvcI+wGvKnrJNSMgzhR8LDJVtVSI1oKFdn94bk4t5YsVe5q7BhB
BuvyxeG6mdx+GHgPr1B0gJ92/fT2AOE/y6ddwKfl6pvaG98jPafCTbxxLLW54qyiXX2npdDm8rs5
qYYKbVl+ipZnPCXeIsdXfKV3juoI7jMnCsKuTSceTfDlZidAkHfxo1I8g8A1jDSx5s+6FbHwud2E
8iF5rxhRmgrpdPMff2lijSzzFJ7XaaUj0bY1L8oyH7mIg5hm7UtQpo022BBK1tXe7I7p27hT7gY/
nai+d10FF3IcyAtPkByrBvuAIhJuXDqii51Mhz8PnV3Q2IbjtykRB7uP6ELoSMdQCXkYT1QZQR2U
UF2kVdfQUJS4eRDmXqgQEMpba/ky93JBZIdq+ayoDTTb4JibV9+pXdj4zNin+L9CuiD0tl0j7fLM
kXhWtcRC+jh0mz+aioOnn5oE0IF2IhJMXHi0qEqymp2Orz8lcfduLdSuaPr8VyjpzWFM6u8iF97w
LfXynD7o3IDviVjg8k88AyYvneJt/TFscH3coRtoIOlDQh+GWDCLIdirXJOF0nTUaS1F9yrV/Rja
braDFPAX4WFcA143RUDe8MxBdz+kX95E5p7wRFWgyNi46XMwf/PkVCJTl+kPWXr3poDyMcrzJfzQ
112nqJ0gaTjoui62PdDodTzVJMrd3djm1O+zvUEC0LylVy1PxHz7F1FXWF178XHeYkj4UeAGXZ6j
/LW6tI31GeMYRNCl+gU1aOLar2FXAbPgHU20nxw4kF6N+JCDtxSvRoZo8itxhNGNNoTwuIZ6WQ2R
6XC3IDUKtnSy3D3t7yWxEbxesYh0SxlIJKq/lQM1JcS9pBsDwTIUxr4GZOwtXcNqIGyuK6frox+H
qBbg1m3QHrtepKOCrs/pyaRSQ/YPUwjipOmjhGFydoKACVvYutKKx07NHBgSnSMO1dX1l7wbrwqA
dk90S4eONn4XBS2clkv+e2m/7kqHW0Ix4/7yQuL94hrEYR+OVzCJYpEPVTPWPUM8ItFPmXwaRydT
opqj9ZHvT6Oy8+i3UzgN1PPKe5M1zA3SeDPjMapAH7zskt+D94jhMh3eUbw7zSXtnBEH3a6clcj9
Gb0/k/8OKuzNc6HxxYpcRLYCBsxexsPLv87Yq5AfwfiDndnhDxBrx8+9/JDQ6kfdzKhvgUd2HIOO
epjR37FxbeLbN9/b13Gtm5qVxGO6vI9n2P26QsRFO9A29UCKOLuKO1JsTcn7hlTgL1g9CCUGZgzZ
IAHQpoGtVCB44qmbvl7t+7efd5OQL15TyAkGwoc80DbzVaZeahPa7imVCkL8HHYErtgumPEd6USg
nRckbC7XM0qaqxzOH7OkSYZEvbGPn/YKZy1OCC5dzfZ2V8Q8TU9NZ12aQzVJl+JQb1cnIq13DdD2
W9q6AC2vRnZUJL739YFzRkxZ3rB0ljyQufCiGWgKGONoLbzyV1TNx/gozJd/J/38PWeh0MUEseCY
TRhdgQeEd0IiL0ZAhckeUe8YcA/wNCv6J4KgPdNc3MXg9TsxR6TQqItYXUNJQnSh/hJiPp6hbEV0
wsrTJst4gBIVo6xape8eUZ7Au9/YQHyKI6KemGYWtawNLBSPiL5OQGVkaTpabgZgSbHk6nv3aZvL
LNFx2LZSjhfp19k+/w6oM9X9aYEhrKIncRuU6nEmIX59EdPMcF3ba6qxJKWZnR6M1kiJhXdCa2EE
xVLospnPUqdCCzPTuzr0UDbuYHzrS5ZV34GENDT6wDTdxe4azEYf7ED6SGvRjhrlqo/1dxYm6/o7
kNU0P57qhfp8MB+f6VuEFC8FaQJvDGigWgo/Mi7mVOjNwSs8QBiCHl8p177h9IFr92ZiIQhcSztG
KlbJXw6Gzh7rSQYaie1/8gAtsPoNc5GbCwVFI9o/4XuyhXhSt63Hqj65cftCak9F3bUJBJHC9riM
ZhBtA3EQBIvtDUdIJw3JVIcX8rpnBWYj7T8nTS1NTHOMjS8D4n12F0nFkF2iFVv6SmFQToprUkI+
I3sPOlOSQuJA78r/XIjYsliEZR6pMeFAnOBevGJ+gaDDmzEXnjk77y/3+OrIASbnqylYY8ChLwsp
Oe+kxd0ttA8Y5Mjy6ejI3sURIl/fkePBLMFt8NBlphXmr356vXx1kfyMzlMZRrxMZnnbeq0bV4wh
i9n2ckylq76k2kPyqymimGKTnuBaVVTxuKjUzo3oJMhAc8co3c2QAOzQtCRfRESKWd/6d0thqqNe
GgCHO1XoIYqS/uu2G5tHV55eOwyTlHNSoMrmsZCDCilK1sl05+2Qm0g/1BrTib+2/lL1gQKSAzfD
vESrnEK4bzO++6YFIaTmtxB5dfCPc44yNnGFv0EMv7m6kefCv5PioFTAJ1OweewSqhp0+ryGrTCD
6p53LdRoJuV9ylTaQUknY7ooWlvDwQoT7oTkyv0djJ3+gZ7c29cj6GgE7rNp89869CHirQr0p210
tOwfWte5CG5B386m1ekmU/RuNP0zCICjh5Zyf0hb7qzKBK70U18b9L33+tHOOSstbzimcQwAfAYp
Uvl8GFNm55Jm+vrRB5BP/88ItThsuBrqSew8zcFZU6c662mYMoscgtJWAqZn1ptSoBNVrip8jdpF
Y645b1GmR/Qpu6H5HUlvLHsFDCd1LMdLKvPx19QfBBgi+j0kY0GQ/+4560cPks8EnXppVnq9YTVL
OE5n8ju8fKX56WMIivWjfCLoZvTDJM+/ZktM18LbRnnyZ6rFjR153tixVBQzIhOdumxHmqjOG333
+rDR7NepMkdAnxuY6sz3Cetm+BD6yL/iaz2Cx7MsZWbgAPYwBNyEkYTRQiWX6JztgjxQssruN3Dk
5YRvEGx+AAmLl4zhHYDp+uQC6c3BAaEgVPJXzuJlq3JrjIvt3zpwhOhlbstFna7Ivb7dva6gzk0M
rU/z5HCZLulEE2ZzMnjVhxzn/0/nA32iQFUpjqjy4tPxxKVY2lg8QDFFZdBVYl1z8JoIQInzRgVU
K2N7SmSEREgdutq+leQCLMY3YYFX3cJsphjjvuST7G3sEsOz1dMyFp9VsMpC1b++ak9kYoy10EuC
+e5m6nxp/jqfm2zlTFCuEo0PgownWzrOd0pGlpgmaQo9wml4Jloli+Yemlia0AFsl1RXwJc32iYL
hRIhn8yt0zvXs9G6/ZQWOJOURIGeMT2wfffW6G5TeJKcKIUwySRjlQoUf2kqxPMcHMj/4/B2p8qW
u0JFhlytauBz178o22C40ndcZS7Yn4c40HlQcZJo2mgnWK8JpNsZpVogR3wQBDd8FVTRWD36ZdB2
65oMC2qpVC6x5b5fN+XvxM8KtPz5zvd4DBpFNP003xCqMA2uhgUiqmQB1UZJUMEV+4WZosX9cRnS
Zs/z7IWPrfr7O5gxWKuValPQBG+kfcfuvste9GoFPqpGPN84mRvm07gIPTBUMVUs8d0zjfOIkBkP
4iKqRuBlj1x4dt21SygUeb/wEVbsXFXwkxhhA690I7JZTz1Pqj9ccNv2gG3dx9CvE62ZaVCxrrSG
hHxEP6j4w8MNL8lX+mdswdQouerjlc1lfF3T4kJxQyxkIn/DECpnprfnzvrmdp+p9O6Rsu7AfaHJ
CIPdBMcamlMTU6Px6tev7iPqyHYe+aZy5KFY8/4EZ6MnMWATg3sOQqZdoFXG+MMVi+pOA1u/fvPr
Y5HIOaudy5XDm0UekkDXT9wVnUjm3W5JlMMwndLTo5e21gP8k5NYUft09D7nqeCmbe2savMjkmD7
kgoAO7p/fg2810v6fwrJiplZQnynEm4QVvIehGNB8QyCyY9wqBjXLx3i1RdyW+9XpRefYeUwVWjD
wRznNS4Na70XE1SHkQqhvji+gZu3e+AhTngPtJrATpir46Lyfdg+GDpwSTBd+gFMigUut2PN0pcO
uuOjzweFySSOgWAVh0JmSaSLvgw4CvBilBu3GRddTBPXu9m5q+2DSFSwOjrod8jQBx9Q00exXfSP
HOOUUEaOFuwSuTPOGa7LDdOSFQOONi0HTlS5tjjPDvg7cDpvIShiqzKkoGIw4xBPa+dfh4KwtXhk
W64TJpUbvUxxZ88W6vYXh/ldzyUpG3mvAIhYWeGuQsInonObhcxn+laX3SNgLAGyENjLAqCI62sm
+jjdf4klL1N7yuqIOx/DRHAjfrWsPZeshsR01y5GbkpqN2mIyaITcSn0xK0crZ0P+gJHit+gxZw/
3tehAO5UzAmiNlmPSJN/WC/qFlko2cD4wqMsvu+Gyb4E+ik4sEjA6kygVIkC3vZ4EFYzRWEvLyjg
WfyTtW8+6dcs4n0HOILjxHDEKjqq0Lkm4wsrwkXXy5A+JKWQxIZ3sne+A4UHLYEG5vm9loI5egI3
wTGblWrNLBLn8MCu1XHpsrRW612WUHKuGQFndVZfzb4HY1kEsVHt1OPcbJVh2GlLRbpXndXd9wRv
woRU7elQ80k932Dqioz1V2Yrn6ieOcP1T1/vhV3BENMFT31wVNTZXH/EzmLcn4dxQxG2aA39SALH
uRhBaLsb4GY4CtIukfq7+tgXZgCoj6e66KSHrJAF3ohrll/Q1hRLt1UAEUG/dN3oDjbOtHAUwe2Z
wD/D9t8OpV6wgkjGAh70jONYQEMcXgV6Hdut3xeciCIzhUETLIHDFiXVaK1zT9IhBUNTUeSHiBit
N05G4k9MkFl/JTzK/+ToWuuoXqgZRxkiUdvQihkEEgDhvv2T/Qd7vW3PbRIBMknBnOWna2kcAtU0
lQCeh5rri1tP8FlupTnoPq7A22VPrysbAD5KPKnyWARKAgpLRSWI5wPv/n7FRyQdnm7TdL2XW+Cm
neURbGElYH6C72wCkNpe+QVTaEExZibOM4nl9xx2ti21y1PasvNRjOMhkyMPJnlbFPxbeHtKO7H/
3ChCTwdEAUq4GKXuJAVlTjSAe9vstWwXTaNGmrt3nMoyX7qiy3GtEKFhgxOVZjgW7T1kSWAR5ejO
AWWJPMFX2mvai25RY6AOAAOjZ6LPAmMvIfII009U/6zf/8v7GhKbgIscIWCn61NF3faZEE79zgLS
1L5ilVszsx1KhNjaDJE+otDwgF7b6VOS252mf6S20zVIxD7HkHUzWoDgCSVybGmO/chStEFmLKKb
yRi5//PlayBdq4bq5PmEJUGViM8ZiuGZcTvET2913b11VIFAJqEnMQYySlXBom+VwYhBt8FJcKb7
5cQRJ74CPrw5Kuh3i+yvpJWxogyPUPUUZBGXEK69/N4ZJ9GWCSdtjDE1I/CAhNl+8/9fcNZ7+SUo
DzrfxVovZ4XD/CeZJ7bOMUP2Gw7Kkp2rbtFUzFvF9ZSrFNto64fpXaO/q8OuSgvLJpdwfKyrW5MD
MFgUR7NjDGaIJyCGD0ETAZuViyzi0r1j5QIXy2nudxfazLf1REl5lPwiMDwmm9dzIJIVaiCw+4TQ
Wl0Ym4uG1y95Isvf6nu0QU38p2ssLWtteD8NO3G7rFOQxuHxsRXfcNtJVaMoYx3kk0djJYtxB5nn
Anqu9V/buCUprNuRWHKd5VxKwqlUa43i+r+rw1rtijonB9Xt1ulNuikknMRPWTH1ajXuIqLj8URH
q+AvcfcVwa0WRkYfalY2H/sssTftJrj2XcZZbt+aI4nnaBON+ffVsgU9JKo3cAW+BCAa2vJTqxXa
r9w47wjWGIO1swREvWLXJZg02ZUNcwX8f9LfIe4I36z6irE8vzNWqHjKb3NWj4oc5QrKVtcaZobB
b3bqveeIOrmbw5UV5slNON+SgXxKhGiShx7T5MGnnZLaTLT4GR++phcQ5oBX2L40F3XLyCtDvSFA
5gnse4BsTi7Xr+9Yl9YwxauCje75bbWCRh8B4NP/70DLmkSzImSyzISer5qN8+LEuvqjFZNsbdre
S7gfOdkiabA1FLe+6aEAnKpuUzeYLyAajya3uZYzCxxJQISdb5S+Umh2j0SMVjKuixf5KWtRBIgc
1QO/NOdVyuE8qiXCCIsYBADbmYU7TEbf5vNokKsVaQi/0tMxJxa17xWm+cHsGhOILSv/l3q4oO7P
xWYjHpBWylBzpEhIoj74SfYxRXHuYuDg8WR0obIeHhNaitYAvgTJ2s4OL9DkltRB+34WGnLRO4+5
GjfyG9OqhjdskMbxhYz9aTJNEwYrk2ntIDx2iTKdzU8uxYWNhMCLPqmjBfDcHEUiyVbB0n3cAo2C
C9acfxX2sdvwVySWe1lWDk7BnvXrwzOR7RGdOIfYQgTsuYtoDX/zlA5K5iqhq/aXnfsyO4qIzz6Q
NQ4dQcWU0Lqkej2kbpqebBXUGaeHTMS/uheGAqynKMzEaf++sUXxsY49/CjZ9APINmlSvoG+yCFg
ZhdZ/buFFWC+s3RtByKvJoG1vGinCCO2MNtjW9Cv67NLnUA8HsRVQs00OvdiGTpgcIVD7hYOSH9I
bE1WnjclrrE296lSoRjN0qsZ7v3R5HrkWm/FrJeJl+pHBPRdLw9e7Mrzs0EUHO7WOGbX7Gay41Vl
zJf4tFsjBFknrSPNuq7CbsqTlaN/7ZKbszvfVi895RhzhAM72fMu4SNjcDcROFEQszhc4ct5z3IJ
wKv4p8xsgSDlxbqWSiFDR60oow4V2GhMxCw5oBGmy5X4AHjLu7BSbEXFE6i4iujCkk/kwg6jgf3O
+NoulhPFUaKo8igzkqbKd9t62SoTrZX4tiTdXU+Vptk2CxhIqKBwtSEyr87c0c+pMGIi8e0bIcaA
U9WezVcnh9q+bgrpSYB5kFugchfl1aY68O+LR8yxBFjyh2MV4Z/fZY7MzLJg3SX0VoTBgN/xIRxI
ZmAaPZ67DIE5dCph201eP0R13Fb91ZKdfG75b75JisY67q8tJuRoITfDRLJz6Nigfbm0oaOKZ7NF
cqTBSgzH5iD4xNDjnN2pU07PewSjvEM6fAbx/BoTaskf0s1OIQ72XKn9MssbMmB+CMQFTe4skQhm
knfonWVv8+5QPeynnad+4Pxq0+0JSWJ2TUqZqVVlUxgSbLnEvcqWvAxnR0Zx4vnRxbZajSLY/oCd
zYrF1/JmTKMyGZA0/3q31E3LVJo2iWaWt4DpbPgJW1v8WlRYDfTik7wxlBFbH1Z8PWxZYla3hvM4
TDXhPt/X4ramIKzUslmpkMrnc4xn2N//hxjAAZ337Eo1ShCIN1127TBgeQacid2QZAMm9BHfJu3g
JaTCYOZ4tdLP0KIc4rYMA3kxnSbQYz3U8ECQcdPz939dqQDM+3pCorFWYb5KgUb41DuQWwZOHwWb
kw8+oYMHeI6N+L/yP9ESnauP2hKLhjJcnI8l+dc2hUfHvP9jggImqsEfOEOJ9MbPn8fNBDv9l7JQ
g1GEN35MQv22fuW7EzHd3P5hfycQKjTMj+trTYynVw6crOUxg11GLmU5FKO5p/nNpNVWN9Mn4IsO
DG3kuA8kMgRORKdb6/f64xJgTb/rnkLBnWnHD9vHiBnvujf7nxdcjWLhgAhSTRTQ2afGjWgAXUwz
imiGnxywkMFMGgCk64B9dWf53msttJGsPnzC8+/U5cm4oFcq0XSOe69r0USHM1Q+J2NZowhBP4i0
mbK5DCLfzuv+N5QeF7zgDqEka45BPDxGg3O5z7ge39/RTCynrK+VmcXqg4LrcO46PhnkE4e+FUP9
22E0KynvlH1gpEMdgDpJGj0mM+zH8YPCA4kFwrcVm2IV3sH6d1GkizKchhqQ28POF+PbphZNPzYi
OhpJTKupz7nswduhIIMXsT3EuRFic9aqsX+L90QsZyojuxQC8JyUUANWFQczC6SL3wBPz4Gfzv/I
uxM9v6y2WyAusIlS6ZvcPchXoDNmoYI5ng/M3Ya3Aufc56Zh4FVgqfU0TN8k/y+nug6EA6hIiWLf
RBoZDsFqINuAgqjDOgsp3zZsKDcuwoGdhQ1Zoj6aWMRoqGDh1wmpry5Ac+QiVROOkvbdV0wJ7x0S
saGeTFoBEVq/v/mGadrl6wg3q3aDL8wjZrxBcnj75Ww1Wj3XUDRMaEXmTL9J03xHZq3d9HmpYCs1
HBS7lxPdnW3TyaLBKQkSK3Nrd2l8iBx49/Vy9G+fgB9xFYxUtwnAEq6DGmTh3lfqUHWyi1CQKIhP
eQtMr4AICoYeIr0MEA074c+c5Q2qiuKxrZlh1x/9ysk9w0rTAB0byLb2ByMWd0mpCuCJGte126zO
Wky0sxMcyJGp6gYQtBcKM+hf1wWZkkM2jlib+Vymn5bxNnjgcNSoLW8tG0qsiwx8qd3Y7JChDE7/
H6jaEQQnnzZvec6PpRK+egPW7atZzNjFw0zFdIKplTkvH7THnY1bxj13C+IglQK1quxQGakbJsYT
v87sCl4TUsF9J9gp3yKnGx3w/xa7lLLtuiYMz8STp7mvXRZQidTovTmDFQ8JQCt2E+jpoq2qW+b6
K0SdQkOeuVY1jW/up/TjFhcwZSBFhzQsMIOv/MBk4JwqA4EsfR5CbDxjDvODulSolPbaH20NgAYl
V4dKJpH8f7CthORLyzdtrIWPUBn4aWbXuRhnbe9g7BAJ9C0Ambpv7ur5knlyzHaQioze/gEdD/0b
7dxPYf8P5kCfcyXSymE0XFW6tp/dx34pnehwmJQVn45RSb2Or+RLeyOKu84bbSrtROS/8GPQSelX
6LVeBnLE9/LglqcEWIxyCnt0mDwiLf5G+qQwt2VUfOvnSN3I15VNLH7QS6uKu7es0W7JhPobcFn3
AFgQ1ncLveSYcCnSohQ22b1Ct8aNZUK9pGEphXEyoF7NIVpFeVhLkEG6yOrSY2ChM2VmPf2haTCM
iRlCpdAtPrExYFN33OPM8F457JSeO07+XfiNd7JH1EjzstXg2jogUI2zN6QDZJHRzd8OqfUDCtGm
hJgwLcf3VvcU6i2/FHaxBxJXgbSnu2VttnnYAEhaJkNPZ+iSr011Uwdmy9D0BRnX2z0SPWtrrUm9
RADS0bEePb8xzV/r30tTycMF6JIBbBTpbkqw3itszpB26AEG1gpti7VhcJRleLn/+nX4+5tiE9pX
gL58Gyy4H4E0EdKeSJ+PX00huTWG608//abJgZRdMlZ8oCD5PxLNjoHe4l+MqqYOgVqJFpSdz4mL
R8ygGWrRbVFYxLO0ZXdSi3xCKSeDnIsnuU6EvFVXmKJqMyiMe2ciL4ucDC31RBg4V0Y+diJvQZ3/
KCgQ4hzEwhl/qCEury029f8htYioCRau2PQS4ULjGhjRyiSC3ubh4Dhxn1kUPFUx22fhtw9dR8yC
5ioSK4zbZPwdjpSxdPR5nnDig0X3j34TWeekFZnwgqA8Oj0kQ1QfaPurB1fAW38fYnL9mob/HBPD
glUAZIS58ajMgQxVINqb1q5TE8oMJFVwnGDtnkYz6hw+DNRtxxQW4MRVqlF3hwfjCafz2+WUQbUe
tRlejh17y+hwxobSR9oM8/1a1V2hvdvwUwdT0G5L3tgdmalEXvFIX+Mqkc+vFfR9i7gi8xP5WoPD
Ar87Ej6Y6nMQ+7MciER4x9S83Z/x7+Q93Il16oaEqK248Ph7rKnAJu8VxsUIsw+0HSrJGEYIRQ7Q
OO8v3wXn/pw6ng5aIKJCtnn+0VOcG/fMZHK3CqrWPfSh4CcQIzwGO3TwxULjz9+PFzSHouZl/GhE
q9tQXBuiMCARLSFoxvZOBa3w3tPf2iPycD87r5i4J56+MtT4u+uzb3Odb7X7rmxI9Jr8Jocf2Nce
xH8ZSXHNpCSwBa2jgx+FHMsbtvc7Qe5+2sRnP2h/+HXJQIXfEPBuEDGF/PABwQOXI3OXP9o/drrF
p19nBcxSSp/s90dhd+t5F23WgpROpi7HwPRmj5l7vV8IgQV/L6DpsITeC2sOnagHDuGfuzlS8xMg
OH4vZH5e6pn/bQD6nZpc8pYi1ai1aE/7NtX+iQFDCw9Ej5fcYSa8j2CciCTmj/QIrRmzmmwjqJlO
wN0BiNl1mcWHtaLlYjBI2Xo3M6xq+04o1TcgZqrX8i+I5sC0wRUXSkVvavFFSZv9nMlVcjmckcAJ
R3HzObqPFm5JQBC5f8tr4PIUAFcphsmP7xhH7Mxu+2n2GGFlpHtd4/O6UbC6NuoG/Y9R1HpYIJgm
BNFaDO9Ip0E7rZ5Jy4i3D2IQGa0J9RkwKFOT2eV+uAJjcvG2UBT54sLB4JIRKYUWDchSU4C4/nPZ
Xqa2w9mC06PeCVfK9g+Tsu6ju236jrH167h1F/dPpw+5YvS+2EB9kadU/De4xkybDF9iMZUE6Tuz
vS2MG3kda0ukC6RoLMg7cFU/7WyTIJFpyATNyq9d9jVcWm9/ezQvhKVWluRNL6njRuxiWfSyyROA
Dr9CikcqlZQKHv/FOHc38kI4LDLXprX+gsDVWnVrbakOuQdgbT7zpKKBPv3U/JmqY8O/u89EjuXV
HAFjEX751sR7qjVOq3WLCtjLho0eFRgeJ+vUGdwxhb3zIYCLCL7ztQ21diuCDZEB07z2yXQCJm7w
Ab/wc93qdqrW789p6dh5cnFQHPS8suRGedAfWrfgLvVv4AjDiO0HkVO9CQPQlKxlSRYXCgXCWnUY
28WtpGPers4IDEiouxQ/ALadXo+Rg9G+TsrGGDmfcRMSX4NcMMMD5MP+nFiiADG+WCiBZdS1slaF
u1XgyXFC38u9fkRbrhrpa2GHx8BhAzTnkh+RPbgoAFXbvWZ+yv8HSQm3ZOU+o7ap5LaD5G4Cof2D
S9gjHUGBSpC0QQprA62y/lKHIip626zJ1iBVJSYlGuZmVOXNQ1I1uSliz+UX9TAh2PPQFrVYlLZZ
1RxzC3sPCpqoniW8AkoqB7G8tdIxT5Zht6ty33gNISWGr71t32mF4oJVl3nzpVKTMoHuX0VQmejw
CWaobhcFcUBRC+v/K9J9Q++iZ7AK5WFN0Y/dDPDRJ1LR7uYwqdTXxxDfBbsOsZiO2kXsgi0aadUM
iePS7dkZXX44hS44JDEBRo1qd2T3CP0OSxkscZlnuvSOoMa92eaEEc9srsQDkLqsfF5R7Vfb0xoc
bSURnsIDuTROWkDX8NbInN37vTNPq22wxZFeYvkc+5sNrZADaCkwkuZaOuTujvXWTsPIjWEuD7C0
g/xfd5l2ZW5lFMOxBWJH+3UarBKeTcYqIHIBe2i8hq1V+oHnmQMeobzQt7aAkf9nu62Vz17Ut4dF
1C6iKL83uIYT0s1hVm+UgCyOc3IarBy6TY7rsQaPe9p3mPXhQO1ZQGcTrccze4t3cPNs/tVuF7/y
Eb9w2CyPKRY/AQ8eelxvpbGsasrYVu1KNRZv67C3I5/h/QINgnldYxMtibKNgSfHYb9I7GqlNhc3
PuL2w9u6PIjLPj2V8mvjauI+QEszuAiKdGRDQ+8G97jVRTB5C/PQszawspbHwHLjKYbxYIY1mUek
4LdLnZlNiDvfuSWFltyMnUBEAn5kHEu1Cm8fyNdNMzDfaYYyDzRBaa0CFL7VOI7JUURHgcn58jOY
LfhksuJ6DKNyLoC/e/caEqKKPZPMDYYMZd0Dye4k3d/bcsPDI1V0mSLNOrIvpidiwd6Yv5GHlaLS
cXIdyEP7K5dSOlKyGQPWnzzTLX4ZRETqc3HWdSIcE/JU0oYN/5kBVJYh+bC4Km1qmfQR4vm+AMOB
YBatsR7F2bnmGhqQJhvFplS7FJJFy+TumWmA5TsiI0U5M2t6GnEdyNDhHO9RAhypUjw2dHGpbME6
JuRyil7roQ4KgHNlLDkckJxQogppTLzvpNUOSJbJhb0OFXnjywAmWzwI7v4Xm0Yj8xPnO9HepPdq
abtwMKBbCpJvLl6+G7HCITEAsU/Q3BlUQEw4oeOR56Qm1Wa1zwDK9tAy1gsm7ROHEWiPfteAQLF3
hts+JST8xAmQJQw+4lhSF4HQyRMyrT71PuSJ15XsTm93n1dCQ4MYvnvKzG+Qfc8fXBhGIiKifCzg
lBU99n1Rt+cWOeg1jkjGacJpJIn2VemSMBZF6iAG0+axNhcfHUUqKHmMXj+Hbj4SCppTR5lZO3Ra
seDiB4Cku/iAAjIRN+t23J4lfuU/KaVCI/6XoW2CfEApqNjKyBHTaWIrMGzekIQFYGzeKesoHcwr
ZUTt0GdiOnaT5gEgMYynqWFjMlxBBUAiV+q6F+rkMjbjRGWfoKSfZPuC8223mi8VUbJYaZAZu7yC
CCAZNEGoh+PLOfsEhXi/P3FTqSi/9vcBI5TOfWlHchqhvBZnlmVetWptWjVTzBDUrgpmXu2BnNtW
n9ceKv+DjgngeusreJBiXGHRtwbH2Bgj/QfQ+ahAwn8vQR2a0KtunAI7b1M1GOoRTvvY3VheXVX3
Uw3Rnpfmv6L/lrsXTb60nvjgRbTIgZAGudGh1EuwqtoLSy0zGiR6E4vm444xtUX+h7KJ32jdLjIK
vqHm0uFiL47wZZNuKW7Xw0R0N7x4CnsNVf68O11kaeckJMMtc4DYVsPhoUSLnRwULfP2pOivQUrd
lMbe6FNKRBMxmHihJrSYsO2Ky12/cOdrIAqgW9rOrAx+IMc4DpglEKM3+hbwrozYuoJh/B2pbTS3
KK3So/8eNeEp8oyLc0D89D7aKmHAQPfqZ3RozKN6cJ0PpQLM+4EkKI+4W9fuwGLWcfCMZHan/N1T
mIT2RTujkcaCbv/7dLfXSjXPyTYevaJ4nf8/XKEups70EteqUm3BHxU5Rcv+HLKRJJMjekWA+5v4
OiusVja9kh4/bCePlBO3p/q+4sVQ+sA5WTvz0Ty9CbBqPox4mcFwZQiO4ul/MjYqpKdQSwZ7Gqzo
5SIE5ibLhOQm6uKoQykSl6CNGdsTXdFBVRrD1gxGgzp+OYjFBiE0KajywlbEcV0krYnWPCjOlAJS
B8+qxLytoNr9hBpBwB/IkPEempZcU4vz7JlRAjdZVd4bjMrmaiUidd3/U96vvSSEDRLyA8IO9w2A
IwqhZjN0WFoENi6WwTi9aiLDcYj7QsOYNsjV3SxtsJETBiLt9wBgIdt4da+UW3gPYSLp3Sgx0sg7
2Oq/iHjTxV2liV+yydX+COG8a6wB3vTDi3Qs/n/qToqNkxYTNXwfbCb93bqBhz3Jw0uSaRSDEBFA
/bqBI5VgxMYH6mPZ79Mzu65Fv1Sx2IZ+PJChbmjq4FAXvn8f7toaM/B4QWPRNYOnGwZT3CE+XOBZ
3AEDlmuNvjJQragK0EPDpHDPkyIn2SYY8VzCynUN8pBK13XTTFd3isMtHqYG3KspkbXV7wGE+U8m
R3BtW9YGZWEUnHAFWzKvYQUI8VcLWwdQXAZ3k9ilthalpbIzt0s8rChrEA4vw9HmND2hM8DIsyFs
+a0OmxxOamQZ9hJFQJ5FusxmJF4g4juY8o9JUvaMEOEED/cUKuda7ziGABnt8NTON6KNO6ZhjyO3
gj+iMJcowDeXaqwBBQwwq70m53rzoADwOf0x/0XHtEEeL8z9hrwngX4/D+LF0DwxIoli7D6a67Iy
AXjMymjE1n89yRKcZYKgwDa5+AwSg62dpMR3r1wYZbwGP4Mw871lO52fKkuMWR4nF6T13S4kMQKL
/O5UXAVRn7UzmmKPrZb34M3/ai7vMCAAybC4nv2iDIIJwSYsd0JD5leof2a5oOOt+bbcaR14bdlU
qQl+AowVDckETEbmkjqTd0nJU+jFUIUyYJR/GTTfdlOBrdDi22bH7oQByx9EEsfgfwvdu38O15EV
sRfpnuaIPqiSt5fjtByU43erUsabAXCBHL9vOJ8uh/ozQxQ9ql3xcDC/OaSGYLz/8KRWjQOUNoe7
IBU5Gs4dpFGwMox9B5iHWsuKBu3OdA6+GM9kKsrS/tiWbSDBOhaS06p/CAyzA1GmFI4og8XIR5OZ
TRpej0iULfp7DdLkQPT6q0BKuQtzIKxwnPqIuJJBwsHSwJCz46zuNkGCASx1RxDtXiM+6X7M/NeD
MNcAITMK7UHvxv4G4h410w7Ezst3P11QYbVmlfG+pPZUT1BCqR3b85AV09LWFWBABw3SEsipQeSL
rZ2Yu6cNCTQnPXynp8XrNUiLJsSFMe8Zb/vcmxKLJcgfv5z+zKqum8tP8Hxg6KcSe9y5hmM6TR99
IiIPqIagyFvwEA8SMJfezds1xKHmCa5xzO1uuc7NEgGQbvLHO0rnbQWMd2Blie3Rd1KGHt0ofWnP
rHcpjRjthAgRzTqX7i0S8gajhGcKL3WO7UhUj58rbeod+tVsEbLlkZTGaUOPHn9rBd4OlVMLqQ2B
K+I+kqzBkqmdJ/PkLFQz1P/rSxYeO9Uu6DBeH35NLgFRCM0WSQyqDj77RFrxzw+OGi+Pz0k/aKNe
n1Wi37QyJTeJpIg1kkTwla3XZ3yDuw/+OgpZWtP2Sa+t+TY08xkeuLNn2CGdsCCnxQCoytKODe4C
cV5J3Jc78uoizYtFtAolkSV59naBOkj+POlIq0K/Pp6CBM6dVj92udhXLo0SnE/UV0PPpvoK4xCu
fPqcp3MZMldltDnhW6Xv2/k4HgjFO5xTirwdX8pZurATDk37NsKCgU6CEwlf7YMNCVBYCnPYXBcp
X7Qc5VJ8Mg0LT8Rdxjy2kz/PPBCJZiBRiCOTq8zIwiMFhxdxJfSz0uS1SJCsmMcIk5zMvv6S9bi+
NmWwS7I1gkOd6iPwvLN72tS3wTi66VM3oP3uQD2A9kjj9KbLNx6JEQ2Ec7XTI3TMJrEzA+jInBRH
vtmCJmb6HQGd0y/hvJta4lYIZ6bM1LF1wsPENXl94oXgqKdgg1mt/bbB+/mQKNw7P/9+NRUl6clH
iYvx6Beh1gneWpeDDB0pOyNjeVmq7LYAiNbr6ott4dJPjZ8sicnzqmW/XTWwu+O7u/G4UhNx8MCs
kpqDIQQxWz5GN6tLsC5Os7o2LOTq3ZE4Uw/tYQ72W21fAEQJwMFGC5tfnnwpFksM5L+PJ14Aqb1E
ntw/PxOhVrDNOgaXQxPmuLaN2Iv53c0VOMpOaLA5OdVjtYNQ0XXTfUQijfjKJPjD+mtN/58LozuA
92mXNv/2o6LVG2Aet6AXD8J3OywqmzgRtuKD8VyzEhJD+Arhpk2cago4mSkoS7FO85X488p3wgoF
AtMFBk4HODFipxk1ysgo/ZbLe08k1XzujyrkFhOsmUEbSPkkV082qGoHH88ZYcoubC6g2hsrV7xh
ZuqUjUCVLo+ljn4pT5tyRzYAMA/H+5f26wL3dmnEmTGFcBaCYHBysl2Bj8qiPlEiB5CYTdBMeLlz
e6+WgwEj+0K1m8AqfqNZxrvczrW7xpE+J+HzJSGiskZP9umxTg6JLQlXe2ALCx5/fxBPbluB7/9r
V6+eSbPtlCxTI+1jpOLIklvvzZyzHqzOTFsRjgGI4ry/1PoUZmOTGIgRr13AjOwiVbs0A/flWEQx
L3Z4/DoR5JHSOzRA5QnfMLz7ml2HxaTv7iZwy3KtxdlP6XtnV5F9k+HjwTRBVnrBtklrniNZP0vR
Mhbm8pZLkuGSBDtf4XqA7m96c7LA0lG9BfTEN/db0hKwID31gnzRVj4YAJH2F2dV4udEHUNhNtlz
951Y86u4PbtyobMXeOourzXWHNR2Gp3mZwwOQspfD2YT362wZ6Fj/n2RJwFZOsNezpaAuYGrRVtN
lHoQnAIOcZ1oKwjRYuCkhzxBoSfhkt1O+y3U4U8TmnJ+bn0NLKgvaKttmULkaYPhHzkBVuuPz8iE
qR1cP0RMtf/cPId2OxhI4aqjLCQKAlrEO/a5NmxKFs+WOSlOZNNHeTVyciFEGCAh+iyVCqIiQ19S
iqI3wZH0HP+UrKaeGd/dGRmoPf09h2ekUJVOscAGR4GQhp3xVH6cd14pyIJkAxkCFcCsXhA6Qssx
Cx9FN1ZZGhg5C9lugaX/gJyx66Fu9Do//IZMMlU3jXX+lYInj/jOyZ+VEYuDNOkVeEGFMC2W6D+Z
A7AnHjsZ8x8J2acKRIZiLP8aNv3qotzyC65/uT2hOxfG5XIQN1W/A2BP9LEmS/MR7PkXaEWyrI/4
v2wsPWbg7Jg8zYUfghsYo1atBUDpXynCrMmDPrOxU8pV59XBULGJNVTmSGCLhOIumabZsUqDWgwM
MDTrX4EZ3RkZ3D9TKIZAWQj0bwHd07iy4mSH/Qkww65usYZHE+OipNOOGdsRYBd/2AdV4vG5G2h5
w/PcCR46kADNWLh6WAdCJB6he8HuAoYda1rAYZ1o446Fub6KX5fRsYdFb08swdiRqCDVYxCw5g3K
ZtmnE+CF3JNC1HW0ldwDrsvJUOxJR05dP+eBFM9K7XteAD0t4UvZcaHPVW1CDi94qF3aLkDwBRtp
zvv2OJsVtSg437t837XDqv9SzOImpVu22Qv0oio/jZpXDmz1MmTNzBm+hq7xLysdfyWnwdvjt1rM
sWei3DmwGe/u31YMUQ7LWlYJTfoWNLxcdAEdQ78dqZlNJ/sEXXbqEvkYX469AfsbiKRE+drufehi
mBvs+0rTViGbjvUUKCfXtSnYaPGfqcNgt/uyk5wgy1KqaYUhbLuHI6aBv4euFOMlXFZQU7EIbXjo
DP9hdzbgMLS5DBSDSfGOyi9vti+7ZTJRRSCTrSPu3G00ZcCSeB1/65UBxFMLX52Faq/GwWULs3bJ
jvfxvK5WF0y4UyFR+RT8oxbfhqFsALC5k/oAw1238eByrB4RhfzbiGQmLDhBci34j3OTAOv9Qg71
vx8CrmbE9B0yP3tYmEB7grOXVSbmh/zK5eV6HC7yiYZjTa0SCmG9zKkdr8j+E03AQv0MDXkkUTMC
CA0ylHxUZbvnrQ7U5jTXBlEa52N4LmhvBq1hSrbYO5HbJvWC9S3/cSlgE3kadMkwPtzL2tH25ZAl
t/UdOURdyuatJcT5Slkne0FTItrG4Jk1u9aXnVjyzbZOGcSlMhvJK0R28OJMJiwzRisflm6CwYqK
Pm2eT05uXlQqgFyS3biWTSJkAxmo84arukanxXqKBvcMN8mQi6YV2nJwPZ5hI1gmdlECR6bNSTJr
AjLmDBGwMHbtS/86TwRSzEKRmIcqIOCVKhYpWEPfgVqBEyzCf+9F45e/wu8qwjTzdmeklktcGOzd
b7eQuspc+/DAxbZd7XxaKe7ocxVHO2/KyVfUmZAzLzCpoxaxS9nVa0sZz6n8G82P+FsCefo/0cXe
GoCT+1QoZ2HxndZQ0B4DDFHgDKYE5uMDqgK3zPWDj1PdnSaCQlu/EUqUJo02jBNqcYkZIq/JIP9+
N9zipm7f+SBz0fkkq4I/XQw6CafGceHhGr1wWqcyjHGpWyNAGWxeJ7wdFsLf7krHYqhXA1pqY0Gd
AiY3lrSTUbylVIQT2XsvGPdA6OJiiYwkUrQdXXLTwfkGLwyiWC1vDgDne9u7P72tdLr5cDEy4O9o
RFnMBxvdYg9NyjhQGif5RrDaghZAkXRGCkaawI+F+vium9H5tpAYrymspzTmkVBnk3xi09BFp4Am
M+bVUvbPynVFnMPN94mJbzQJag1dgzegBEusnbVAjQdn1RGupHVEHopuw4X3uf1k1IMx00C2jk5d
bUcM3LF39tNewP98IgadF8t7twQiOthPXXxDnMCMUNrXi4zl5uARN8POrwBhbYJBs9fVSMbInfgH
nx+lxuLR94E/cOdOTM5ornkI+l3rdIOjDjwU5Ym2bW6KMsUjFyS8HfjPPA8sf8D/tefACNH/gK/R
lXlQivJHdCi/r8bLFQSRxYPeW4sf7+fbuJvq9R6UgA3/Ow2Dtw5i4aGPd7j2R/YoFTmqH+VzpPgh
Tp5oy2frezP3PO9ooBhgJUBM4VKTVs6ofFjSMDaJAm2cCxcrEEvr4MtqScWTYbTqGIwUdAwlj54K
HcPXd5icmj+6AnyAn2JSJzf6egEDoagxFKqNjtq6FGK8zbVvWtyDOm25WMeXgJ6vrP/naKFGvL2a
D1Dsb/q7n0B4vt4xfcMy8mKEkBrIrNXwKh3Gdp5QlShxFqqPXnFwKkrTcXojF/oLL5OskvCbJBGa
oO2+lRbmJnkP88n6peBh/I/KWmF4rEKfGS0PcK/rABvCc096gaPYrqGcYShSHRE3ERoOGrObvuCZ
lY2ChIuj0JGiBF71JkFdspmLHafiVko8FYUGDge52JdZXyRluv/PLLXRocHZfAnz0BkKNV2JONSF
INYNslo36aZyZ32WbjGceuInSfzvbcNkrC7R5Tn2AzHFSsfYjQ/TirXrZ76mFq5vprosbyIMEXoZ
Cnfml/nBJE+cvL4bWP+LnjHHvZjAC9YYDWit+wEXI4V6nn2zpXw9N73NeG38tlorncI5xQ4WDu+k
pcrJPqDjPyr+lOC42SDsSMuQqIY+ds1+PtQInW6ypp3G88zuC5ZH27KkPi/iOlGpyVIp+j49U8hF
jsw+EpH4XN+kBlquiNjXDuJ5r9IWU0sUI8w9xmicFYquIXI7Szdqlab1lKdCURvQaoJjFm2eZVpc
BU0ZQuB5crPyZvpbzyHLgLwcOJrRty8pSbvQ5KGygWqNTWiwfA/A7UdOxwzY36Ha4wzKMq7O6v6B
Zv0GpVAS+bsF6YgYQP1Wi3Frk2Of/ufv8lz3Rl0ldCejPMwYSLOMIbhpiQLmX/942vlGmGVRbe69
iVeTtiICihCzbjJs3suWj/e/cHl24lDid9mb1p/KdW5JAPeqtH93fzW6NWGLWTrwuUzg+grUwt7H
HwcCs2pEfcfpbnmiOrRNL1qfkak1ob3wW6jrQPkK1YRf3HgrO69opwR9Yffg+ko4rnkNNgIT3bSm
DuT6vW9wCrv79suBgl8FxDprHuGRWejKIta2GHK1sRjQG3FNpgiokIVE2elokejvjT1MOmnhlOzs
3QtPc8YA0sI7eQFull0CpzeIIDPiijMajNAPQf9Nv4d78wWrcZ4zkny7JJKIAVi1y//enQvh97tw
3O6FReVz8cLzxVuLNLkuIPp6uzYOfdkS8djD4X10pfsSHLijSZg/3tg1N39HkQL/zOqd3dL3EN15
E2hXFX/mA1rpNEaVbckCje/+y5sFSfRaUvNjzn9rT+sTh5agFLr9hiTBjrHOO33nx0pN80T1UTJF
/OaHDMAOyPP3ifEBKgOH8lrsczRCN49giZQlNZYbtPMzGGF9TuIFjPQcGIPV26i/Mz4QIR/Qq2xv
3ailCztXSnKFFfVFeTQBRievKh6ayVuIhp3c5SOXWvWmXnF7q1A/retidl9f7fTX2M0HDhU7m7rw
D0YDzSb/j4lkcQdrFux1lVuOLSCtO9kh6pjwByKif7eYMVkHuLU8ogazYV94MoNiS6gv/+PH7J+a
PC9POWnsnjKxR52Nry3NVgHQ+yiDPMMqtxd4P5g9gUlfZOFFX20rLk6RfKEr5gQ7oreZUItUL0rH
F8IH9ZcD7c2kWY/wvnzUrOfG9R15laOJvivVtvwnKfhOQRd8SNa5EXMjBMNuP6bs5I3ylv9k5jYb
+ltSrh5gMxQFBpQUYKl+CUXRYOLFQbdqI1RVXxHSUFMZ+YCYxoqM90G+PzYcWNatTuHbvYfrYiYT
YMOilfsUGLkfxQvOdxCotkQ5/ZSWtEaWcZ4MCMzBn/d69bWBCT9NKYpZKDB52b6R4PUyyXo7IZU6
ua78EAlpekBpGglzGgpEgKlG3Hoy44AK7FnWm2XPhs4W+mC54jKrhIhD5XGvhO7GLMCoFLF1rWUL
lXmQu8Yi8NkbM84mi/Iz8PJ97jkfJDzEJ4QgUvVGk0zjmHiG73SPsc8SsWlCh8cLN/bSPVlIWzB5
hmC162jY+t/dYMrawbsAFl8tYUpA2p2R1jQigMusQu3vTyBI0YVFwNj3/eOdj+3y/1JJOPDYL4eU
GHJviPVdgKYnqU4Ls3gbJc2Xt30fJ9/XZnxARYDSn1frbo5CHBwX5IYEKF/ST5vbnl6WqkGKCzu+
hxLaQioftNsWG6GTTIEP9TYKV4Zh2Z4K8oSpFleyIlhoV4wrMZ6n0O6bRq6bs5rZdtOuXFU5RZ9/
42kGUxlsnm0lsnfWwF1PcYaAJKXLZP9k8/TEVBe9FoZSvoPTEBgktz0vkA+cZNWjXcUdNTByzqHl
4FY8+4LiWhqu6AqkHnoWbjbTBBzLnoutpt/7XFjL7ADQEIIzaAC2emPPpp1J+Sc2y0Mz/OhYslZw
jOnD0juA4R06fgkBtoSoXaMaDsGSKosmrFSWQjJTUH2fi6/vp6Cm7uV/cIzzihOiKRPsm4+WqlT9
/G42XPT+Onfeeq0e5EBtThrvqZX9xJDXzdz5mL9ub97QK+BU2iEndAYElh1ygFYgDN9tkjieMnei
GHnijgZ5CVJckScGUhShXCuH3HwO/nDYFOuWj2l11n7pVrvi+cl/ap9rRRKHC/IhCAkprIU0hP8m
OQy/9ZWkzPLO/gRDf52hzkuj41GW7E6DIIgFUkLPoMxQ8NpaI54Pcz0KDosCAMZBGcdVBeUp9pwy
wb07A2ZrjEO3XuWrlVlSUlM37ges9KieE5q0KE4jouDD3gEIPny50v9EZg3g8CoWdG5tSVSBJzqi
ENsSlyWLdZK5wmHehQm+39v6nt+nCRNKnSATgSYKwtY9Jzv/4Bchj3U0eKPSAn3zMC5jYVcjysN2
87f3OtgYGaFH0uAGAPYLNY5cSbUJ52zUof7hJTF+R4N9hPjQ7XIGW6mUX1pPtAra/wHBHOpUtHxw
ebo8dNxPbRozv0uJt9ZGzJJgCyRGrcoPQ4wGeXcFQQyDl3ZCZPYsdCi7PKhCIg6YHSEmkz48QeqH
uX4ZtMgP5aMLfYgbQEZwU0nzdo6esw57dyoJ2uF6bXJMDZ76uzwyixwlE1TJbY2t+MhiWe96Rqj+
5PeQM7ZrNzHD6jk1EWRcnYlgnMNJeMY0oRlY/aE/UAhNH9MNeaNO+nAIbgBlbFN6QQ+sHRpi4hHm
72nqOddjiFtnEVRlGrvqV/9mPY+VA8rtOt4LZjHBTBn9WaVhcj/sdcGXYu3jjAvZmpm/db1kUclM
iUq/vSlPn86JAxaTy0gIAreuPnTT8mJ3Q4sUs5wFbkWIakgKfU4J3a7ARLyTKRrXUb8zAYtWoCng
lASR+zgePIfBzwIxlk2mWb41L7SY6yIZFPZSdzupKFzuV9nTrVxrbNN7bRmaFnqUJgVIVDXR0lYP
0ZeTEKI2MqDaiwwFRxjauyKFa9xgrpc8Z7m57TDMOmAaH+C1HoRglOI3LFH1QlaEwSNj/MYvhWGu
5D0x7XcpQAmCSk4o5GYsnv1T7lnnCgoV332VzxQ3Ei1eirjiOBVv7REanlOIMLn0kOGW0Dd1HP5W
Zh/cDyDUVIotEwFTc1Oz8to4nF0GzRsEV5IbMc9inQLG0Cb3oqy9HfOnXq1I6FYo51UgdhHLJNX/
o9eMKDXlnwXJhvgu24V0E9eR4GEblqZPGLq33RuBCcwBdAeDwFX+t3kD5XJ2MqABYW1zMh4N9xa0
La7L4FTfcBK+BC4LRP+6OsYnPlY2zHpg+3tviuTWGmPKnf2t0vsqwcgb2Y520uE8K1yrfuT91Yfm
eIa/DmW7hFiy5uWHOAJFrSWI3PtnMs+yrGwC2Qc82A5BuAJsszDP7oUF94+fnZ0jdEtqMbA5/iy6
S5rpdtskqBxFGQqDpbSAC8tg/lHPLe+2/R0Jj6aUkYsKLOeNrn5AVZswinUmVWj5BhUzNoZwR84S
BpN5Oaj99drvhHr5lcVr+nEI5lpZamQIAOlp2SycoLixnjItsyVlgUEhPNyBKqrXYm+BW4dqH7z7
6PRfvgr+/rgExPClIk7VR8Wij9WQf/9ACxDrmKj8IY7WgAm3VPMiWziwa8yNwLPddpErKg5g0Sdr
hejJ88wAlDeaDFad+6Iv8eyIigs4NtJuNlSFSesaPazQ+CJT/Em+5NzxtrCypREwpvFyuFVXfg3a
xt1e2rMNDlHb6C5TzCx27htu/cgAwup127WKKeXpO8LdjrpJbMWviKOfFWGoiWEGCLo+KjOKvzxO
z5Dt7p2Wi9jXuooucTJO8y3bOBIFXFKs1HHbZOZUAKcsFUV6+zBPYkwyu7fQz5sKhop8VbFvkUtu
P+ApF8McUlChiB7mZZuum6sfxUrRrZ53lcLWVUtene6+QK4m7VRn8HClJAGFcrB2BMI+08AHK+RD
/ygDGhfh3vePLX727fwSSyCLuRyAXXra6zR26RKrCF3OpaVdf6Ou//O4Y2MoUUugkvbXTFp2zWXS
XtDKukL2enpApePRvoWLq3TtRVqhwZoU30DAolxwskDYZWV7aaiU747X3vEPfCDKLX7BETGVrr0C
ocn6lTGqSWaL3r10PkNsqwR4vszuH1fJNi/KRm33OvLBjb7jUefPvDEdbLpKe16i/PLUf6GqZ2VY
pSkj06t6iMyfpbVtTmm71AEvHbeusOqSb1JmBZp4kYIvDjpdIB7n9nZe8a9FdPergAQ9YSpDewXX
TM28hTuy6zalahRDUdNgdxvaVlWLw4mvYI6thx1l0yUzASvS5Y0J2C+7EQEuOvRSCkVc5bVksy0V
At2ApgSCxx43S6qCcO8X/iVpUKYhx9jLUYs+JAwqOMS9r8rlEFDcc5zBFHWRsN7SRpwofP2Q/Nrt
x5GChTO7nFgHh5n2hZQwAsav5gpxX4CcQdaKVWjYUZMuNGtK50/dMofi9W+exagH8ScwkeltowyP
KOBtq32JvMwFaVk+lSUkkI49amlyBvAm7LspPwGp8QNPKFIJpulHxCy9BMEwO701KChPb5qBucEb
2g9DJT8bAoArfLireeU0RVBj7XarsuuIxFlNhi63R64AH8nXzAP+28cc50I6DTPftyw9s2mWoxyr
qWamOo535HFYCD2kH7EXuo5j38MO2QU6JTn4PWBypuMmmhpMIG5H5YojrmjNr1M+vdm5NYyyaeHj
ZVTaJI5eZotMV0wnRgT/WJvhfAVc9n/xeE7lN3mTq+p7VXZJFsGnVohStMlqiUeu81JhvP+aAHgq
TqA9uOzaFE/aRfyih7kYTfhtNHg5zbs7uRY2zbqhozq7MZmXP5ylK+bTBZkP2z6ujh6UMuOJmI9O
FZcpEnPw0vxjc2/Cfb6jbE6XrQk+im5cmteHV2oGjZDogN2/CGqDM+zgkTw4YjbJETJVV9cMvAzI
/8LaG6bvZbVENz2vvJRQFEd3m+onNa9mTy8N9IV9ULmYYcEpbGdWvnyKbQ2ewiL8INHTnJNV5oz9
kqjgpX+4reypc+Xuvaq1U10UsuXaNWoMe5jAHqTrDCzTgquoK/9X9S4VdpMShs5qHNa8wKFMrikx
19lottVhrkVDMQ15O9GTupowYlA53c5FzfOV4grIL//KgGTF3bVC6+KfJjtpkZ1d0aublKCdl+di
J/DkicDwUx3xc0SuOYkBaKxmGLOjEKSpooFKGWD+bGS+GrMLSxLyMRrAaiIBBeLzSBKbNPdgNewJ
TpoKvtBrUUmIkRUlGuajFJojC6TrH03D563MQDB8LNw6QADdNT49a0cdkXmYFQb9J4VVa0MA0xD2
QUzAVqNiTHSUmvZBUJ/Y81SkdP3uZkXWdoyy+sM4wLXfXzykSznxMxHE+UR+qWrrYsQMkMXzWpNd
g40qweFoG29ffJmrf+V8a92wA6QkHlMebM2zSUDusDz1JUevmyYVi2fTf0rqoVvcGyg2qH8D9UMh
0qn3tI/bV3aju3DaqRRg0M/i50xypCKmyURCtLJ3wdiijoDqrUaR9CePhawT3pIuO+g4S6UBhVgL
b1PJ4BY1VMhnVqjqZ9uR4i5b/m5CBWLrlkKE/zHYLsZunfz1xBZZUKAihG9aa5ckHRqBJOnyrARy
fQeA9DjcgavEBzhi1AZ8Ut0VJL8u2U2ud2oqybn7aqicAjkoCV4DK5ZpvNVtulOZiqUE7bvYG6kO
OcyQDgz6fEWFKhwefosT6S/VGVSqs3WXdU4vAZ8yXBiS6KzQ7fLwV3vl0JhvJpM2mFlUlKEwd7rV
BHN8PY1TTZzZMYTdWPtwlbZtmjA1bb9lH31jnLk2P/V3L+deIv/GJl8cGcZOXX2I+xtOA/exLpg8
GfNK4MIzIg6FK9MetUv6Py75Js5RPn7/InE8EZMlUiJGsWrM/yw7+KQ+qYOsarccg8K1/P5HZIm6
2FFzn9gBNQTaLKPd/JCxufjkZ2xJ5VmwTA6hfX9Nddu/BgkqgUG7FnwIrNMFDxziP75unPQcYntS
AHKBzW6qBKhc4cp2TeND1nL0UC7e/kMooNz4ZLtp2SKHwmMw0Qb6hI/Sb06Gxge5qFhKGeQ0QQFf
c6MXEX5jllhTicOhgNb7AQHaZSIH+Z88wWTKaIYajhrVO19S3QHxauWAvyTF4051sldg4mGd/Ysk
3LYlHMv9KgGTLGtdQdzUz7F07c7P9/VmCsFw902Ina1KDKGj318ao2FtTzKQeHcqosOp6GHvkitJ
F31TvHIaqTMTHMXi+gXs54llOABVJLXtG9xBT6xy/bPIeDGWled+otI1aXn8HpFUEnlxggAOEaoj
Ijmje/p6FgnckWQfIhcZwx5NlWIfxz84lGbNS/xSNB6C87ZI+VIvPUZDn9m0EbjSWEJ6EGAMO8vC
8jwh0Fwu3BPbTyRS3Ar4Ldgpxz17kchfWImfogNj6ajDOFL90auCeK/g8Q79CqgId0MTuJ5uJkKR
he+K7ouIW0GrwzrYbgZCkTdjoQeVBZqlOoza5QiKYyMsDj+AvUmpM5RVoFN6sxd/cidChSjLifcH
RRcn3GULmY9Fh7JpDfdoWfXl+kLuHN57wKs6cTvMxSw6IjIlAIfEq2sJAilldJ4Ba44RGK3XTAdS
e/HN3NkH/qqTHXB6KgwjFemnC2LvAErrUieqfrWKRmDZlfBvLbGBE9j9zvx/PBxzvX+hMJYXs7oK
hlH/BB/IfO44dPGrbYf1BkLCwm2yG3SeAGndtEzmIAu+U5JwV+nvbV6rTSzH2Gitv5PWaWBNkjOF
vIROqAwOleSsMCjAy0w9LsQVuyXVmS9KQExlnYy8855Awb/LZgxLhjxZv+aeLAbVUxBNbgYPEwgv
4Ha4HQwoJgrwBZaQnGagSsOIbzcU+z01nl5weBn2EfESAc+40ZgRcBgTPOobcXFkKKbaS39MUbm+
ngb4s1DWkS7xAzRKTD1f6Epw/9amBGKxTI2lIbdOciqdo1re2dbg6IxeoQsUQit6IlXjAKW56x3j
Qt4B7V0RO7l1ip272W9wP9KfE+wmQxf/PEZTFBLZDVWg9jJGjKDYVoaLasmptFOYfHYMveDPYblw
MwycvkjdQXl25QLgL6hW3EMYePyCsu5LGU09cTKPfpo8ZGz8X6x02V+RV7b2A6XJSD0XVPAA6rEy
3/tjKzLwmr1Bdl2MreNeYw050RWzCKpZed+5Olxkjgc48QQ7LRF9YtkQ3fHpIwWRlMh/awzdSJEO
TmPztWVF5vejqK6aq5JBQ5TaMYq4kI/2qUtmdrdp65JyibQskm/Bgho6AHjfXSq3PrpQD9FDXTuY
RaJMEEYvsDdFWBinXrSqKKA5DgP/X+C+7gNRbd9PNqPyjwULy4EQoaKT2o+MwmSar+LzjODyLYgm
etNpeqcAH+hv3mDd+hZ5enpHQpkuwd8HYZTZEsTJb5sHIHD9wPTrmpTOCT6hgoEUnWbVzWHtoYLL
YOf0HF6OcwKy+rnovVoebXjgcWbHtW9WGLQqzAtddeyS65aJRug8WGmsBS+4J1a4zm5mSgoEffBT
bJxCJpikPZBKoPrUkfASb8XtSJEKTdRhEuovwfF+PUSe42fVXMpoGFvM+7bZBOajm2hxiAGJ/TOn
H7UPFSkgRU8o8nMnWB21qkNrui1/2mtRYPVK0oHzt7+bnQEpwavd+gTRqXaZNfb7z91tfKH/uIEk
QptPQlXFvUv7AAKAcPKwu5IxnoF0RT0srQLRhZ7BSU2FhizCR9uC58nMbGNY4dLqhokWTCa9NJAt
tpPMKufqzVpUv6Z0S1aBL2GU24rgS0sQbcvuGIC9nh+7Y1YcbCf8Sn9FpHoPgiQQ4GxA7X2DaJxw
qp2nA+w/enGNUfGICpEseHlH5dJ+OPt1AraGkCDnlIbl4pHw5TrPi1blwNHoEWh9KrfMI+W+gsPq
30GmVlXc8FJW+SikoUviN8KcRAt00io+uxJHerRiMRgRybrX36YGxLnB+OGGsCqjW9AhdXDgltUn
JE2GEekLhIvVDlPpsIw+G1x20aacP9PkAdU7F5l6k6cDIxfqe8MT7JOlW8iGOnoKG0gnFc2g5F9u
jCECHqkdcGc/lEVE4JquNhveOsHePWwjVUMBKeg54POyce6QCxR0UA4huvYn1kKD+97l16ImVA1K
HezOhevHoZU2tm6iUiIAKIHSxwkKlkK03N0MVik10gMQ8O5N5hK2RrMEv1VDQnCVP4pry4upFXVm
6vZlIxPE3bwMElL/ughxCnazIOUP16IWaIv/CGJhpqc2z+3y958Vr3YUqqBGJzJqCpje4oDW5mMY
V/8YAs4xBphvZpLzI4BaGGx5k9QzA1Rs0Xfpkap1BIMbIYusjetbQtILk5YghTB7rOemKbe/8QTy
SYseiNMMC/kaRuDLvGC5tX/InkqYyvY2k22DkphVvW5x5U/TAc4CnDcW7tRQuofoH9zyrE8LQZUm
0/CZC40L2c6EFItY+eThFUeuxgK2CwCnKNXmOsFdBGC1t3Os7mfrW6cAvSCoiadsb7g2wdtQpWOu
Wt3xxVM4hfRVYEnaH1cPiZSjYzXBbMHbsgVUwwrDwSD2GJ0qv2RD4OG67kz4iCozQYJgB8ea1J2e
1SXPm6h2rY8r7xjukPUO8PQm/rjw3up0O3QFOZCrRXs8LgZJqNBwh7Me7+R2LfYGfcAH36q3ADka
VyGskguzlDA6yul0FLvmor+iCc1uBMhJ0+35VddiMgypdswrQY5nU8iU7CUGzFAD3uvdxqniSSjS
Z4xoKeNoQh0G2ybN6mBnpTHXP3UF8mwWuLJ8eTlq+JkqjXnDYlO666tSzirfOALAgmY9cye0D98C
avgatiGDOXjpOW/f+hwHbj3a9MMHGZmQ2kd4KP1z1mxO5Dxq8hBqLzDZwQx8bq0OMNFz6dlmDJK4
RA++p7ExtMAKGBDYUfz4qXhveiqpnMWVPSvp84t2EQEAWax4o4o/6LzquP/3kIceDcnGAIPPp4rw
TC5G4qxFUNTm3pmwAdXh1f6+V75tAoQObSE8gLRpyZv5sctyZaJNg9I/ulrtQj0O+GqYGl3ERxXu
qqFjfOk+fP2kWj4ahIucKkX5NNYShhNMTSjCs/gT3//n3/rhftujvwYseVz6hw9bh/Suk2kDarFF
ZtZQijtvx7ax96G3LE+3PpWslhoVwx95t0/WKwWrGFwIpo/eK8LHo1qqiNHwtHX1VY54REG4NeGv
1pPn3yak1CxK52ViCEFe9WAFrJcfUmcjQ8IIHU+6TlZjuellnd++0C8cx1bDgweQNoxWHI7qL1YM
UNtPQN8dXEc+xCI2yP/vn2ph21WTv4VZ7TsiATZejjacvkKpUv/f8sN4m/PKvOXrpPJQ+Yf0Z8Ia
VrkLZMmX3gaV6eZH5zNK5lqJM7Z6+ylmheMpQslA+s0kZr1c+PsLCZgciEpTavWIoSFjskWVgCgn
9VA0NoMyltz/qklxm3mJotMIGZk2XgRaX4+5eO3X0HMpJt0S8n3ZQa9cL38z4+AnnszEUd1s4uYD
QNnO4a7rDulYGD/Bt9gnR/KfWgrY1QZWphBIqjQQdx2d6rMttd7ThxfLx4qtOVA4xjPttdw8eNp6
KiVOocEq8jSLHSzdZEfSeZKQWVuGNfTZmVzE77b9KVO5wLcjJCDgwrM62dAip9f/ZUx0hc2uKbEv
h0bMU5pLLir1YwHI+Mm3laDt8CjuE9vmk7lLY+NPLenRBmVtLqBURT3i3gJb5cXdrRWO1I4CoEOO
miv9ke/6FKIbP9HCdPrQB1+pl/Xkk6myomihwFL+Hrz2tFO7t6ro3Cd2prz0VwZJQplKL8QxFtA2
Gf/5XCOPwKchqGexgLE0amBlnnHqQe0/YZACxjGt0Ds8urMd8QGw8CIA43yVfS7d+2O2994OlrWH
CWiNdobD7rdx8olGfF+uRrdRyAFGzdIIHvh5asRLwOdIo2Nno/Rgx5vZO5ReuO6gTLM6eOHGwqKY
jzZy55P6CHZzCl3gcDT0tbgFdvu5G/GHYDm0JVjEQhQYcMRAmRXxfmziKnCcR23HTAukoJId5g9y
+a1pEIrmxoQJFXYxwEZ27uXA9lkmUw4cQ3RzLG6M3229tSqeCL+a+EcjJ+AWTdo6Ds6nyWnz0ib6
VwV5f5hwMMzqHTFRKeZUVYLAXYFCZCgRmr7HQGh1CVwnjABGz3m+rhY0AME+neVmlUo78t0comoq
Do4SRsAEAJBCqLz8DLHZEoloeA8IGqSLat9xzhdg8BVP4Wa2HyiEifxSUG99/DRxx7XkNWUpspmU
VxIxwBcM7lzJW6FKDc0WfBm2K7TPXyTv3j1QN0OjS6LzHCzsljPL+L74le6dVk0G+PBAm3lXRl2X
erK0HTJR2pzttcuLtkZBuT3GRQKQNQAIo/qL0R4JpYilBNY1ora+6uYeMt33QNhZvV5nlqlV/Oif
0CTfVtYRINcv612dFu4KhwL6O30kuUBuDh3Df4Kk7Pcfg/P0CnoTK3XJGRJXgFUuae8OFzAehcMK
bNx3vHLSQPx5b9OX0To/H+kXG7kxRCKMUePQTtb8C5BaMWbCyoy3ageYFHz+hwHq004BP8yOiDe7
sVfGa5LNiSHOI7sxOvaeuCsYe0X+TLjIh8NQeGVciDJzWio/c3tBBcP0AC4qXptq7m3SYRj6hKEz
PdWnjAf6cLjMFxb2z+Xm1X9ZNfrinwy4Cis+v7bHzDmaFsDVHScGwOa5QlkNKH7Utc48JXXMN0NT
x6+BBRFY2zjVuQA2ZNxJkhMt41u89yF0u8DtRJQx+BCsA91V21HbzZrhseL0sKR+c+FG5ap5l4fR
LLT5t3+gsrF309bBLZ/t1j89MvrCXuoAGvGGxR/maiY4bZ20dtSvKZg6eegl507HYm27Da6un+3S
GPkmFHPCKzb3qBrPyXgSrYU1ZvQjX8wBJ18aqihaaYdzH6nBceRGEBNZFRSyOznkpV4pAN3Rn034
IYB3Z/pxjGegJJMWZh0LsWrxeqkKFjuR8GkoVgM/6zMU18VT+kHVbOPsIqP8DkyZHxXrtHOd24kA
Y3dXSX8tDNAPuoi/LESrdFxc5BBeFewytCttnfwH5jNcDYyPliGowMW2rf9QsYWtRp9S0nXIvMBj
8OLdyuDMhqoVkUbg07N6E4llT5SDXiIT6ZcGAd3SDtlyEwCXUjKjds1yytiCg6nDfolG22u8Fsp0
LWWQDux/UJz+bKlqVe02FVtmOG7H9QG6ZNjEajEqfD8+ejPIJ017tfYXefhjfU+borDo9I0o2m76
kkXsMJ84An+W6GNkPBphGrtOZPTz7O4U84sxlbrcGeM6WKdB1KpNliWxaHUN8OL1dYCWODTvjN/y
HoYiV8mrECUGrspwCifFPonogX3FdcID4A0lgYhkhUC28rM4bem6UMP1YLZUO8BGl5b+RIHivkbb
0mxdvE/GwquU3H3/9m0JKz+LgBHffS1mn47+Vxa47shelyjiMSnay8s2NIvBoUEsOsKtGCkOb7t3
ahwc3NXoTIaUdlovcSoxOV9KODsXPb4Y5TQXf1OUrE+xPBflVVUpTMysN/+LddGI0z9L5jNwQt8g
S/zL/4NC7+FeBcDKDApWCztO3M00ivTJdIc0zEutlfdDqRwdrbpmwEtxDqcnLjTSzloAq2S4spTQ
pyuUlFIFjhx/JVrOhB3HN5KJuNr9BD3OkVufQ3bBIpTDzaILnz+FswnnTMdi7ukjJMvWzLJ3iEz4
cAmRkLnrCXWN/uvW4EVuHAcTsYY74l5rWGPqRjHgjrazwxLzVIdWUiGQcF8007bqMDVYCaqN1+sZ
v24von4HaxBwyKcX0qzgaV4ZZBvAnycL9pdfUgoiAmKsOvnKL59JB39E7PPSfhCjD0QPtbvOIaoo
1PgC8RWg/Ijg8+xWCUI+ZusYegY0HWTkA6OxMiSZ0vdH8uHsnENjXPyh6YUClBDfqznenZlsu5+T
hjIhMEYznLdCDzDuTF3slBHv2FkFzVYPhCavgUErlXwwet8esYp4Ux8KCo7cqp+58EOAncVKf1tl
Mn577VU6kkU2Obdnzd55bdSC9kZmMwpUp2nWgE4yBLknP6mWsV69i08kgRohGkI7rU8nlid/ckkp
XmuYR9mZYUpJ6ZVlwVCFvYF6s2CYGZYW9AC4oXivTjkGo/6LjSlhiRGpRaFV5JwLDcZK8kJSzKr/
St730ANYyNH3vx/JUIe8cRwVbLJZ5Zgr/Foqj23TU6iYv3dHU4Cdf/F1ZMAVmtsqmLXgc+HbevOs
fKySr2uEx42znnUe66jHRa3WLaF02GZKu/khL+ImswpBmsUmp6hQG+9XFCy0LnyuaMjAh/fi45tk
BCrK8aj0D+fPVhIZ3PAIxV1sFfzEWouu3TahvnDggIugKl0SkFvO+wuiGiy8putkryZ49YslPF8K
hw3nGq0lZuAnzyEhLpoMlGGVDoYSHN0TXVMyC+j48OvTqGwFYn7gSDw9k80cMAIpZvRrqhnfDCpk
gAd8l5kvT6sfrAyTMT4bEffk1YgwX+iCSs3AD2pyhGbCZSHFKiOOhwXUoG6BvpBkq9Z7Fmz6/RLL
dWy3sa4zoRYZEImHsuS1MHcjj4j9Iof+qaq5p8+ZRnhiii+0mQ4kFvbkCojTCfQsltgQT2JBXFvZ
6TbNHJS9TRBM5DoFQrs79G9DfeNpmljFGeU91XkeFcetf5/aPjIc15zxzS31IwGV7r3BeB7eFGPL
DKMaNcvLTmdzOJX352pnvsVTbxefn7UtYL77KYnnoUrCbjMAlJBkQh3sreUM1mEnknh6fXH4jnmm
5m6vEaZx6jOwdfYw/Kgk/B7P46CTjHeKLqX2JvOQPksq3LFGpL2Og6WBE7cqPg9IecVntvJg8bYn
nxBbuGBqdatUBI5DHIMkhb58j0XxiQhP3kkBvXqLYTm7MqoTOKxEetTcygjP+/5sL1Tp0Fnj+Cs8
Rz5XU4Rad/HkzlEHmB94KEvTPVCrTvhuRxsrjmEGJK1pt62FkKhRGn+QQJ8tJOymnO8jweemZc51
S+OZ/3XQI4DJQnJrIxPg/4NAAMsRKS3tAWaWd1bYmbxmcKwg/WyYWplZ8nnLyWiaCYmsvRJ1FOsy
UQMDjyXQob3fKCXyy6Yn03068L9jFuWluE91Z4LepYhFSl5PiMNhKp3URjWh3+84te9YJHQrkqN6
yF2twe+OsstquR8rHD6J/KmCaJmDGCcgVshfc6H9et4y3iGSJgh8dA6zT3CQTeB82DxlNky20ql3
fnNiinrevdxa0fP5StS/NjLccAGcdWkdHH2VJiYL/DCFbrgAJ0du7QjfnsnMoXyg1UxFANoKGTEY
ovIJF55AfcuLvafGCOCJCIFIBBIl/ZdvOX9TvMGdZdbFZFhbeU71lTkqmsB35+rF2MzMrX1nvA31
yM2KczxtWvldn2ySrgjUDm+5mCbgm8A6JJIPnYmEALSBuc2Peof7CAW3GFEykyJndm87pOgtkh7V
UE+jbD6X5b2kARBenl/VUhm+YbGESpLT/l7Clk+B7WNlazBURgsdRPsN8mZN71rBYhaDKnfgrFfL
ff9znctpDET5o7Gp3MuHPTkrz3v6zpXyHpxI+CWJkriYAxlGbk/VyWMQC1aQRE88g0wk4nO/KM0I
TnYqpw5VmuK/zYGdTcN9BbyIUPYa4b5+pZR78uc/xeEHMmbpuMk6AcNZ42SjJ1GLq46kNlzkcPiP
6SZSpnESlp5L3k489T5b8yx8kuznp58/LblKbO+xAq700jpPUYUHgCp0oRU7sibQM5+7UJAyd8tU
1+0ETGgnn/cOlIZN3N2C1OOSAFwXBiqBSctg+YhMt7Ty2EgD4wU/1fVcN8W/7EUPzYi8UzS3adnY
JMo7o6ez2Do/mRhYGiKpjNpoNZelMGCDWEyIgxobCqsj/84SCxm2D9nQM3IlrsUwg4KzHrXpO5f9
LPiVAk2dYKkGOGtsrwGm37e010mDo+eg60U8WLlxyJigX5BrtaMSnHm8d+FL4CBowX5svi+XVOpJ
uRs9Rblt+TlHvvNv8pFBK1SF1q8KNke11Yw8jMLNb+lQA2ppkID8hEtUacNGLGPXf9h/PKgEQ5Mh
jjTbfoIUNgdTFrqWqCMVdvjz3d+lvg/4bXq+ynagLBCtvUskxjBR03mj0vz2mJx20Hf/zBj2/8T8
STpQ085Ex5vGs3v4xN5lG/L6leLNLEifk2yHbL8bkWmu37Rx4U/mPVDO4bVrGspQif9Y/XERMHjv
PcTJy1LU/eAZt6Zv63pfw1j2BZ0bmCjtxpH2pXdVgn651Ho5n7Z9/mTimiZ0cBe80WsljSKr6CGU
waIUzu66oQ/t5ZCYsKub/0Ff4JN8SIZjUPRo4Nm86GEul574nf9tshfGLxJFvsbqT0QADYbWuSHN
8Qgl57LweqlJml3C1I8lKwsgtlMdlj4UKQteFtR9vO2KOWZv3KTvy1vxNt5HgWr7pZblRTOdCESl
lO4QWVYRiMooQhP3EFvgTY7h05e0rns97+xxQTnxAQqQeDl8QthJDN0TXWOv+X8dsnIh1JSWzMXM
/MLl1Ne5hI4JQeWtEE65Tj5S/qwrPqLYYvXChjPyJQ13M2xmFAjQBJgrfdVPEC9KRxrE6PedO7tb
wfqA+npS/aBgtsizA1K19cYbHVhBm/YK6yZIJh1Zyrpc8roYYRB5sWQDxPBurdcMzDqCiDe9uCLQ
js8KLc4/XXJ7pnsollxwuE5d6aDQKBUIny//uFj4eWUw8/nbHmEsY2Dc+rZKjKO3fkLgrKGxRMvm
BDBuaPhk6NduGUmyO8zJjxLe60UsUqo5vHZvEhZXW/wralXj+Oynz7PAe60kFjZMud+oc5fQN8oF
lqwrJs7STB4BKsbqtiBGVmJgxNkCV1mQMCO86/JGPhcRHWlboYF1kL7bBZPEB6LoAw6HYsrPc44/
qtQbiSDfsIeVYQz0fVaX6/8wTba6S67s2cOExnkGme8E39ufHCNo+milBdM1u9PfORbv1q8TqLT1
tTTV/hq8aaDTsVMKpu40c3rx2RUhBRHvSi8BgsFjTdChgAutd11/qJXBdEh9Fb1wtBR1f6QwcwNm
Et8uj1LAoq2jnyWZu5lqNr1OmYRNhV2EIrE4sAbvHD9CNYrlUoHvhYNzRy/S6921w2N5QXeuHOdI
pyesCjS3i63fyNHaQkUIMDa0jCsS/bV4EDA7Dufx9xAiU/eu8Itaz30XnAOMpV5bfprON8ZzZlqX
dsgv4dWzES8CGmpLocKgAe19isBfpnVWSAUkXEE8X0ubgMIoy2ez/dcrpN5nfbR+Wl7tIPacCws1
OmZC+mHkujnbp1VUvl5a/UKQkLr4zPTZJiXHmBH9NAqfxE++k8kRaHb1+uE2esNR4e2Zx3Mxyx9S
viUkNWxM1HHl9sMealaLXau/sT4q++oHcdD7XGqMg5KWkPL9twghmtI3ubztAOYYbpsjFmwFZruN
i14HmoIZzAInygTNnMvX2oiWW5z48zuQ+9RQsPRKObtI2b/OZ5e/drOftki/kweFtoPNDsiOc4VJ
tFCEL7x3sO6JeEsMn4T8krk8nKuoxWK5c/tpctTH4XZ6ZmjoEC39HZxwvFZ1jlPSJv2HrZcNtb03
/+BMl8KDsu27/x+LzSrw82FFUNVgXacLrE+ncKd0KF0KauVUYOoaXuXfImtV3ds/hUTj48bsjJwz
RAr1/Sxano1P91EJyLAoRK/2Sl6LFbAQJ6e2O6GFompcBXCAImCJnyF7RYcyGCID8h2E9Duys0+G
3S591HEj7l46SMMsB1wwULI3vm6c0iHvKZD74rULjL+IAMYZ7ndxEAw5OU/gkeh2FJciHsHFpO6w
DMlHGnRf1NX6/pmC9n1ro8NfL/P0RfyuRwHT28kdWaNM6fWNkGT9YSp9yMeSd8ugtgvOA22N1wEA
ex+3fLSKLwbHZrL8QBzgzjC5CIJieID/DIWG9DhtXcxRtK7q5TFvxnXZZTbTyBbmxFVxHl2M7+dc
cqCmN3Ka5/kmuP9HaSIo3AukN5SgwBhc1sqyi7/ep+NlW7z2xMHkwxP40YdibkDsXRyGdcuoXTXX
vapxY6gjPTEjCTZqpZxd6slMIyN0oGQzCEYMfq5HtJ2TUZ5PNhj1XoK6/SRZlhc5vkyZrcSdNqKn
F7i2d8y3mwo6OCKQdOLdRZhNAMV+ZTgh1PVLSrMnQM85yEzmAFE+B4bciv/SAAZs5RcKMPEblVbs
52fGSEH5BPxwVdkyX0J52SbLZj9c5KdowHsCid4htN89cQ+uDXn/rZ/5chKOkP2ZxkJnEYwVgbuh
9uHGexlu7StAHSibjdAXep+8heUP0IQEtTn93IsPA16HFt7fIYOWs3bBCKa3KgDFMOi3L88Rwg+J
3g5F8mv6X1ebMoadONIONbY2e7TKF6J6wCbxJqpOzPf+EFID731h6mRQn2ux2wof3FpSdPEmmcHc
xcYPnOqpsZ0wGVZ3q7ykfa7dlpSqwS/FaJYSnEMadwvdq9GnmkpU7PN9ir0JFEjlJ86CkDFSmHQs
mdw4vYMuXIWOwpBJy2VekWyw3LAsn3cOYtNlI63LatjhekQyS3XrQ8lnq9Ddk5R04InFITD5zKdi
Vu2NGfgEOPbsdK7c2GGu7D2YHLsL2IWOx7OrdzpkfGF8RXBBmIZG/ZcvEO5Kmp8UDvEvUbHD/N8G
SxS0UoBNiz32cpYcO8W//vKt2ZsZdk/MwAduZznsSLX3kFAp3DDRO7Eo40+zaQu4+EbUjzmRlW4p
ebbnrBmcFDQw7nZglcAJXJTPVu1V0cdsHjTMGtOMFXL+JrI8jvp2AwnPlvgMUjkfZQHaQUFRipOq
rCirxKohYhVp7Sg6EFhXFAuNlvSrgogo35CC3mqcO5v5RF/byvpRWqO873TDRAtkCjr94YWG95Z/
zaOi8Ada3sl2S7NojPz++UkSEmmpFSPqKUAmv1GjrU2Yi2DyJr2jkhjoktkIdUUrBoFvJex5gxOU
829Z/JdwWtAwaVxMsYF+cvYC1ca3H5HXa5UsxJkybooCF6D6R/hJEDZA2SbODjXyvER1COxrnbus
ukTE20j+QfGn7kFQiRUBDTp20ANYo/n5hDr+g7SHHoLBdh/nYrC7LV0TpXZdM5cx6dzaKaIB8YnC
gMQEFsHsktoKfESTAScD+zA352m9LRuQAP1iacqRbeQYeDsuqX7GLvBC33tcP+N88vuVaMLlDCa/
jb07keYS0Sgi5t9JfxysjydE5H39HM3UfEreIBMp9Ma5bKjYDU3ueynWOIv3a0uChOMN9asahaOv
iZIjQPgqiuD38kf8lHkHjZGN4W8mJzriZs6Dxc0GhKMJnbgnbWl7ApEtESn1VIR7+naADPa53VOg
dDTHp9T+WmxT5VX4NcF0dyGYLEHDcp7zhaoHZwE7xprrMEqkAykMEHPBCGOPh80NZk+JbOiaTxck
f8LWL7EsZP13bj9PLX5cCf83tWV6LAcOFjGNi293IX8p8yZAQzSYp3NW6zo+uhxWlGnuZoBXwLVO
ALp7I9D9kDxwhkmkYG805f0Z3bgjwnX/QVP/kGdidz0j53kpxqsYljhREBP4AJ3XKS1MsK/S+vIC
NjF3ylcoatl9jdlIFvhOmKcO3r6dRpgDdynaNcQFW1FKWAHclF2TJh498BKNfzaAPskZIwyAVv88
+6qB9r+GRE/ZgU/3dUYbvNr+oK26lSYP8sM1LmDAJKgyTcXhV2GOEGClBnAphFPlB40vtf65l91E
NEZKN5kacX3wiZMgesUBhFxL+wgcjbH/bgizBBMstc7xs5eRlg/T4oR0WKG1ocUVCqQvJ8WF6Dqu
sb4eT/lHS5z2gp/I77j3Vd/d8gUTVo5MpJGD8RoPtxMUaj1cBVCy3OtL2/cBe6vkBd3eRFMx2CLV
oRhrvC/bXMuTcYgLDaC/bW/7u6G+0GonAymbEV1jfhPI8oE03nd/PuGgTJvrlpxNoAtFvrE6+9FE
2ZkWg5bW9zQgU5C1Dr39WtoPfFQqiD36W1tIhdFyZC9M9XSyogXQGZLCOfQo5lZ2INHX424MPt1U
r8WWWGhOwc32y+ELtVkSPwGMl859ZVzLqjdQCwiGci3yoQfY4ZMkF5k7p/aNIsry9BrQ8UBhkBnp
BbSAsAe1Yp3hfNWLWs+NRXKe2qg7kxKVKZVlm8hl4wGtL3l2cr9f33rvo2N+BUvqygFHKLqzGBYN
NGUa8X+dLY1yL4fPkoTzYwZFJgT1X/FFfcUvoFZ5oKHZeYlAQWzeXBC8c4nygmb1Hk5CX6NS7WCg
PZSlFKIGCgEq5EqMeBnL3nC+fio6BMIOgYdh6R0yX8AefQZn8A7efEfcg/0hINz5+mcR3crJTjEq
mpRSq4Om04mtuLmb83V02UEiMTAJ3eDjbVDBrW9U6LDVL6ECJ29rNpt8Yv4i/weRMFUdjIajZAZz
tqL5TsY4NzgWg7HSaRdTfypAH7GTPSwDpr8NLoRvvmIdm4kE9QiwrXBXYd+Yel6Qgf+4ka5dAT/B
5EAYg0WJ+3VA+e/cNXotkhrCqHpab98tzU1sYfS9ZtlUNTxuYFgT4sBeZHeDQWkXZLsFPtw4euFA
1ovH5Vr1pbu/Rk3uoia8bGOgqneiSNI/22RVe2M8xcKjKvnQdZWs/s77qf2OMIcD1zU1DqOLmOEV
V+KyWruD2Bv71XGrhyhe1hQTUg1eBBeenwE0xZpy0pLR0njaF3AeaTiv7brDG/gDAZVaRH+aKqQI
e6/64LEfZMnM6pCiMlpujt39od9+Hx5LHMBa9tBjROJDdSutBpTaNDfcjpYgK2rn6AmFInv2Bpd3
6EhVZuDSFGm83t/9QkwUzC4xae6NBVVdSxckclkvr9R+9PojeAggm1SqO3V85yDItPy2dkxrbjtm
VjyDOKeSBScM4FXKh23J9fAiMa47FkZaIbXDQMqzUNb8y5QZ1yGCtIuM7LX+Qw+j52UdE7cvWjvS
het85n/vkXha+SK4uKdkNWZLu12y0kaInZiqTIaVWAwS2QR3tBDDVfU4yGokU1EXISCOncqpeqdz
UWLYL/ncmBkSW+3i7Pv5jdhweo4Pa7l+whGxp5lpdwtMetjn0ypPaTJ9vkxt0sgoEdfTQkC/g2Gr
+WqWWltR+d8RYFyADi9JahD2vQTVhgSkNbUyceAnHGfAMOCXyTQ98TkTBBCaDGtziTfjiwxlPm9K
VVHo+rec5tud+CJPBYW4VLERMhS+P4ntjIAYRtRleDVYSv2QU2tM4eHeQ29BNBmSrdtYgtnNagxc
OPN9WljMVHYU8blnTRv3c/Ri+ddR1X3bsT4IPSAEGIF2c614jnuZsjG8RprNTol+hgeJ1R5W7uTR
jN5AStB66BVREpRuJ9rK+Hszgr3WEqYbu9EvqO2SLk+UN4QjXOmhtq5zBMoMzQFl+WaHp3wt0JsF
sINne3KQzCsdJV+zyfadw9boQNXqiwSREwetp1M5zpTqlhYxg+voN/wL4sZa8sCXne4pdiVpXhnf
z/gf0okyCXXsKxbCI28HvWOJc1PCBYcpyWPBT2BX8RoIljCFB4pgKT/v8NZaWhEZWYOq1+UmNWt2
bcVCiuK43qL5n1bctxWhvhtS4MWefDj5RfY0LQOAwMw3D6RvUUb4B/ykfUZqxFWZ2YwLBqsWB58q
Np3Uwb4KaMbF/gCVFhnf8PrGDa+xPxthma+b+Jxga1o/LTqGxlGNEWxcnma757JM6WawjF8ME4qG
Gaqq0TE00jPBC/oCe2hO1qAFYsYJWt0RiTciaG+jGrMpuRZpUK8kKQKKAu6DC18C6knPq2m1gGvr
IcSdu8cOTqhRRebsMxea1wdpi1bqDFMb9T/o3ggZZPdk56UtyTP1GEcrGZ1hAg3LVMF4ixQhchAw
P8b0FDEpCnAz70la8SWSQnQvHA+1Sx4KaXUfnqwijy8Frb892UEn3Tl/mxbKrqF3NG0H13Q7+ZVX
QqilrSGfctrMp6RkjyM+wNuKT8wxI3fC3EfgDUmi4mzzLSUEG4LdXdmYFm3NSZJDHvLIzzZtBZVu
DEV1Goixjc+PNHWfLYxcEwZw5lgQie5A9009gnqt1KZwXrYhdQZkrmgF8YEYG6ftzZadl3hoF2VF
eleJRnTf9PcMQngwJgSBbND9SBiIefk64gThlr0qSYDc6GYBa5OMHPE1ak7iAomQ9rKuhYH7/yS0
IWeL7u7tYxRAORwweruG7KbVn5kQnd2IjDyAN2XyQz7vuMVBMWaXKjo/uf2wX2ItUWasI7YwOdMJ
aucC4JZikeVnjTWk5gAtQMTE4XoQbYcyHtVfW2zgs3GeJpBNYuiiurqmp58NTUZgZI+VDk9bZb8Z
uHOab++RxYrVOjKqcisVsnBIx0nDQ71+0Ygk0bZgeKPD3xzvi7jbQO0w+Psc5FcSa29dYkvw15oL
lDqEmUlSQHS6lSNa0mIRPeq9pnjR9iTjZknP3xlZ8xHB3FByJHAHn1KRWtaamOhBQoEZGNOcpiyg
7VQyxCqMZsyUcponDrLC81nCPOB6b/c8Q1A9hNz9SlznB7GldfQxyhXi0TNTruzO200/qNjiLrjE
xz3jLix/rWPdZcwwbjLwp9KLbiBrIq8TxG3hNeamGF94qreONCDvkOBsxZR/PFlx/82J7dHPKE6A
Bn2t5s9cm2ZfPIsom8/efb89E+xA2STe26cG5XEx7O6Mzx9lGYG8DnW5g2MhjGKhBwtUTOiS380Q
jQ9RYiLSvxo7xvuGjlA2+WV+wvFam1Wt3a3BNvQOl1SCZqlrZHOLs4xLknV8g1r4S+8hSo8PzZP7
SbIhEgLeaNh3yYBnpka7gAzHfU+0JlknbFX1D4evagTjTfyc9idELvh0yW4XA8rzT1UEkrmwkrfO
kqDaERPO2dWOr/KEhbRCuTv6aglWyNiMRQcbrtG5lwD34e4xRMD0qGvTqvqoaazfj0ExXIjczMRC
+8VTXGBqfmGtbGM22S3oAqtXL6pcC/NDxKoZb4uZMQxybbZOCYoqMc8NXkg6AgmFP25vLtrkNPHf
SinmMhdP0AWuMcu9v3ayf89+86L18IanHlIkmwRF5aNv9i7SJTnkG9AiDykkEgagLDWc3D+sdBsd
XJ8ahvd90UDg9DZDB05PrQSAljF7I9yftlsESI/w6ZXITP3UfoIj5vPv0k2Gq5n3zON767KNhAiZ
OwzUjAI/DyTDELGuiooIFPNcYiCgluFfQNzlDWKJuHqXtsFfsbHl7lee5qlqmyE3euJ7vrRaJ4yt
KKgiP4tBKFnSCxryu1nXmLHgUdALjuuUYqM65WTebkg8IGC9gNzfEsEsW9LpxbuarLPr8GVYKViK
hQlY40366ejBp6MIsvIHjbeWlqyc9m+Ctcec9xY1LsQ7nYdX59QXqkLpToKCaXSTfGo+EAHuwBiR
6JouYYNwH/AdpX3ig0aa+p+aA5hWBmQkE3ChWO4gfafCYmXvxIzNXWA2fvvYGLYxkUK+q9/CXt3l
xZad74pJKwWhj15VypX8nl53hLslNr1+TVbU6VxKrGu2cDnDPpIvAz6UF+EESspVq4274fkrcot1
9MO6ddTnJ6utjYYdhcDA3SnYCjhshk4CpJoSLGnF8hbGSxb/TWvX3vUFUQtei+P/LWihyNf8ZRTn
YqnSwXe+ZnRXuCJaTYaoCOvhwnISA1CKt2sGCsPkIMK8FDZk+mpwyQSMK7/uX1PiY5QL0cxVlYE1
biQF0l+YNcI6y76pvMRg6fCT64MjVEgsZc36RoMkzaSd66KO/b+R2rkDv8bCiZjMQKFkWmCEF/I2
Wt7crp/bd1T9G69I/IJQkD/ZelM7cySvQonzs1hbVmSU4mOPj3BfA9BNhf3tjnV3iFi+q5zjQblU
+XlcodosBXlgLEfAtNyfao2omnZTPKU3+k0EO5e02GvOYuAl9JIfQRih45a/y5zbiBg3Q5NF1zB+
TTUO0k3ujMd9GsPf5Po+BjVQasyP+BixUH6LIjn0HlfQ1HC+WrEBgudDT14mobMqAVIB2XbkroXw
iC4WFNO/BjynaiK/fPT06eSiiEHFAGXRGdW9d/KUsmdXvQhAuJNEJPIsCkL2XnKUXLIF+SEjVftT
qRll3HnOmbOek8uLBrV+aRV1Xp8PBS4Arj5Fzz58c8Ve0LnvUQECriME7DVmHEJhbF7MQEJUvalu
0485i44Kux8+YCoe0n82QVc8uxd+asAtXIiz3EmFT4KDCPgkYxPjpuHyAoFyUvg+vpSctRhAJcP8
MteDsUiL/LuZl4gHc5mfXqcM0n2DCyiptGvXqc0If1b6hhKn1ShtH93ruPinmmtLtE6wiX6Q2V7P
+oP+XiK0MnE3gW7qktq72aXO9RnwA8BNXQtqC1iyee4YyPihboCgirOuP3eHbUoyBwZpnjvoOexd
yRq+ksRaB/IHlJ6cfD58dT1iX+AxEcUTrQKSBJ2Oi37ueJsN9hlzRs/R/AhtQNfKIYc6bYEgXm2l
a+9LZfb1SHwwGqnESAgInhe5KLrdYtnBt94rEzEoNvfafC3JgXT2Z3y1mZw++JzDgsZPSfNz56AM
WgXJshNCQmmPEW0t9hdd7zU4Ppd0hAAfKAddePmYPC/doDdqwKZxsAZlU777MZqNVhFEYi07Hfq3
kmPOe18XLgzhnc6l9RvByiwUM2MeQUjLDTKnxJ025LfzFqCekSx7VhTEWayKwWEFLhYLoFIZu8RK
2TzgvGKKZBv9qaRevFTpaOeGbY5BjFpC+mmAatfpIQJbN2xtSgtIwV+I3qZ8fx9VbId+VUtZlf3P
FB5XzRL26B5th1SF+NYZYCxXFvCc+uyJAK1Oo0jlCQFOhWVoM2ToszXNzJ5iROy1ev71XELwED2w
1Rwu8vqHdEy9Jf2IH3Q7YqMhrRyDMjsuhN0Dq3PzcY3EqlINb4JtRmw4PLScJ12AZP9meStklGCc
GBl4elA9j7b/l1st3bOScqwlc97Aynksvwxm2VQPZC1GVZIXH94idDymm4HEcTvumLHE02bZH651
qeNsS7T3pyR1XOcuUbWnUgdqXySpm4cWk69sn6i+a7Q/Xij/OTUMU2AT5kGpYvaRshtRUWG36ABs
lxPWoFhAn08w1X+BaSi8gyDQOOLC0AcZt1fr0OY4NyZyzBxE7YXoW6ZwMbVs6knYuSSJwDpVo9cb
HmXYYHSSQgBOarZ+3D4Nf2jojvCo/u751+pqyzsGLddIKVT5pRzr3lj/uoRRlTjRF/Kbsa63yg4F
sjQFgEJHBOjTKcgpBo7FgYxoryyLR6Cu/40JuSdyJhC5SvGAQu5FAsYvr0xopS4VGu7ZmDNH4CyZ
sIuukRqMaMxt0SaHj7Fu1akgyUwSzEhV+mcMILfmO7F/Of3OJvrmfpr25PzBWz0EKsbRB56gN0Cg
2QRM9xu3Wd1nWg7TyZQYNh7tk6mAsM4v9+4/UXnIcGllTinhEVHjzeHnOvVyWecBJr370G1nt3/m
bgXbBo9dPrj+h28YXk5S9lPKNpU67BcVI4ifAW/CvagcRqsnYO9VeZ5+bnXOGRW8aC6xCrTJG1qz
YpgXnqT3REx/DmhB4Rms8h+VUCLJqX1SKe5YQFzbGLVULEdRsSwYbiRv17bAotUnRjpZDOl2z/67
qTMqfd/ou+VsONEH9LsAPM75en8KGir3qYeYwvy48plGf+evs+mVjbi0FmkBwLmBDUOs0jvPh9JS
9nnpQ7Dx8Oah/zR9whWgwEez0209MkRwy3cpu4cdMYtnQOmGQcfD+E+IW5HR2qzvX5qHSCTNZw3f
iZkApseukFVxdSTaTUD+lzrEU/rI31BnAYGPGBMleW1wdZSe8Ozhxm/p3GNiIfyYAW2ZYvDC2Gki
zJGWzOgdIIV+bKA0N9sk1nFrdYMbh8IJUoO6zoNC2P1wVVIciDMvi7Owo5RE6u78gwfSSQkNpHXA
YtZxtEI0bHCmc2k5TIn/pU4XC+joXNQsHyGExCvb0KZljUxrYDWDmFuPbvy8wCryU9tYgL7sbbIR
1CufMN89Ar8bVz3tmyWE8onTv4L2OT/Y8aJ2rXMDKcuIvzy8AWTdnAAoPxo7oGjp3Xu2AXxlKZ+w
NacW5Oth7RC55MFiRWrKLCAS1EbphrHBXTiI0ylp9cMn5USKn6s02DJrXXqGD1zmT1ynqM6zNd+G
980vJx5PUbbWUdvXQuUFeIUjxFWXdHkE9CpNIjxs9fM28Ylabs5OIb49NLRYIfnZFNrIkcEASft0
egiTk9sjxw8N5+6STFnqfcWA3ISW82Fr8MdQhVwb9Ha6SsgJX7O1tA6P8mNwgkmoKeXbWzRVNi2A
08Kfdvjcj7l0WpfhxdI3X8zaCkp/MkWWbq7f7TTyRF1MZqg/QoKVXE+EoQJnB3CMNv/8qP6/b/ww
cBZ8kmnGM83PZhG27kMbpwqO0Z8VGClLuSvcYNcCPF6V5QEczziMIhyMOfI0bS4zOcgYUmGCZsAo
be4e/KKd0t3vr49xgXILMokCiaXpFzYHK+ES06+KQWpUgCljsc0mgN8d1QO1kU/Og9RpNcsc9to7
05LrjMP6iaTOZLVEPc/E06Hmol0LPdG8M11VN57/HFUizMHymK27la1OTtrPxLqxSnuWKj2h4ety
EzgYTJjSo6V7s4qYKaKPGsJzHV/hKZBUk2j8oRUMrcO97JPymZFmBUYDg9cT4FzeVxr+4gaOdpY6
ENS4HLl2fZ+rrqSe9hV+uz0qqegEObl7lyA9IQqioBcq6FoJx6z88exb3agbviQssN2GvsupcXZA
HqZG1Pm31hX+hajTnzrq8p1TMCAGOXgoUq0Yk4rwefHGVnXb0fQdd+cAk+/Rj/VJSFPDu9RHG1+g
9UD/a+zIjoncYvuJsM2uHxd62Dvi4OYEgNvwsg3GdoCTPwrG4rxYWd09pGu/TBRAiIrnPvS1jVj9
AuIdwYdEvqJKdccjOtsbQjrdJjnroPNLW6w8mSjXS30507Bm1tda0Xb+jeZAoVO3X8xf5TLJ9lgm
IEV4SC+ez/7LBJZ0ZCsSxhwXXCyri1EehGqzgTv4Np/5XCqNQnWCK8BfANZ76QTq4mCcf2yi7rsk
nqkyzZhvdoRe9TTHJFC4qU/sKSJQpKE/KNRDIlHCThqkTlSthQ/B1FTMpfQEZb2eANqDzyzw+txi
iNsJvYgPDHi402oR75PO7Wo9ol8uHLZc9D1LVGmKN/b5iEW5rdZDM0XOliVEjLGwlZ2IZoy8Id1j
qP8rc9RB9Vi2LnfrJxLLZVn/8aAGSdVh/8nZT1BWlzuVxVLHgYWto+0vlykjTlKRjFGByLNcvK5e
ER71qXQd53gI1u4Az3KqnRXbmX/6VVNpzgu5jjaJBKB/tkznTOkHVnOQoFtHhZAMagbW7T1070ez
TJibXQHeT+pszdT7h8JdzV7W6TP6QYL3b52Ib1NyyZIGF0eCfA0ZVW0GiNbk5rVT/9Q+/msFwiVZ
VPc5LJqPq8kFL08rzk+6DrZSEjqySepHYwAXV3BisX4L7IjzSjYjiGXgKabPTASogTiGR1SLBOh9
AwsPSjWHVvTgSp0+X8g9KVzwnwoJZKzctUXvyBNb2URvUVMRdZ51cCJfBAhv4cDiv10MZvwZVoYZ
Rx22bCpYjIy0mnTqaKlgJqM3O4mVlbD3xIjy5XCyYJL69aMvHwB+FFuo29RmVea8zT6XoPHHH2e3
4YMnCtGfYOmkzQerq8Cx1h+r6tFop45u2XK0jr7GzDYkqWqYhVtaeDhXKc2344OdXs/RqymQXg+/
xXHf187CfOn0r3DpxvoMKk3i4ksYI/oRyaHWhfRCCIo6qIifY30kWawSlm+oS6JY35TiYQePPh89
HRDfetWuUKLfk3jNYlv+tFDLf/40Iz8AO83aN+jS7Ei2R68D+iy++/4FpaFzrneE/GwIKD9qlUm4
ROAY76AXA1t4KsyedjzeocZnji336exUBFy9aObnuhlHgC6DHxUe+gazamAjR3vbEIXMsz45Lmtl
DjSbXCnAe+wJpcD+FJWVAt5WRIvUeDWXWEhqzZrxdXVgfKlf8j50RwHL82HbwopFfrr/+gTVdzp0
b+yxYMWtOStF8h2BaUi5JcyMqomkM0VWgQcfT5fe7SIcnjloFaCtv2CZuc+jM4cvWmXl9r/RkBmE
gmn/VZR1M49qYkpoHVB4UUQ3yDTGNG0xZFltZo9qytRaee9bBc1ogNT6Ozekf8hM677uyMyXsVV7
82/k/+L8Jy79x1n9GSikD/l3KIx8LdQTtYbDrHiGoo7L5vNMavxOpEJKrMX9XdWaqTEH55vQy94m
xJkaPMD7tRA/kYp/FiYpSIHeLgTceQCvrVP8r3FMPn2kcsH25dEGaPyAR/P4r2MBtBK6gWS3byuU
62R8uW3gAJWHvR4nvf6ScOAqv5WC732Y+84uwjSw7gKd6vNtJYm0NL5iVavUCazVFH0n+6LYTshz
7QeG6qWnDVGy02nTioVa+kLL81yOf4VJMB4LdYVSFTAtprUTRR1fheyxNBXM9LuKET6z3aF+WANo
WejoesZYPG7cVJ8ajAkMWS0IIfdJs6mFJPcRub6o3MZyeFQq+pDSCz1zY/QqbpWnGvvoKQTz8jLz
IiAOz42YC35XdsSOXK2Dm5OIb53vYxP3SzgZUN1g1l31c23rs3LB3sm21YyqyC/5Xg7oGLnzuzYq
mJl4ST2hzPkCdld9b1qIBfPuMSoIzMTzgKoSxzCztFzmk04YPgBzZ0jtrn5k3yo9nEAY6CDm7br+
oCgozjgKvrxhcQoA3Jsm8G55l0KBVCbNvJEEh4QgBC2IjWBC3eR+VhHNWolKgZN57Qd/ADiSQ/if
Wxr5xYJUeKyQ5te04rcuVJ/fpeFfwpHk4vL1uaCZQjgRjZp1/MJuHOO/LgQiUnN+WnlkbfPG+N3U
ppIFM2a1LdgxPfWAc8P99bDPIY90NY/jsvfxMVnVxRaRz/gc6w+807Sa3SCJk/DdeamNE31rM8CU
SNDrhavuVEPfAgAKcpfvGbw6CqL2LuIBVmvtMc5K5EUADGtXz2Xx3IGNmymG7/5HezCalMJxGW6h
ejsIZ66Wj6GRlvj8yIPLfG6Sx2LRU5hq/CXopnGqD351wvbqsq7zKM3+TdXoQHWzUZWm2edURpah
38nnlitxHw20tTl5vhZRW+L7hGDXkEQ8ZjK87I2D0uL5VNJPG8Km+ILUxZG3Cv/34IdM2281Yms8
SJbhqNwiJk6M5VNoClvF2W52oih/4jf0SssEN1n7Xgq2bArytPccCz57JM0sHOaINzPejEBV59yF
RExgW/STQpg+wXT1qL8EQVSLJOCmvdJ3IkeX+iOXE03fLsGQ0qpmSH7JAAqA5f4e15x195kRAwVy
7EKBXkJvuTj4hDmgcwCtotMbXal2VH8agDg85YVQ7qeac1muWSWk6yrE+IZ26qLQhDOnHJdSN/o/
JTW7fWEIjA5H23I1A+YEQPIC6NolZHqWMnDJEjB4ofpRSLfa0vnzWPGqSAqj+lrLzdMSmC60hPy8
Mr7zZo8PjeT+/kr+VAX58DeTn7pwJMu2i70BIxB/PAw71f8sUq401sszIC06pHvCL2Bht63k0v0p
ynpASmDLBQdfp3dDPydiD1lWIRNbH79PWelJKKsboErN+CsXXdcQgFZU1GkfAVaH6sF2g6zZ+ICw
A0DW2AOaOYXmJCf1n+WC/DV/EhB5iLqLfNH9uK5/aVLftlILzBcH1zP8/8qzRYrdej+1EaGVzRsN
gD0G9yiK2IgJNef0eJJeenB2VwPtZkCmyoU7VEgBupfu/IJ/g0g1Xlr+ez9VNifgTPz3f2Vw/Iz9
st0WGeDfmFBN9VrZ5t/nNIMS77LZuDvWOgpj+yl9qJobXlU2eet2OUFVPT29YedKiDLD+xwnuz/V
+mqJGfWSmO1pcVgGumgvT8e8gsDJI2+FMa3tPJkaVjNJBXMKeg5Xdue2bdqLQw/DiA39AhFv7fmM
R67Q1iRffBPGjxrBdsg981x8vi6horpFioZYEsiCXxSKcKm6tXTQkKEXjzL1P4yl7zIzQLM1LqGg
A56d6N/Kbc/JVU4bx6dr7Uof65Zu8ZwHxt5t7KAGXxNwIuG6QVjcW07IyJmK/5NZzkXHJjND6WHT
ZI3Gk8rWOt9Y3lgIorxgIXlIx4YCQxAIPa+alHPSU7m3elhSFO3uwByTdpn85xGFMy3fRSC0eD3y
sDR9chnYcbBt0InpMa1bWc8kpdQJKa0MFyHzui3wdbmF6N3Rk+uOxjw2DRlLZuvlCeMFVx0CXlwF
scbjylrusWDMOCtcd4u9YCRkH9IMlB3aY1wRmodV6iWuhDut7ej1icRBlRXGXh3jfFdNpTB67ygu
ZDIXHKY4cV43TVVoqZCeYEpdmPKWYGlJqaimBLrOBPXURn3giJqFcSInnFsJrC0cZoZEsRMIjJpe
wXo4SffzMekanjpdi7F18dsu6CCHR41Wnjqq3GIPfUIjCO2/MQyTUzF0SHjv0zf94txpaCOq9L17
sza97j3slTKOi4A0FwekrlRDycWqnYHjk7mNUNLGM6Lh1X2jfmcNn5VIln+BBwdTF3Ris40Q5dNn
gb++RRD0apD2OCsr2nBpqSc4+Gy2bTYK2g6638K6peSh692yyYjzv15TUHRpEQRZuOU5YiJ2oKwv
S92ypDI7RTj4FQQS3f+reBy9DHa1t9+FpQiAl988buvqFkHv8lYYTSpRjDYv2XF5ko3BAH7y2uZE
5jub/E2ELffdkgGrnkBRtPdUd0/ttQ05WDAzGmcHZAzW7tm9xe67UlnVlVRBOonVpyhMEbsj3beH
D9BhnEP8kaL7WuIS+1qwrOJv8fuRgbR8pZosE2hxUvTKsPmYPOhXey6vsdVi2Ovhk3OJRnkas4EH
L8D8pQDIXh84Q9TDpIFKbIHn3fa6Wp5fR1WrgmNrDjyGlbnPF+rzbT6iFmyupoZd8Vf1ycHxcV/H
mNA5V7ZuhjHBY7eUJ+aKMOC9ZPgyIwHDpkkgGrgCijWMAQ59pSQgRf0cI5qPWnBElYjgtQdWZOMR
Jc28QoVaosJcHuDXhmoz+4bB1e1SaB+6zU+5iX7Q4u3QOnUsbsNyVgDnB53eUtIv8tYtnXORt3Y7
qRxnP1qLdUcG3KAWTRgn1EiaTs3/PkQlV0AI3aMGLoW2+ywlEtWjN7s10p1DsT8hckA8wCTwME+9
DS8HPsQxjLJn0WHq86oSr2z27loMET8usA3B2TLJAk3tEmKb7ygAi9KDsFOU9aUjAHWxcJq3+Zt+
xBuOe7CqOvang5ZjVDBKBt4XyiVbvpKv5Qu/MimlXQLxs1b+K248mxK9jh12FqYn7cXO8KmhVJaP
1pVQ5Y9HVqcOL8qgMJYEolOwNGlODlVyWy+uj+eV12IfE65j5u/YwfXtPtGR40yoCe/47NjBmw5P
EE25Y0QFOkgcaY67iPOL9DaEjCUIfO7WDTwdkejQcmUlL/w7DYfEPiWN8ygbJwT2yEEqsJUrhHzH
swGWahUPBPN7iROcKGDq4GTKZSGMSN4S+/j44WtMMW0/pstuM55bsQKyNUdSPAtsaqWpaZ/75Vit
3Z+18V24vhbidOrI2dx9FW98EeiiTLjeQN+btkGidCcvqWOvypiPiT+pjp7Bagf6E4HBctbjlcSL
+M8iP9LlcFkH12NwQfoSRuFY01BbkXlt5uNnRgRlsDzWtZ0pjX3VS1Nm3gshC6clDcf5IbEqGf4g
QRRw47t75FcEmZrRZTp9tleyJ1haNkQHuJ8yE1g5I+H97uhVMuyqC1vbGRahtbczN8UtF84zxa3+
KnciLuMzMPKobzScSefVa8rp6isig3jzTV960uAaYDo1z97wx54C3r3kguyOBhPnEHTHinFk4zST
Wh619unSqT8414K6uflWD3qWA9klhXMkDTgRtQR6eB28EJ3HNePDQfUhuHDmV3hEuZkfp2CEAzsM
7UWlMpfiBohQHxubZkTN5PmeLZLTsaLQbT4RW9tqLHBbN7CPLXIF4vTsD7ECqqr24uZkzzKKUNH7
zUQM794AuHzE+4NXSCRVnsYUnMieSx6m5+D3dKGHcjofJqHuiO/53644g3V+2zExIHJUO1mSnvun
hO0rvHLALUvzhum3k/GqQ5nDj1+2WFA6OC+rasO43XDjHyLTSer7dTUWkx8xAMBQlvxFwdA5jvxI
4id23VE3cDZ6iVm/N8YGiaOxdEQai2V2WaMKZOHjpT6IAiV+KAugBqMe5993KxhIumnDoqC6UDfh
e3pDm5fQvwXRmcrbBMjy37uRsO7fdONAOalwF3cfng3RVxczz8iKlEip9gu0Uk0fRyD5ELCzv/TL
xebGq1MNXKA9E5xYC+7qSl2xLsRgo8Was9BGtZ/kKEsChwnYoUKVeJ1QLo/1zsky8aPhF6wtbtYN
EDfCzS/5f5HBQ2fjXRWhLRgmFZitckcr01AI+TCFMrsS70dQbq3B0XeW4dTGMZaCNeCXUVFHylNP
Q9yWFSkJjxfiuF8PVbQaj0VofBHHsHe6Ed6xVlHsbESdb1s+e8l7S20iqkkWYgfI3uerSXhNkv7F
3QqE8K8mTfaIjmKmbTIGHMJt3NQvR1WitS+YxZLmP5d4zzu6B3QYysm7YB13vwfEbAZQuNw+MZMk
spM/ZQhb6RygD0oQI3tEvmVaLXHIfI8KgEFMPNMpSsQKTXDIMKpziIQueez2bDe12RWTYopIWQHe
m+WTeB/zgA4hTB4MeryExl1bKRXAKog2qJvFLguCAM5XvioMrzdKo8eDAGcftXsBBAm0+4dBlt0P
5iIHyAxattadZfrqw3bhS1RnMJgVCzAbJWra0MbKobd88tFu2jZiD1OERkEmoVFaQtUY/+i73RlJ
PIb6m3F1iIgrXRA9EX0dAOZucFZkYQRTnmgRmdtGV9nUi8SjfDGbpOzpEcKYEuH7D+2/jXBobT3n
xBlzr0GkmKzxZFibdWBTXX1SKDLAPQz1yr1EwLBmC4Dk8kVDZ4s1YMy+/Vc5Rp/CopZ1/PUXHuwk
B166TY1RcHO1L7t7u3qpEMewfjvCFrP2e1xwxlkz6L7ilIo5WmtSZx2XfMaYZdyhzfAs1w2LIye8
NdIx4Arzx9HWbAUwfJgfCzQ8QBpdWa1mZi2GmI6CcJqOkOVw+Z5YAesOjVIi2pBvpOKivqJ+qTO6
14NWZ4UrZMDjPGYOoHvEMlBRAR0uk7kLph4/eiRCkf83NY7zybWLNcrHTECaMPQiWquhWkRG3jq5
q7mYlkTdE/ELtWsrH7MkhC98ybxozPkjBeVGgtS8Xj0dZhsTBchI29JsfH5S+OlBV9mpcBGHtobn
qvfOuE2N299ZEbXHIgqopTRVnv4MaxLj/MAWQCaTxh9FbeiTq+hpxD3VDekgU/tEsiJlA1lhTSIC
poLbT9lXWpxOM8h91cbSnY/S63J4kPBcaV5uco5l5xgYWKeO4HYrdb3zxTMWDsuvl/EUAHcS1kH6
GW/h9VxCxD0rzmhKb4EWfkhmeHkJqtUPyClrnzOWPnmX5gaSSmlO4YfLYVH90SSG8qEJpbsgbTfe
Fzbwby/fAW7naudHzCGEqKsUwrbkbcgsEUFQS39nhpzFGzpRC5tqKIpW3DbELd2mLyj88Zhawhe4
K4vGJGtbnO4tN83ofvHefrc4WQjCyKsi85lSIyC3a+8bhn7mEFH+KiPFfmjchhay3Cz1PuaXfo4U
oRaSeoDMIPnuU6MMAfzYxtMqLzVF5Un/3m6pFCphfgQHBXskcs3PWYGF1yCntUTeQZSw2hHUm8ta
pJMJAjW7SFVUUCJ17xBdZlJLjoZ3YoEvyWZsEDChtq1l1T9AMAjwAY+CjAF36rfRl4GJB3WXmIW8
7278rBZjLOtxAtmCy2y1g/7gtpq+iGIxKhoWr7K88HUf0UUiqMPawF5kOWVoBH8VFWNxVXgzpxbu
fUvnnDBkPJ6t+oko965GCS3ZyfuxU4WEKd9qSwD3S3Aj1aXLwH2e6oXgj9oqrl2uLWSZpaCsXSjc
71A5apc8xbtvY2xW4iz31Em9+HH3GWJTVStOge8pz6oQeMEdHBInJj/zNFo5uLXAIMizh2JlUY/o
is4ra13EQRHAWLl49fs9avPywKJ+0nZTHAh5p3kpL4X5F1DQ3/2GP/PS3XFBFtPtQVNSPn0DOhrL
JeRxr5vywZ6+yOe6L1kBUEFFz+qtjALZoh3nBHCtOfK7Omm5bXgb8C4J/cDSTAjNP2bKHB5//VDh
wtIezYrPxw29orQiFJA8EUmTK8cdNbURyTSfixW7s9VDMVBvyF8FKT4ZwtrZhaW8zt8T41qqRl6J
Q7GSn+JSc8opyC2yO/D8vnQFOzR1cpv3QvPDg+Hv+N38pfxU7yuNhyJEd79HCxTJ/xKuzxI0V60N
GcB2f1tseaw1pPwyFLBglnH51tN4ikhG+doX8LGL1HTtrUmU/2Ar+Sn/XqXMgXrVxCBi+Zl5br9M
Nc1HI3krqSRVB+3P3c96fFiPBxhQ5UjBhX3G1iu3tTAlF10DyteBladLNIKWtMT+1reyONOiqYzn
DeWhQsIhXEpgd3+/g/R+CtUKCFoRAtw9l3rN42Y05oZShzdBSNI7dE8FD1I7SiXk7LL7hrGZ8puf
3H3jEIRPRoci/1Qet2PDvCmCOw7LA4V5HFkpwOvKiMnszxyyZR1XJ6dvxvWIKl4wGa8WdXdkFWJK
7J5XbPUZ+WWTDt0CunlXpzzjA1D5JQGGUTVQRWuHLr1LTEhtoHyTrLjulFRI8q4nWTxa0QaTKmw/
3iDxylmMLY5j5eI49x9/9hN5nS0CXChJs3XKhvWFhwXzfL76i0k6CUjibAmjjl4PvAazq7Z1SKfs
iC/7ByydlQdM+yWx3DyQzZ7c6AOO3saXR0f2sKnbUGF7OsttVVyDMe16NHe382VaeA2dtyusCDkH
o22a0+A+RyisH7m6pKBFoBkKY0bAJQhqochivWriolvL6sN7wYu5P6kV+p2MwoTujttdz44D7LvK
WsaOwjI0T31G7BHWikrTzf+WaIQseviTctqdo3DeLkk0oALxnbdhCg/ImqQcVYJqK0+lN9eS2oOn
rQ0lrDaP3pgrpgm3pSpDqWSlVteHJ9UWPLJH6mlaZadGNgZu/7YsImJMkLpMwGBgrZFiydbOkU/c
mz2MLPQ6ffmaws9PvU2hkmMVseTr1MSgpWJ7SeKIS94o7DYJB0xHSgI002XeLWj3dbOdrJHAFpOh
pDg6DJEd9nKByCqlGlX23YlyuWhMY9Oe40LiVHkuSslLDezPxrPtps1SeaxkDdaAs4+U4X9COepT
/zGwIQB7yHOvKkvUUFesNohm3X3uiA41IfiuY9II6WrZLx5a62NLIde3Z+nqEQw7uEzN8QKdO0zP
pHdPzZ3eACefTxGh/7WRPH47oKqB+4qZUZuxzMBRS1eodxuWM/VWWU8M5r0/0zaX+Rvcz08X/tMK
nMELSONx8aWaHMzGabe2cFGEuZNUo5miy++Z1p4FPlSwJkw/rxL9KepXH6gISLFHhdYMctuUK0z3
oqAaqpJpLPbMRBL6Qh4LQp8j8PpBZ7iAuFFlRgIG+D0AgZVv/17ytbXHgPrgsm+9qdpl9NEpnvSe
GGDlALVKcxFQIpB8WZLo67BKPs0AKHgaBelXr5Cq/ixBxjNYpN/+G0YLw+WPSKyTAo+hBMMccKZR
m8E3vuqGve7TqcFL3lIQjdCttHldlnhNmXNdUO1HCh7oNRgLNAg41adaiFGRF69xZK9Fsy/B6rb2
Va3jdgAOtWp8L38sS63+dPv1lQEVv4mfYtNuSscjz4/JkHh1HSVNlujiwTlVdjM9FYAzp/0r2tqP
pxgMoWZGf4t9Pd4u0CRi83oPSKiLCQLl/vTJtbdrW5Fh3Lwptw1Z7ncIQpbk5sLMZXuwQI8PVQOp
BdXZaWn685OacAFwpIM98/yFwUuBhho+VEKnik78ZHMAh9AzgswS7sxAFlnJRk0HVAjy5/DS55Kc
zMXVS6HF4LsoaWhoObf4HtFE4LFiMlBERvFmEvw88M1FBT+IYqjRHQz0ZF5x1F2lxRM8WAmjVM3L
HIy2aqOl1FAcvw04GTJUG39OLVblMRC8EW99Y3sJhr0mFFp6Mzp5PaQkGvs6EK1u6OFfKU1bMMFK
nwW43+dwN7GTo25YLGJCnRruRWil2QMxRp5p4sEJXjr3ZrzxgM6wg+fGtV2Q6SUt0P+V33bMhlC4
OZciOAGo8VZk4kxcrK9JCECqcoCl0G8je6wbUKwopyS4UzCQwn48OBHYTvchIZPBH3mygxAoBWSz
/5dhMKxrA7AJmAe0H1sY78o/j3SQPZIaUoB3xqUyV6jUO5FuAj3+xF7550s/ZUXD7x54VVmT01Vn
VUzJjSHiFUOEGCVnDwPcrY6mGJmQoB3hMFypAXaFrVfUcs4eyJY3aR4t0WpdLMfQfi88jEWGS7wE
JqEp8yotrFmzoKX+xJ4dE7eGuZ9IlweU7QdZOfpkh1h9KKpXxM6UN6SfyuCSAd5kyDumnvs5mgxh
lLqECwd2clO2ZfA87OL0PNhozeICX64JVlh25GsYNuvih4WCoTkRj+0L19C4LbEHRr1CWhETITES
eAAHVVwmj7r9xo0RxFJyVoH5jRaz3sofSN3iWVuPW18N+dRyzp5GWyEYJeXZzoqrnRBRrNHzfsyt
Okci36a1Lu3K+H96guVnT6akHCBALryVMU2MW0cwDfhNg9470KuPIwVyHe33jTkeKXq4Wqqz9SCJ
Qq0tVOqlk43RosUrCtEvJfP1YwcXoGHixoKRVvxTXkA9ALrLXnvY9C1Ugb3jqAxlqK0hFz6Sw4/D
uDP0fTBSx8jzRn0WO+NTdtkHztftg6v14OXLWazsgavyMmZvzWrzqQD8sGRfoMmDYOSo7fyXUOv5
XUdBuCqQqV+7GsCqVbudT10lb/AIyfpBf3mMSca1uM2VOh4kRgzdUpWDZXryKg8rY6d22k6uTnhH
pUHJLlc8gSGdpl3wDcf+WFwYOEC/7FTUkVe7Zizi1RT7+7hOXR1rN0T+DlkMsDxCwgW0yycpyjgg
ygx6d3p0zJeGJX73hDuwH6aUUnztMzP7VMtdT5HlouzDK9H7tODsPaqKxEhvH6QTfNiWl0J7QLlq
V3Maz/PgaF75UsGsNlXNp3j/caNnNA9s98D4IW8OEtF7V8si0HSETywInWYuazc/n7RvoP3Airp7
rXp75aops2JxDOAuQeVuNtnPszmVFxESH9qHBGzIixRU19mhgIcUJmuXOREm/Sjx3CM15nS5B0/w
XVlN3kS1EyhACIfLLtZ/kN/dvznkjEHpsXnuGQFvbR7bTebqpMozZNO6j8ZdZF9+TnqoswKooBOv
e7dUNfQ65W6Li+j26y1JLmrJL97gdY2q6qeRwFajuiMOVlj1CglulVwyEagPAkMx2BZI20Ag5XMe
1XaBmiPV5/FHUps/ksL0ef8rX+aY/9Qz6Q7E2nqvVFLtGbKFrN9Jauqq525AAVoBFSwWZl35q+t4
PaRZ4YzP2C3l2KFpShE8CNoX+YqRchyZNOgXya6jSY1hF9EYwIkX2cyNU3swXwitiqZIISusqvPS
FAG3oulQCyrlXsamV79FYgKgzQl6OUJiWPuBpVO0/I+b8PMr7koTiMkUs0FkMs4gnwuWBxGE1pVz
bkmXMjBa5WN3nC7gaguB4QBAWAF2N5broslZma2JBA1epZYMStUXJBOyhXP+zzuPMc0KsvjxQFTh
wqBIMFvIyRRZ6C8ERsAlyLn7J93iAZXnDDdhZLo42lKz3G+Ms0cCglx3UgLcMy+pFAoSZDbtrzr7
243ZgjxSqZjQUfNl3QbsNGfeldmHOQnOJW0frd6mySEZK4iyuujyVaH2H3YBve+evHkVQNFPPeE2
rNLcdxTpCa3dgbUMdo+DS/vH5YA1ObtgetPADcJFUE4hazahKVmoyBTVvCe/IgINwGs251jTVEd1
gsiesbh9PZZGcE93g8JaEjLwzyOJgxqJSNIgY6hAW3F+O7yyzqX27XQJ0N+L40Q3GReAaLFsZ21q
USamFoZeXlrA9x7lpZdx4sfVm00pwoApeI8hqT+BBfWqBlEau+OCydWZ6iKl+H/ga8ifTzlD32UQ
lOWHbsPCfz3sJuz5d2sQMAtyuDiq8h2Kb6Oj9ZRfpQCyhSWmnvVtuM+tZ8+hDxfLZAzx2VYCqtQZ
+Dtnh8G+i76vaM/y3GNY16S4GtJqPo6i85PvjTRzfjfRzvd0Sv+96ciGJmaDLUcuua22s6SbOj56
jAI8lIUZpjJXJBIdetWlPYgVpvVPJMSanNS2QbsnxBeTV9q3ncu1ktD2HOlBcXYgaiUe2QGStCAL
XNxoMxhI1bYjg56m6iidMoFT8RxWRiGUijdA5aEsqsmpOldognEvY6cFlpbnRoaFlrY5eKtj8nuT
QpG7I61j6/4jriCzesgJuZ6KtdE5ShKhUTTlVZXUF+Qy6dbKmqfV4D3sem2t12Fn5wim0tRNnUWN
3Xg2Jz/OBSYNXByMsGZqT928YSZHktMeGCeH09fyfMqa15LidVW88FgA7cyPsyW5mT+tHwaPhY9g
a2RlNteBULIDNOac5azxWINs5zpGDfhN9JVweloEn+V1jfBNa8+dXCfJ6RfNEC6W2U8+GGpSYhOj
xOZNg/DL3tPptXnNF6L+ZrNTKdrwmmQtUvJk2VLGhiZlLvmkvDGefXsXW/WgDiT9kwEExayJKPm8
3YgEzYj2xhhOmtKrZZBXOzADez5w7gaBuv8GBqigqu4BrYJ3iHOWaTYrUkciD/4IgTogSZABGW6d
jqZj0Zb/er73OGPcK5orTdhi02rEVEOs/j75lt8F0pgxnS6lHeBSzdtw6O8YecQogKV7biIew/d5
MXb1axxse91eKZL6+oLHDnZj1z4nrHY9aRci+7+3AChi+cDQbquH24S7WIEglggz05mxQiGS3Nv8
k/TkMx75QtMvWuG3vqKtsn+ymA2qTVYGcOuBmjCZHqz9moJyjWQ4ZSCYQi0aQAz5LbxXaMhqWg1T
I4kegMYhWb6EC/dSikoHEz3O/RZLDc+S8gUYb4bhq4NetqANHX+r8dc+ZT5hu8XnmfEzs0c+GDvr
SPWmQ8UXazGn+uPVoFWSXpdRdhIdpuL0IPKj1ARCgjIviB1wsggNzkWbuRty++OY+YwzBB+g0Jd0
NcRcm5HyGNjFCzTDe/H926GlLVSb6l7cqedc7PsSQrE1s2KO0Sr8uiZmYVSmd/b0q8nX+ICoXFJ3
GW5JCn9HoldmdIjYgMRmifsK5uQEN4dETu22nUhepT6LQhmX6WIh1lWLKzBhVoKJzCPqm4xGMv6b
S0aoRpjFFfMQStI7qutQTfwo42TpXJG3uMA0xOM9mX6Opv/pcI7EFx3GZ7pPwGc7r+6jXq7JgL/N
R7JxAwIW70+btRQhIwzcvgE45SV0CxJeIMsItkVusci3CoIOqvnMpB/7ARuyj4mpzbeWWJpxYUK4
tUzLVbXgh8tE1J8A7y5kvxc/EW3qc4/iaZfp8P3HDIFTdXFm1aSVC4k2LesfL9PMv5NkspjQQr+l
vA6CM6BEksw3S8y5GjBM6N/gJ++GTIJXwfo5X5ndYiW7oQAGUN9DIcdtugQu9ZnBqqZLKjpV+tx+
uRpZ5pa43qdoK5daR20gbdAq1a9Iym04O+nILtiuCEEbZrYZ9hyRi/0bJn9mYuMKf3RVPAQMBaPk
xltctPtbcbYmGT+RYLiM9izS0TsKDgxC9Vrkz4B9s/S+nXbATWI3v6rm+iSBpYHWcau6OvA7tUa2
dqQ6mihdAR0G40gtpc66LmyUAGIZCgXWe9+cC62Frf1lfgtpiG+lpHvo4/4iSRHVeCfXPGCBSb4w
o6l01XouNsESGqy4+cJOIfTiP7eewsmsjRspGmLntmNkSc6brF+GZG1gK4v+gfZAuaMny7MUjGYL
+AfA2SFTCc2MUb4iGKn2H5JQZtdkf63RZls2baSrVVRoCNe/L5dNUPEjcjI0zMSRwIZ58cbEe0++
++T0Ja/l+9L7cXW5zcKS2vvDYyZoY/5n0VDbtRKi1glXOi68ZMZhsXkPVMR851aGtqt2uDnYCw6T
69kOrYUVN6A23VmWNQb70SE5vhgfmCBAH4MkdC4kydEYpmjgAK6pM1mFnY++wc1OHWgtx8kBuBAx
82e9mP2eSCASHWzk26WIF7PR13IFibOuovHzAmNKuu1jIF1wWnE0A0ugj0bi+qN32pGHKmiGWQwS
Z4AaTfaaamHc5+mc/Zw9LHDdkN7HXIATQpw8i7H2ShA/JLzkhHvwRchTw6QdfVAeAjvlPV5RxPSx
0ZCp7M2FyqWGLeb5PMp4APbNpZU282nWER9XY+cKT76OX9UktAMJw48plAjXVutf8iZ4AXaxmUrR
vzyBgmP0siYvl1hHstsplUTnD6oO6ORO1O1ZVomRTE9TCVx6OxGiLTKmSCUDtlA2o7pJ5Z0mQEFg
7bGs8GGIuZYh7W3OJZrmNNsl5O6OXZzqDjt7zDFKrL+xYyXoY4T1edPyS+4qMlEgBtOfeVpZDSOR
rdfjbgzOo+c2oqA0dv1DDXBwZ0y2FAP/zfr9TBM9TiuBvql+G9n3JwOSLBsW0nTygV0HVbgd4SuT
R3VowHR7qFhnlC0eQyYaA8KzQ5pW/JegLdllhnVvW6Z5UOfQbaRr9C8KH+PJYw65jK238Nwz7GDO
4c+BfnTSlK7Fw+EqvYK8EUX6mFJUepFCeAKLbCXcqoSq9Ie7QrTEHX8Wl+THMnkSgNktvMX/D6TW
YynmKAm21rZjb+ZakZGX+Mv2wlzU9OshinXgcG2/S8+NWPUthqs/EIdA2Eb4AC9otJukOPtm+1lx
nKi9bWuMlVtpZ6+v/hu8RUf4g2aKeSQpSkkudTl+FGOPdEyBEs6qtHd37+PFFSzkxaVui4b4y6G4
QwwWn/cGqjWRl//Xq2LhzK+rO08o++1hQqL3mFsrfTEVVmd82MZ+TUT7tlU6SSzB6DOlHLO3k3r4
HG2e+o/pMS3zj4GKylg05FBOnWlGrfQDw004cGVOVupTh7+3y7IkwxHGM++tFzAamlZO1E6W6bU3
S75Gpfu3jHb1bN+9iWdQCdQf1+ADMCximw3VS0WrdwuhbIqmSYICFZcl95/7Wp9c3Lf963rW7XLL
OWR49dHG4UxJZogKv5x9vHpW4Q2iKnrZ5tMUI+m9gC2w0p2/6YqJjsyK26O0VPYoHvnG7tkPMB4d
WDwcCYnU9+u5thvzCdTq0BfSgoZtvaR7MFPgm86C3TX1tyEOQ4g72iqHgxwhIEfD/WP3KU9F3L7p
5XEqkcqjWDXQsOmuwtScQfyrQEdJNfFdHrHgk3N9bkBPLWVjIliIpp/HbQHLMzQZ1zFGHsPN5fv5
s1FYUwS0m7P4912cn8KRuAhRrp8YhiYp1BZnKhDWgBJ03AIZsArf/e6ASy0T9aTn2kSdi/gzVPHK
GRtIDwK3FrKGrug2F0Sg0MdlkGVI28xr4Fc9O07vcbTkSkTuOwPqM6PzI7B9dE7U5J78j/OsG8hQ
yNHN7kwJbqUkAWMNNCDAEftWkTajKZL/KQmRNdjoYMbn69j7rIkLrFoIuR+0i91BNz9d7c/e5xNH
C8CPOOoZWZaICFtDP0xqA7zpDXRVWyVcO44XFwijRGKzxFzYYErE17sDr78TmNDf4C80cGOLVyD4
AxFq639dxP6cNU+B+ius6kva3EkF0fx18uXY8uVHINB44aBefKXFqUHArdsqViCGxk7TXR20ddka
A2P9w63kLpcWCzbRs36CZCjKHHwNOs5fESQJHztmzCi3rzm4ODRk7fLzEKel0itQ+36ytfbQrEpI
dSBK5Eij7T5tjkcDiCoRWal8OPC/IwhpABaXyE9HqmwSHH+O8Esog8hSw/R118n8WqS9VNsAVVEi
JQuOxTZTLhDgP0hiF79xwOJ10/MkPYpV8A580E5exZ/CPzO19DvxbqX4b1DtOA8n7q2CyVL91cZt
yG0bAmvKi9Bvpwo5Nz9cpOTmsAN3RY/z7zl7qcHx1y3Gq4Rlg3OwUHAEVrjljSpbk5odTGYTcqOX
stMzBsq9wrk980l4/yNnGN2YD5D9D3WoU39/aSsOPDtBXaG+ohCndClKdiiiN9PV68cUD2e9rLAN
o9QGmD3vfXiFUyoj0KjeLyV8rbZpFBSnuMuTc6YHcA9uqHoit07Q+4tJuErT7EtAEvFf032Fukpo
o2UDGv6Q7cY7YRFwzA+0/PQcIALHKq+0EbEVny1aIFMmIc93UzQav6u36/wJ7JQm2iMeRbmxl2DR
WLOwudU1A2Ak1KEjPZ7voUTRR3Vxv2yNsf6DGaSTu09YyMeGG+GB+5bxuHDg7jMqoTel0PR+OqRY
9fm9MbXi6oAil6zHTjkKxlOlcbrbmgxh/1gWcFnKlgzw+8xGagsVHZxfKvgqcRYfHikOTYbTBCen
Uo0N3PpS2zkRHbhP3ZuqTW+jurOCE4X1zr1hQ3ztr597vY5LU6KJgZjk0kcDvIGid1C22ByEbuQI
F6+pQHkl7mKbc71u/LYVYYpJ9KEhhOC90aFHsrQjL73F6v4gnAxnJJqn0neMKmnnLIPsyW6ePqko
hHKsRvX5nkuQ3sFMPkEy7L97FwFLpH+mcinwX8rzVGOv2s2IJRyumAVg9HdhzX75K4LaKci50z4v
+7sfNTs2j6UGawjAXQ1uC2GzIsuhFUKSqX/aTZA4iaCMfCGvFMmuzRK/Qb65K/C/KCGwMl2Df4hP
QkaQzYNHogpCqRUU1hcfdvIeGGecHc3csQcH7Niy8Gac7SjjM6tTMXzC16IBIqNKIZiGjkT/cGUf
nXFGDBnjnwxyp55XMw/bCvjs9MhXlMbXwnREkWqE5SEI9v5ChY+8iOAAbnviFkNxg884f/12RrSv
dn50/cuvXiiLpyYtkdPF/DMvF4y5FtxdIFopzC19wvxx+vQsZw4o662+/xqHKgtHU+08oLEjA3n+
ntwhlk4W62PFnrTcuoB8kVkiKrAeVk7ZFz6wBEU4rDSB5QpoUtYV5iVNV3PMrJ7t90RTc0zyZeZ7
GokfOv7x/mct2dUT1nLLq4IyfZ1ICqup+zduuB3WPraizSN63ecqwBtoFlExMIiOjFkzqpwdwEW2
CZ9GR/ogQQxWCapgLGqbHwWu0tNpHabzCu6kfV8A7hLxX8IPijbjJpi9+J9yWBRiNyUi40X5FzHr
pYlW8Bmzy0bWrgK/z+ggTk9aRCD/woa08+tMVgHpw7rcN+VA/UAfC2eqLsd1PRK1NtpF01WrB77D
gaZS4Fg4lSLuqu/nmldMNd9Zegm0SAsxm+aXxV+5NRbfbG7RW91etjok2aG2c7kEckYrRhaHUW+e
+hc+7J3LqPtwP5D9hNiAFJnWZcWKjdPV6QdPpfFBhjp/TRsunu776hI6YUCDqDyaAHtFD6vUJhsx
OerSAYEp8CCj7icVO0eaS4S5OLQsBnJmCOgSSnh/cL3NNgJtpZghIDz3OCwoLA+4JXvDIhiLpq1Y
mkXncuzaVd5xIgYUmPXZyGDUr421WyVaiOdNQM4CDFD8WVkFHQY5mZIIH0PpJWDp1H2OP5nx1mnt
wkcR4PPjl7Xy99Kee0crGSVCDvbgRSeVulQIHbW5ld6l0T8xBQ5/AJQjKrPSsFi1VQBMJfkZpiDG
f49XoSOtevjm0UUzyA7MvME7wFkGaLdBp1iespNIrtv36wc4EvBrOXjC1fziL3Lm4w0L6uinKjOO
a5g+/YjauMTXlCUAffPzUAlUfLAXYgntzBDaRuZY9rhOjuUOMbJbgd5P4yR8Wadp/6ETT2uGeBeB
T/lHltixzIlGktamunKXiGk93x4v6+N6P3YE2t0bctQ4o11r2m0kcwroKsujUgMmLIJEf2kqgJ0o
jXJtEyzTxBBymQhDUHTBQls7ZfR4h8DE0uFq7Mz2bOQR/Iolm76j4h7OPTJwNUVXLOx06f57Pkf1
isJEY9aWXzDSG+qNh05MwX6OR+FEVUtBsnJswLlHZZvnXIhx0PH+ONNufmQcf8xNMONdG7/7PxRb
6NNXm8XUlAn07buiAtx+K5dOAVMzNQg2k1iVTDwwF2wQGKF/qni99A4KagdYSjnIhj9EuyJgckDB
oiuudXLrIopqn4ywvsduF27su0DaAJVS5AYBhyfMy9KTOAO/x4Ade00UEXWCk97vWCBb9XWS0XXN
BJl3e6MFP5gsL5gOXD8/5FGCai+celrCp6H4KU4YNXvJxRfnNMa8/RaAVuCHkob/TcGtcNgY9jmx
l2DpG3MwNJk2sSA4NVhKMUEyR2K/t6mfJVLJCg8flU8uwF3Ew0b93eNzXtlgT8/24ncmpFYMfxBR
x2BD7ebcelDominsFsHcYSHUDPtN+YpwvT724Y6KJ/9GXtXfkicUJQ5GjWeMAy4CHZyvCmBCrYkp
Z8Y4j5pnurOvRgabz/mKflHuybfS0XhlIA7waMBrZmEsl2Hh6mQDaBuvJ3WAhPZ4udYnz1QNxP8Z
xpOFX7zBP/lcLLPEk69UTC2pvKOMudK2kstY7tNTnVvMrObB9YALaCOdCscISsaG6bPmn3i4EV/o
d7GiJyGDo/TyF9Ls9D5Q8xRy/ItnvoB7ei51pda02GtlLOAvTa48qRCJYQ1LNCETPxk1ibXBYR1o
zNYFdS/59eYo9Fn3UILzA5J9iLNECl8gOBK1ZNxpmHQ6IWTLnLiN1z/jmN+71JS583S2LR/oMptV
YjSh1YblYGUTFNH/2mZdQDUiHw1q5p0PPazAdcodYQkyb5iovbnVHAXtvxfcQZ1jom4Ipl3mcrsw
JxPPuFcE4cPCin3WD4MUni3rak/k/iTH1Dp3nYMjEjlFnoRsVTKuzkMM+tquZNYYAwRD3yCzNot0
Iez33smQTyT+wi5lhrxeFMZI1ikAlaZqegWUsUwvwUktyHtmoreJS6u+DT3c7K09XmKNdxRqyPZF
y953Gt1Se3p8irBTb+NqRNJIpFkwB3rkF6ZmzPKlrwOskarUcgYVfNJBQ5grEBDa9ZIrHaPXRS/e
XHVah0ZFcW+JluHN3arnGZ67FB0xZv7F96VVLp5+EM19tgTH6+7CFDWYopVb+4GvtIPCpiMHG/7f
EaXX6ADLAyPqPFXKxU/MIrEvfVAGKLRel5D0mDWp4E2RrY+CmAgogkQJS5/wvJfVXA8K6Fiem8G1
NEGjT122DywHMJLY6t27QhOwno9BveE/1OmK5Hh6sRLY3Ffi+8Q7OmooB1xlTIYEtvIStDiv3HQ9
gdSl2cRE5kXLD9I2KXrhAmi3mchlT2mIbiACOjYiNpTc8LcNs4WyBtwAZyopKdQJFgaHOGLy24cI
U4UhBBlRD1lt/uu9QVIticSzOsaZ1DQ6aPBkcefR+q2RqyPGp70x0GnME80kEz8Q2MZc7CBgIYFu
xoqiL7zN73mnZLtKp+8lm5nxVK2AVZT0dVu3HmQDeWsSIFYo1Gss1sJ4Mo4USE90K134YqvzZlmf
fAU6p3BCnh88wnuMM3Hmy1nmhBytL22ZAVYaVGwr/S5etZ0XCkp0xJ99eOYTMmdr3n5ZS5TaZZNB
AbZukwar3DY7e6Q5KuYEoW0WWOmkJIF6Guq81eqAiVfjIOjKorLG/CaazhKhZXYm2lJD5aSQyCtJ
7/ZpIpUxsfKR3cfWnJBcRsQzVLhmCrqqzK/uOOwXU8K62LOM+kqjnFSiV3K/3nWEID7q2gQV714I
OGQVT13PJdMPJENKNgMmc47/D3ZIwH4RArx+bH1Sk58nHhlhgffsmKunm0He0pOn4auFswI+LAi0
p8vIl0P7ebVPgW4BNUz61kl6xwB3CurLKeF2MUvh8aRXdI0t+XfeB8mITt8vMYPCurfDiHoul+w3
eiUZYxD3tu+C1r5S+3mMlcXSRsZ/ZNYhFySh1K5Mprte+C5BkpfOVzZsluP+64vLhQPSJn4QYDnH
mm7Mhk1YwAL+eUnjmgshMaZ6/fyrIMsP4zkgVBbwNMw554mBUwpxp9YxjKu7Rd/fbXQrfBQ5QPsS
fKED686QbwTRkoAxf4yJmAqeYslyMc3HxKF3aVquWgm3CxYlhtKB8NXy4WsrPcf0+Ehp4A6KE2kV
YItEc/wRMEwt1t/5bREbE1FjX0SwykOyUnj2C7VUyDkYN/3i3YPHS0c+yKkdC3UtyfbxIcnEfvod
IEjeJnvqFWNQgyHYT1smTZCxXn2QiB1SXAbPyQV6mcWWosPnRphnQ21nsYyXp9oeuR0RDKArRiYs
ikSxTH8Fnzx7MgGT0PKn4x0VESEAkPsKCP8l+jzuzeg4RyaQk41bA6au2R2BM0hKTL96CptWnL6N
YjIwmWNdtsuZ3Bu3SFmb9X7BOhfTB+LFwNa1jWyhO+ftGeO4SbmcFdDpk4T76gpyS/XT5p/fgrqt
Jkzn63GvmdiF/073bFBPHBaoW/Kl8XuPSTgj1qzgPw1MKDlD3jq2vNCeVaTt+CdFcgsQcXdQ76tm
X2ScMUiY5surLQIqeZWqusUKr8fkCO1SnqQdpAr0lLNAxzBj68GDg1s7RxBbstMj/szv5IqshXB5
P8CUWrJ/GF+l7PthlrNKJnCXyPAVw0Cvnpp+kionOmPf4t/TPWENUhckRSVUeaG0cb74yEo1Hdqv
j0xnZg7PqtBT98gWnbIY/2AG7Gtdv6sSwvEGRo8abPKhK710H3F9e/ZOidpKK6BwZmbg0hCIXS0U
fs5cDqSg7fMU4ZWsNQUOIVtZg0MiI7VdZ6OvJgohxZVER65WKlIYJYqtrxzc1rqH66CJIjHiJBN6
fxBlM5rNQb4aDPqs79hwvYPrFjLHqRTItdfmF3ABBu5bEQrTGUpI/d4QR3Wf5BI2TsitrreugdlD
PuYtvPsG6A9RTYGoMZ1+a2bBNcItrDISGoThtA7lB2l9m7nM3YiW83uJASdN5PFxK1+Cua/L6pCA
wHs/QNAEm/lGy1UDkLOkLt4qW/e/NIfQjJmNsGwYUQGi1ggSJpkGMsyvEjBWGvsHZrkoLWkzFdqD
ksC5vKZ2Pimux7WTPGl4DH+AVWxJcAna4IJg3qp9wZB/jadWN14X3iAylWfjXGwlNN2WsQMikQ50
u5u2VLt1CJVSNj1iw/UUDOz0D0cF7efxPd8xXZuFkXmTk3aTIKOs2XEWpIaZZYtWdlWrMvPp3pUw
E0TEp1c8/hQwIKEBzzW4kXGh058ZIFLILxntra1nqbhLKXd/XvSyvF2tqeaRQ3f0CKa3Qdvp72xd
TOWbfwGKTQ5FJX1zJ+G/OeR5HDisS56IVxeJnUg7XPXZY2H6a3TK9wR4kLXNQBnLKdnQ2p5NfMlU
CM2Pt9D3+f3o31VcDn/aDkgwR72cfnelcXofUGugI9yfOatNi+ny92ytu8DLxnjVywA8Fd1HKT0S
Eypc1s1o/3RV6jFJxXmc5I2XMHtuMumu2uCTmRs6hSiJDnB7FjziwW6B6+ih7WdCj7ck5+/Wp7b9
g4/QdIodpCSy1Jh8wbYepcoT7jOQsyTpM9vsEgAdQ7JDOiLy1+q41ee9ELydU9PbaL8K4KcFdEOm
bIwbyc6W9qzdCBVRkEViRqjfKF5MnwZJbTOyPzXcKwqhThQiwq9ffno6W/i4bGQI0lcxqHsntpiB
Lp8NcrVvNhrqv0AoytpMZZyB6/SguteqZQXqBzuTu3JS3tzoUgUkyBfsj9LpyWgDksGl+LC22Yy/
uk/o7yVEGEGIxrWZtP3PaGZvyZjYxzMHe4pBI06tkiRZvArt1dwbMrYfrjydo30oyPkdnWUMGLHb
4DaNJMJImnDHuGokMrvKVZO6zyTZmhMUJ+0/3hbheanS74UDOQf4lUx0N4EEAYtn4EnMp+ug27/T
TauUeS1dLj9RqsuMkVy24D5s8NcmhrAt/zWjfEP0jbIoh7EppvUoweJakdKeDtyUqSgAJalnxuzR
gQ5z/4dur/gwYQxNuD4Q4gA4IxOypZ7J32q2VWiLysRakE9UFzImrT8bAjHkoyBipaHqWn4LYiLQ
bv88POvwYpEWm2jBsQreFAvoVmV3F4qBabuJpmGc/4QEGztatHxn65HR/OJOWn0rYda9gT2cN+iB
uAdzf2EuUeP/1g73k+podaXcaPR3Iy+/tlMLbjMpFJM1Bq9mImXSilFeOiBeoDKH9QDVeycp/1vi
Xr7ppYx8TBBV3s3MMS4Jbw/u3MjP5Em21pde9HASiTRmCsoa0faw2Hs0k6ZjestPduAfmwxTOhjh
FZrVQP7jJo9WeW949IV5PVlcHAekNpR3NSto4j8tuCU3/RYXTp7Vq7h+9vjShuJDbrlayZnKrpqo
GzDVMl7RYAKP0qWlnIutzIdDUPWtyR+A3DiqY9p8r0HXAq++fCXdoGLFobbFadjskI1qENKGbsFt
+rUlNcvg1OgcjPd3+LFweK33hRMTlDFRXJgG56gqlZ5979hgNgISJ5MoQwNFgBl3e8je0h5HsHXe
jNdIy/Oe8nSoFOnbNeN0LLGhwRZTY4JhR9K3ujmPUJhMRt7znLv7FXWjyyyv7HXV+tX07KqIteO+
XQhNjMlLnipm3RxgFeB1CcjgNl+gxrV8ldhrlWa0lMt4Xp60aYRAUOuAS+sMReE1XYJRm5I1xMuL
0Rp+5udMuYl07De4o0SUbKHCxV5zmdYf/DVhSAOyQd44HiHwKqmXv+MwGh1FYY15KTiPriqzNuga
INOSMDlOtHFgIl0oSJirSPFvfxzHfLf8GyXZkg4URFrQNHV+r42jGCNyHUQSUlGZk/r6BeaQkKMk
GlC8AAW1zjpydG65p7dzmMr3bg+J2vW2ekr5/5mOXmmtJ4alXhvE0fKm68rHFzJ8rH/DqXcg1N+d
RBob1Dbg3TpIpXjBdcp00g33a8TjveeFmQD1ZaEmx5Sc5Yen6hZOgIriRzUjfuHyxgD82Hj7GymQ
dFu/mtb8XO4l603EzN14+Qo3+MAhS4CgC5rN09rq72KwKjZIqTUl+uVPcgG12izOSYs3SncCf2Ki
wMIdom/CjnQxY1nCHTR25H4pzpxSs7OgDrnLci14FfieizOsAX/b8mRkc/j/XP1LxgRnCRNhH9yM
8Vy1w65myzy/q9hDcFEaJTc9ODsvSoWU6x49noNboapQDOeSv18JiNLmEdzjDqqc/Wl+iv4vvzN2
OpvQSvS6lKKcB3fXxQX4EJ2ZaP+rpJV4mavRPXhGApqvJd2Ro9Hn5F1z2m3/Os/hhKaqSZCG+tLQ
mJHijIcfkz8Q7ItwVfESnsHO7mO/iqa2lMphL+yGhtQIDLUv2CocRS8w7NHXvepRZoGdb4TSfzQo
nFNu58dmCwZV03eYQDQlNgrI7DU0BaePLSuHuUgUBI2NpCkMlLUV6cTx7CXOQWIGYQ1E03k+UXh7
d83ugs74XoUhhi1nFRl0/fV/E3bsvqSspFJiPzFVs0hMkne4FJiGtRZkC0cnl3MB1g+HJLxMZh2a
ESCCZ9BMPlxnq0AgkM375+6fX3yvrm/ntRuOtPRDJxik6FYNhAhVp6/9q8l1uv0ASxgejY3vi2XH
l1bMCSB3U8BMP0k92+ZuqonrvL9D5sdgOyQq07lJtWxb9kJ9V0icFAayKOIcXfoIJDsNLgrnEYxZ
d5MGVQFfN+uR62qfj6wSDNUAIuo0NraJne2+D+6ahF3BO2HXvM7AFHcgDmpXTFLIISHLZTSAwKRd
h5YeyvDTdqNyFznBHM/0K837LCSsNJutt1+TCey4A6Z2V+UeiscS53UF6mgR9WxO7ntqnaBdLVKc
9TEvxy2fjgAsh4eqnxTfkjXUydN+/G+6HMOrsn/wIGYBFGE8RqvL8rn7d5aREfQE0j+im+lB0AZY
TG9LVXgzsMAIGG25Hzva+JRVomt7SoYbcoVVZVmJiiC0nrALycEv3Lxo9Me0f+QMwIOXC0izRrFe
T5Vfl2+qSZ4VvHNlYjCzAsIDn8cgJWwqy8roTgfW9VNeNF8sm9PATXXail824HV+11Ae5ltw/FxX
S3XxprTMSEdP0280RZm3B5st7KjhoTiSe2zQW4ZkoBX2BSwzh5IpF8W9u/a4x7FStw6A7DrT8I7e
3BWkyY619lQUBW9slJT41mc/1gKM0p7vRaXKgSPBDQ1ahsHZU+rrwEnT3ZMBicR+atus464adFyQ
i9ysz/hZbyzQKaRzDnkf2W/tO17gNp+zBOeHdVMchBHfFSmSO64IfIArS4qXNC0tKGtC05hud8Uo
zPNpw3JITHOVgsz78TypI/icIxMCQTSjfKqbrXzwktECr619WJrPwEVNgBQpwVALORs6H+umwn9D
X9mFpH1UzKIG1DV1D69CeAzpxsNNad73i37ameHk/RYdjEDwTMX+9tbhxsYH9C2AprE9bs0r67vt
8YjnizeY/ttO39tPR9GqlS+lzGon2HoLbeHjPzk+Dqghrd0Yv11/iJTUVUaSVs5adeauoJfZZJ4Y
maObNaCZwL0KGrPiuv4ZVk7zyPHMHEUHp6dlB5zQsLA1A4DjMCUigXWO/qwUqjk5aghgDe3+TuGv
cRXi3gPmBIYenG84X9oEAtzz9CQpenBsl9TWKcZ7Lb2HHM8n13UfxXr9+KkLUydFyPMb31EvO9H2
TOOtAh1HhRtBnSMRhYHV+ZUhcTzeBMoEabGVEf6LkeGAAFja0nG4MfEE3QUyrL/pH/DqNOx1iNM8
HNuFjHMUuk7LmPJDLSG4ywEmq8DRqQIXOXOuNJSgZXmMAxen04hHyA7D2PU9Qc+4TOeXpfxgJJ4L
gXfZZBRObepJn70+LPbXl8vLoS+oYMDZPqdznpiXKcfUOt6rLLF4MOZxaUMSmOgpkDRl7bAmP/Sl
v7GybalsoEd8C5NVinRsA3OaTHDuUQiOmvJhJfKllU49ri1GhFX2BAQCtGwJaNnmIoOXUTCskPHF
lNywl9Obk5UnDY+vNVgMUOKlC1T7/INUubpi16RJIxAgz8fUYcvHqjzoVJ8f9ZeiOCN52SNjoFOJ
WdRL7Q22ypk5i9Xq6sW4kfMPXHtxLZNqusjAHXGvqsDiZRg+Oa5K4rkKMvtBc7NG4Qso5ZQAAEj5
jcp1lzA5RVhgXTzFD0WagXm4acToEcFFc0vlm+ENPn2G3EctInHvZJxy2ydGhXvDg+aDbZOwW+hb
A9x4lIEIESC/0gr4xMF942etNlxDMJQt3+3FZl0bErKi9QauhVXbET0usjReZAN/BU3Y9YMgfRqV
/1Sw/ymi2JjRWL2ElZc197NxYXRdTVYdpAY8SOOMKnKYZJtt/fT+1Gze8Vei1g6jrSHjtRSdakxt
s7oQYsibl2mq+5SJ4e2w3H/Mfa8jth5kjtylMMmBWCcpIRygrNOHAYEO6RsoEwP6HzFEQPflOi3/
ziiweb6C0plnp0nl0fNUDGpIGVTQI7emvLUw/bFq9r/fXcJLRq4GQ1O20gH13xhWxqu4Rkhg4c4O
IAw/UHnHcN2+0YWsD0u1eKK/2crrB5Fg7sb4DMpzmsmbd+zJCi/8OUO8ghr5bbhMyQ5mtdhHaZjn
jT7OZumhfXfNYiU0onBDtxi5kK+k9XKfCX4PuZEbsxlgKE+dyiN0PtcdGaJnxOiLd4/YYzLam1Z2
PzMaWBNBkvOn8ACD9gZzBv64fn01tE3wnwjZ1YIEuHNcR2ReTf2jcODFndjRsYJLIhqNxV9DNNd7
Sok56n6FX6yzkee7PH0linZr1Y2BCjU64TfCV19U+Nab+F5IB1Q2VC7SqyrcSYYMyV6NCemPz8ST
c38+JwAU3fol25Q3vfgqvMRfqvds/5LMduJk/2i4YXXBu1hR5pkUYQnNGtEF8d04JabpwTq5LDvj
RAyUpvXxeHyyvU3FHuTRmJlh7rrZUfsilkTqhy5vIoLYkEyJnt9j6Xa9wfo6QepPzYh4IX0nHPnR
8cPXirxKPtz8emjfRj8Bz2CB+79QjoBVRL42gM1YAWyntMo9HFPnJYXrldvPdOOSWKafUOrvmQ92
1r9L8SzRalfW+l+tEYf+GSJhnuWL145gupXFHqMpG/4mViExzhXkTdgon0HTleAfh7iCj8MhVUD3
GET22UZXC5xoZtcLdPcCHa/XgnTLfDp9DOhmg9XmAfqq/9vEc9gWSe5dUBhERYaobN3HsVwiOnWr
GqqG73HijFLOtGLLQ3xOgxhM6eLb/wCh5stWpOwXrfFn3YXILQZwjq0RDFPMMKTE26wkuxSIdtJy
bNWASAbZRz/3bbRkiz45zx6muFPbHz32vHSyv0qrTIVrazFoPipSEKGPEaJ6r1l9/mJrHy6uSwLQ
2WWHTZGXL+y+4Hn2MS/ddEONrICxEX2YpCJDKuNfWVdxkvfm4u4An2hU6A9OFIVHILM1d0x9k6ve
d7kRkPpeRixbQSCjcVChSwBrNw851QiemVbnakImHmEkLh2zo7Q1Oe+PKXJvFzLSrLyiylVvqE6y
sI/cyLWHCEAmAtxwAonVqwathTKkNxrns9tjLyImgp73wbochh+TC8tOIVdpk8k/4fAApdInSZvw
wLGzOck0LnPzt2buHiKyCM1dVe5ww/n6sVzVfF625E3nw+CrxtfX8FVBnuhSLRiJRLT6jRJXuuF3
tM4KMncu8r+DnxCA7rXu61veG59o1mcVX4X2WX+sjRGDGBs7IW2lyP6LlIPV34j1/tQQx7pRStZG
Rvnn1ukKV0cs0oR7AJfOI2ejadU6LyNqxjPNdgpz48aq/3Bb3DeGPRTIQvCv9uYDEjFGlXIMH/yy
1bJ3vTBgMjhQqk6emBzbliJQYS5Q1Qi+d/Qas1Mw0zDxyOIoRa0spmWESyjzFuSdVlOnLiLSzfru
0Nkqc5lpjtgxjlxkpQeMzC4GfJlE3SWoXTNe1bgaSgcedjw55ByBtqkOzpaprFb+L4E7zdb8Leri
LOqLmwbJYY7FWkxUA1RL9JFAcsOLh8MMWtPa2LfFK+ysSLgU8UikGhUUrzSFy6JkI/staN6DQrq+
Q1HqHYHz/36ihmiIzFstwbeestbDKfxq5fOoshuyjB3+aVx1LirSx6EIukwYQEoxeC1H3MJJvaDv
D1TMPqEgEMrxqN+k5/VCudIgkJH+uCSdjM996X4jsuNX8VK1m+RKLtIbBKl6etufIEvbRSxrSpID
UluPQKWUj+9HD6v7rCk/UOUao7Zrbhbvu0ihdNUOvq4Ip0qEhk6+DX4WL9BGCdtexZeJt2ekaA7R
AZKCbY/1SFe//tIbPtZII6zJ9qDigdtY4qMM7Y/b1O6CyBUFfDuZ9OY2RuuvkREz7Bgo6bSQlPfD
8H2lNmoixYjkxKGIkq0Qih3gvGKH3uYkSG2fmmcRP1CykBwEgzbgzuBYx2xUL+XDKMZwmP8X8SMy
ytJJT38FpATfQon8bhY1WR6pLSANBXlcJVTJWVkpLou/o8Sz9erCe36TQ22m7scS1xCmHpESOACx
5F+ffOr6xK+CtUqVIju2GDwwUGRn276qwmpixVmLkQGKQaL/0QXHnxKk3ITt+SSwpKtgE0XaBi9F
4QJ1ZT96xUKAu/UlveCRKjA7nNUiOda9bbDTi3NJiqoGajo3jItaLYLYUCaitByehEZQqr2Nz6Uh
tA1NPoh9rkUf4kLNdSemVcQaPOquPwgkNGyIC1P0gszSijkauUkhl2VCaVNdCG1jB5TtrqDiRXLS
9KuuuA4v82KEgFw6TXOda36ZpxGZd1PgCfoUeiuWIQuLgkMniPRldyri4iMoC80OJBC42AV4tI+b
82b2yQhjUEV73NC/awyw+A9PXSHNfgkLAzA8sJnbh+tO/+ftdDXsSBiHLyCBWOdPIQFkOA/g8UAM
Lh7lG2kkquOubKMp5Cp9HwK6ZmbK5mFslKpQZkcOEz8xLBOXoHoHSc+cfPgebqgUD5WCJIUZjzZ4
RX1AycFD1ho//MDBy+slTEDyPs9stDkkgV64zoEDFNoyO87Z/BSG13ojCoeDGFxqTw89evnqiX5l
Ifs2EzdYYMHVMgIAVEJqU4B3Z4DHwA3n8XdPTvUYJyMLIizbf4l0D7+3ylU0wsnIP7zbqjojnLW5
GS1yTSqYNJ6ZMPsAcvDmEoXF2050EKEN+pLY9K2sF3r2ORj1fVOAn9Iz0bAC2s3NM0C2fyyBHLbs
rJKO923yQiiIsnyb6T8NODcBC/GuJ0H9Ewme2O2Utm53DFRIRa8gXQTxCJGsiAEKl+wDyT2G62TN
TgsIbFykDnFUb5ba/pYTDMIfT4U4ng1aLFYHSeuOvcI/uPVlZaWfcEfToStSsHLMBlpjNM3NSqby
RdhKNU/cagPHSOp462xGPHZM/QZojuY9s0nRJDAM+CIZ/db+ope5KJOytBkUJiRSChEV3A962Jmw
szwdyeNnKVu8jpGVtSl+xBC77DhLAV2ZVwU/TT93K+X13KsIPa2xSApg/y7Jo+/IqwPHTTBrM4ff
mjrGi3IMKEWcLd2GPMTDhNhdE/bOS0yCNM580Le/l5vN4PW6Mh2Ewwspb9cZvcdJHyZkKAzGLJYO
+bb8/W1V3R5cLODGVh9mb8hMVjgCz5/h5/Mc+o1PePAQCwFuClZZbbuDcogf89Ctki4p41X4sW4j
sh1WPqNm527kUIAuVnZ38OyQhyJS9zdSCuBT9jpk13VT044vuGep3Zpy2NQneKI9kp4LTbaWupkY
cKxetVoWlMpCSPvHaqQ5fNYOSk6MgtbPodW4WqKqcpaeYg79fK8mkBlqXDoR9YlhJstCq/Y4P+Pa
wiXChogmO8/fsb45V58X7qEQvFXRSkMqxGlYMpSnRHfJBMBBE20xgaXUOsKuEy1uroBzDp1ZUi3D
FCdCMMEqP29J7IlUp6eLuu8kdC0Al1sVvjjZt5EeUfxgtnr6ZEG55EtvkzWGw3T6cPlNLrumbiYX
i8+rloW9Z5XNVLbcazYlBi3a9y8oO7KVVSpJBc1wH89rso2LoqtsHySVmzOd8f52ZzI2icuMXI/d
76Z4/2eDRb3I6k2bTWg2QiFvkMUn6BOfVUAU4fDczxbswqStZvuLcVWWsfElgPbi+7mhrzZMb5ar
PQLzCX8uT+gKH9GcM4dvC+Qc9hyAoWla1917qXqVfaKb4vMT64uPiQnJ+GLE4KN8zDOhQQInmtWV
stmiLWD/L0uyj9P6RfIdodPLI1rCLmQbYb5xPPlRXo4cB6xVSvc7uaVgdl/sAlTQl3nz2WgAe8E5
lcUNMU3s4IRKlirZQgJtsLSPrZgRHkb+f1q+HXkWl05nYLHaqe1IjjZXIqT6pkLTpCWgwvH1Z5gM
U3dIMtLu8ygeR6uSAyIytDkz2IZrN/T4SspyvKCb8nuYRpegq1a5QlAx3MgV+KHF5Of72JZKAcX3
IdaOOmHAIpO+NHg7ofaRi/A22/SJ49r+UC69lk8jrlnqK9mMLhqVFwnv5MLFxWua1FPuo07+ET4l
buo8cMJjjG+j9w+ZNXL74yG353+xS96k0ih+8d29X2XEAcbQtCvD+cCg58kiapXk0MgCMCkMmHfS
tk9z5+ycrfEXDZJBr4wdRiGNrIIIbmoq+6J+0lcb20PqHoPzw+efoah/mxkqKNJ5nBuHZu1gN2Pm
JIW/8i9yzf+63SsgA8Foe+dr+rR+D8b+NA8pBYJI078FiLbg3aviuwga0w6t3lPlq5xVi6URINZ7
SXiivLpwb1XAe9pnPmiz+xTLlEL+gxG06a983Da0IZiW9XudAzxxQNEDYcBWC2RgfheODR6LNscl
yg3KbZTYqnO8nreTtggJnyCbMfTSQjTRCViEYadX33kFhkH5oPq2WsSYnEFSAbHbSKXDAut0dGrk
81mE0a47mX5YJz7OcKTFuOFWk/4P6FIQVMgTgCtCvQED2DsO7LK740BFoCi2jWXFMX9nx4Wn5saH
K8GoTIwv+CZ1Gbi3QVYd1SiG2daEXzndvB0gGPrVPl7oqqfoeneBDFHzeFD9+Z7Uxp2F0B/d6JWq
DXnQtmwFFVWN3IRUbcKV5f0jnTJuB0ARBBoO4RSSdwODv8zniVsiOVeSzLEq99SuNV0QoA2J4Xve
RWsEs3iyaOO96tST4d6qOCDtDI+KOVUkA+w9nXw+bn1twNMhK2UX2yZPTUIaVdg9fL6Z9GSSZQHU
17la9bzLWKQmq6qpOMUjGZEJmbI/9OhEawC//y7TGfPubjUmo7r4bJimyi07euWI3tFXKJvPihyx
X60TzLGflpiv522DTdFYxLMOJCogZd2nWsqBr6ThvmC2LTF2q9RtGw3s1gZAHE/3YriPIk+ROZmI
Iq1t6DDNgTsqDALHfupefPvwujy2R9Xj446fo0FUK6OnVZdyFJP5iYTSgtLXMWB4o7GE2hylDrm9
LKv9zD/RImRqOYY+T+2WvFpF3q6cc6YzF40byfS9zdalCWQAOQhAGQzjNWop8JM7rsTSZWqBWGuu
QGe9mCLlITdp8YUqXj9Df5Jj2wsV10a7DDAA61dwaHqPNciKHn2fyXTAbrvazB2JosBPrtLvYEmx
ouSpN4SAByVgkCNWzzBn868Wo6EzyHz18TEj00XPj2YoCOoABNRsH57c/hLYW/AtiW0vBcdpxlbl
8aWwfZA9jCCDaK0Gf5ouocOUtNfFsLeT8sJU63ff5d0h41hK7jWlGgclD6uieKxMucbDm7q8AWP4
cUOL40seKq2uMs4XT11SZQEuVjAP24zM6dZjfAudgv7NEKnU+DVfvWGjL+vPNzW4oIyL71IhzcPi
uMlWCMvih44dKeM5IaZTFMokFi0jo1C66oEvNWxew11M1Fo3AHc+ntHXg24wDTJ/cCRkbyv2dzVa
PCYjCNmfqAx/Ev0k3xBPdxVoZFz0Mjph1WBx9x58Gotwb4h2ilkukAxgXqgF0QjaslEgcu+HD9Wn
TvF3P6stG/PKub1H7j2pzXh/IjtVIxCbzOucNg/i2wahZW0JWgfwlOxW4tXAsR/c5aCawgbIiSn6
eQchGM+gTJkUrhRrEPJqL+ltquFPIUyWvwqirZUd2CJXf9p0ggxq0yR7Bv7mlXM7pPwOctHvZLEK
EJoqdvnkHma1qnKdZc1L8uRN24/bYHfanIN2gswHMgELv9Tr3ZdN23vIqNN66S4TLc6HH/o7IqqK
M+gPdmsgtKpCxKuHtFISIyLhzyKASFYFh72cwnCIra2Qd7eBoWnin1TkyXTULEoICZZ+OyaLKwfQ
4BjBWY7l+Vj3OimGMrzjA0S7YVO1QYNfq5z6xwI8ePt9oIjK4a2HTde8lkK8Cm2Svsc6kQ3mmJel
oM5JWuq8oqkMdp77NP9DiJHFQGIC/JNvpSX3ZsIVN3LYlSESn8zmSYjRJwQqIXcmnDeDbTcB4WD1
BGa8kCyc+MVn8IF1ynX831wWyn4bTteVe/EmiYWo7FOTudGDVU61tNEnvN94ozcPJU8+ah3b+LLS
rRubLmuPjKvMPTcogfcCCu2zlDUl7wls175H4C1O+xxq10DMa2hFKhdMlbANaSAADCMOEa+3z624
N17eJrjUvDLKTiKSAQD6Zye3JFdQlkvDp5Ak+r/uPD0tsb2P4VQ7PKEXJ3J5vZhSOuBf2mQI/lNG
3O2aZVHhU8ooQn35nLpVaIITlokBUGUz7d3Pqw5nlJrLGHq60UcCrakwwmH0GH52e2Rc5eJbuWhM
HUws6vc4r+OinrZgRVSadp9lqtrGjyT6qFGysxAESYYE+00R4uDYst5+arA6idy4r3TkvM+OtUbq
9VwzA8xAOuvk5gZUsakHHXW9tnAPFV1Ijy4C25ye4FKEQ6G4gZbL/N3zDPeydcaFZhLb4XyLsiQb
d7GOFAF8QSjsXm8MFIIC+T7Y+axgEpzBJaSPzoo7jKB32ifXN3txK/UCkc6NmeqSkNZfA/kEr6SH
EyST8R8mLFAL+j7jbS88DogYAAXKqnr10uOE9SIhO9ikyz5GtGMIYiDjkvTcDcMvzBDGUey8i8ma
rDxO+iCE33AqGZpi5VPXnlBe66YUn+eFE/k1C6ViFspOHCtfFTLIafpcFiLusD12pLfhmVvlPy9i
VKCBbBV81+zRWw3WjWLWl9RS8T44+7CdzkkCgLv4zj3hewE0klNgnlVcd9+QT7dVBFdmMorbjHXK
ige10gA+FAqyVW+f5sJdt3EC+Jn1vmtliH1P0ghE5FE+GlEFrpalmM+5LoXT6Np29c2iwV3Sb3Xk
/EsM+RMnq9YwAuKb7WQNudbg2waRdt+eqF98IKm9qUCuME6QxESPJg6j6lTr3OSAFTlXNZoCRyjm
Jg1EryoHS2y9egbtlupoEh4n3fLKBeUZoAyeRRJ2MHzgpK0vBVUKqXX9JsOJkbdz8DZGLd6toAd+
zlGA6KQX1dfeRxcOdQSwU4m/SuUrWIxTQeiJXCDK1CtVNHMLmW4EEBp1PPOAF8yFLiAUoyzjp8u3
+DaSrhsEFLnl/ls3t1mOBZfTkR5oziZIiK06MNQlzTfSl5DrUwNQstzD/IFrC+jeuw9eSlxx22jN
I/P+yHr2WaRt7QZkv7zAQU+Lbs7faNJrECR6N/aZkFzWTCy4GqJYvYopH9UNxqSGAeggM0VTzJc3
qx/5CdV/16T+clnvuqaVpmWNuMtDY3rkNjbzdgKrO5G8RC5f9tcxc+eY+lSEopSMnIjWQcQXdLR8
uo3F6ZJHYZ9MlAFehjIXSNIl7I1Btomgr8W5o+uHWs+TjzJmlMx474WcC9ZFMf5356SrbDQ9pBQ5
KZAFwKNocX7B7yW/BEm6QTLFZUw3c0er1iaFSzhz9ln+Xtj32GwOk6BcMn25rAnDOa3Ys0kxtkH/
vXBZN3a3ZQxKrHOrrMnPBbFhv40ltKA0BVDkWl/wzr55kQwHoDM1jWt157xn6tnmhLTZhVXHjjAS
GvUw1x30lHEh2iYn5VNxia8uaNeAxC9sXe5NSf+gH3AXegimBUwTcOc82o5qKvTFJ94btbgXZfvp
LyVUTEC8xmqdtBgVhUUkXor/gK7UB66qCf9UoHXTWGzzhGGlxfj2fEWTi7LfP9nHdF+bLZYIAoba
xPseNlVlYVt+O+EFmNj3vtelzCEAFE7OSMOcx+d+KWGddneE8SzzmVCmoGezOjuV8YlXUa2zW6hT
rY5/+p3WTAAFIeqS8X1opDgdcDNfJ6uJl8OLopba8zear87ZN7pgw8eNB/wg274c0D2sT4NXQdPN
Gf6av+Jm+U7xQOOG/iYD+5o+1edjU+9UindwUNrXUhS2tDIg2iNRgrGbidw5dnZnhL7ajVn/ymkU
KSx8K6oUv0t3KaE2bvkTB8mW0O71uyc61vPzqbRl0S5AiMSSxpYXK/pllQuqaNxi+v0x0AvJrr3s
GD82PEgjblLalQmTdY9wjiCYbj00RVgsyXgU5yxNtijiIF6VX+3MGpqiWLzZlIhlCvJS/yhTHLjv
nrgsfubrjxfvob1yrzoVs7GetH6iD9WFaZsZMxcq2wdHuvThWkLEomP78OfOqD5fJyyAC5yg/es2
PcBdRAMIw2fRHK9TuM/LSdmG49jUEIQgL5XVLNn9q7dnbtKxQqp6k/pmEweZTZ5wYr3NMObQU8Zy
jxbwW0AgxVjlK5vm/U0pdWc9KweRZWGbHl958xLmCvQLmWpNJpuL3kDDyUustZdapR+bGJRaaMZZ
sS/kSJjvS/ORdINMhjl0zD1Q1+S4eUJcaJrtp26NXZnNeT+v5gB1BUaeAmTawLkAkuEiHWYJsgfc
M4ndIyYR3Irs/EH7f0/YpPKZ3gQbrxkdePRh8u4Ea1zvb1Grn0dFJesdGxEQCa+37IL1E5cYpPBC
CA8YklVkIZaEwU3xt/CxQd7BZ0VqGL+uDOyORjks0LhQRTEgga7/63yiwHKbjF9gOQMXQaodq3+j
1M/Z7LLWGgkAOfGj2utJou02bmE/bJ1TImrtcYOeYivAOHRKUp5fMGwOKQNRtcBape5zjHrrWM1g
oblLKKFNceDd5RxDMrHcA2mNHMfto+tHrYPsbQRS6DHwhAEndR0bTGtoRm5/W3CooLVj9zsHD2Ya
7/m12ltnW4AvSmAySP0KnsKiaP1Fty9qSyfiPVtLe2xF3Z5ksx+IGyBKpcaD9/4wcnEGdoiYoPU+
buKiL6R78K0Pzr3fqDY8Vx/FpF/MK81MeGT9KMzSPu/2+dQuoxxTl/8u4EtjOow5RWM0/D/AvMfN
VdHRrtgMwQPuMtnMB84+MkBJBQ5Ohr18+Kl7/uaUBMuzi/Q0EjoHGnM6HOaUs4uu+fEBm8oT0c/m
FLUwDjziVmASY9mKnQmJ2nhyjDGTrsLzd+ehzUFBLbQoWhP9gNUqlnzonHfeC7RMSGJ28VaAw75q
tgS/pRg0IPL/YN/KSuE/p1axRHAjuRaC0pwBYsS+Vw4dnyG/YCOhzlhNX9vTpaCKFvgBpPhJEGcF
odkxZlrrdTk9PyqaCrmk+jEd3RjAPSN5hOfTl8BWCx2HMwuFko83hH96b0h+Kgcarwc2y8fS9/FU
xRxoLbs7IY7fOBwUvpBaaGLfvHC+TSGyhjOWFxPjMFvBYF7PppSmj08lO2H5sn+Ze+R/N65/3YhG
ctC3Enhn8JCpQHbqHkr2zRZRzy0p+sADOBB34TVofZ24YAZ5clHYoy0/cPFQOHrVfRHqPTky9ddi
KC7AQMhS9iNu2HmiXWwnO1LKc4FDGS7llkyYvtVD09+clPwxcKqTr/QHqvkS4htnfdE4PIXnbK1o
NhIZDDnjOSIS0EX02N9ouVn6Km5PTRNZLqkTBY/lX6C2GD88+Ex9TxkS7YCExcgnBS3hdFJL807M
WpMMytgbxXctOabYCP1kzG5Fy9jvr/qb+szIz/U/sUPJ58Nrd7/c0L65jSWS9TkP9o39O0hYvEDP
P50QO7HX9LRjgDyvNr65/eOBu+SN0qHjXc4gJzMhENLi24BttZGyQbfkhkav7auyVKJThy+8O9NL
W71VtR1QgeQFQcUYM8QQs4nOPCzl01ou7WoodLTwVqd2zDjcMuYfEepJ21nr84IodZF1eRWJNsca
+hIoysZJ8TxK/5snB7oYCG3BJ2DA21oUsuYq2G0fUefeHZrZ5FEihNjQ+SBQRbE9sF9UG2myds8W
Zh10tc5ev2v1Jcl5GSyM7x05S+hKEVZmfJREZ9pcjjkXXWQRgiihs3LWqwa+38S3vlTJO3cmAFVk
NHco1GDxKoy4rfasr9wclxI11LRzgjYIltIed82GS6wgI0YUH7HJoNABdyJOAxuy9814UVnEUmv1
pPyhhVUyC3u9ORpls8ComnhXzvARAXAIJTyItbU+pZyoit+N+cihP1cHt0oxUsvOYe87ueBZXyKv
2Wi/+3JgjJktWCAMHoV0IefqriZveg8M5LBgVnvZ0LafIDq4en91hoaiGmjCWp2ooQkN8U3ZNWRD
mkj5VetV6CUbbzQFgrFMnqKcb9TTfdamOKJrcyKrAeA5cRv4OA+2v8qerZ2+xt7SW1kL8tCPy2wt
A6Amcu/KCGv5eV63O92QCfAX3YA9f0I9vY1pMvmnUFaqS4MZuEKdL08/+Z/+a83DLIRMItfqPBvd
jzWwS3rBe3IX3BG9wZ/HCHcbJZhryVv0ggYjWdm7+tH0U537Zwhj/0CQW0MjsRWyC46wmM0Z3Iog
qwddT1LRn6b1NrPSSyAmkHqK4RlpCTPBH8vyAT/Ke4RqO5PeFKkY5tBYNzjdBYTHbumavlje74OU
w+Y54q3txW892c+MP9w2MBMiaP6HanXxjWxv6Qp3CU1HoW/rztT4Ssfsf2RfScmRs/QFujzSJh57
kgXGuIA6pg1xyv3DcaDFQvaIfqAuiIQKP2FZBWsZfZ01SiPWu4pdbN/gF5mFzpi/FsY2uz3jQbKc
laHzGhez/S8/ZQaCPwAxK6miOLQOVFMVw9y0o8iTtR3Vdmx6rrDarTy29yXXCOufnC3xhPrIwO9G
mwTFEEaP0dPDZF9wDuisgXfmIss/2oXxtmEaoGtsCihVfOQUrmt22vteDbWgZFK9gv2Owf4ezZIP
/Wh4mSFJT75uJmPKmBg6tXbBlXeQs35AWAXwu1+07RryB6ppItwvV4TGFKSx4kIOgT1y85Ym91HK
0H3rsgteNtAZQpoXrPy+BFwtbY4gFnyXG3xmUhi2a+cHt0RArgQ9b6UHDcQ3UnJYuLUZlU6E5k8r
m7LpzUHE+OPhs32jEYHMa3wI7/HhcdLw0gkpiqctZz4t3tkVLMie2cOYbKwDuCzUSEm9TqsXqT/z
Bb4aJXJ8kDHa1uKue64s9SQcidpMAWrqhCsiJPKVGlopV6HNeeA/nz4MoUTJZFvZLzcsCOT7ride
kpGvZZyDd25/6BBAg6yjF8VrC6zggKBO1nuyIddRiF8z/NDTPf+hpek1GJnahVZwxiLtbdinexjr
UCLMsaTUlyzSYom9NmLhDCFW4JJ47uTjoglqM6CJ7RnbKce8B5mCJAMuiiHED7Y4sN76nmlVlcjr
iP2kbt9abheX6yLcP7bA8Tst+nueoXN/g8CcfjGerEOfHXtVVH+ActpFVAha/tE3vkQAge817QyG
Ku+P+N7A6KjkKZu0lZ9yBK9NQp09ajycKbSTcWv5khwlB/x5T0vYN1sc7cn/5Suw9DD3UP08XfI9
dEatNa4Ypa/0cFOQWPRjkkDe/mN0GFyBpOSVNWw+T7FBDh4/HHqJIasJKkuBYUT1tyRn5PX8vk33
R2/3+048sD9lp0KQ7dVXxuWbpeZ30Q5aJflyPD3Wxj+ke7gpNgy9+IPkI9ljZ50BGImiah2NhP7I
C6SyW6NzEN9qy8ohd47uGYUv3e/Ko4ChMZg0yvO0sTp3isIUfeSmYdmteDtu+9Pgqht9IRhU4v5w
hjS3JRCYL17fcSI0UVg1z1BmqpR2Q+Izbv19u955QqV9HKWPsYFNyIh9B3FYR2vSx9bw9sOfBNRD
KFEv5pnrkvHKWoUw/79kxKij+ju3uw4WdyeccyXhv9auyedfuQqchJY3HjJiIHo0PCVMjTqmq/Sm
BjZYRJ0B2rs2X4LMp3+qpiMlrPKpbUHYu6l3r5u4Yo6vK7Jo0J83BbhsGEryNHh7daucZk5ANQZh
f3D81mzT0LHTwgRFrHMPx/G3MkHMVgFcWZ7WzV+RKdRkIH/4y+Rys0ueE/rLyXO7MKln7RisjUj0
xH01dVQowso0FlIgdAUFiNUL1Tm+SjRn78Dl11+HZQP2kiWF9v86lByauoRGeHklZsvKFs5fvpK2
xDAsCkP/Ml4Mcq/tf4yXv2C3ISLqSkMrCV1TIB5/1vrQ57B/dhL5rFGSsX3W9D6ly2kjBI41xJd+
wJdVgmY8L33Oxtse8ScBuliUrc9hJPaYhy1gsbgGXcHNxP3E+NItsZPqLZ9cp0YV8V6SzMnt0lkR
O4QE5gB5q4SjK/Ih7o2FINm+cgLJ566uScT/G9KjQ5PS7vxR2dfDJN1P0/SGML+dUAaEmIMVJTNC
ZNDT3ZV95fK0A+5PJGvAf/cGmDXacpHMMS/lxNJkE1Pj1MVq/gmbcpLrNVVJf+zGv897gFGv76mK
Dp21K+zUOVmErmDyGq1pNgUwh0w3kZw5tBVYo/8tFDOvMm+8JLsh6RJay1y7AUZYG5puWsNwIqO4
eDNhBJxQHv6bBAFqyDCpPK7FCazFGAV4Rg1VfxviDmw4KHbx2g9C0G6zaeEmEaxc0o0Kg1wYPE+I
/SQeGC1+LLXQG2DQ0+qgfkbVksEWGdMGZWQLisoIlCUGFNrIiHUYCJQLWW4IQHHQAN2Jqzr/Hvwr
ZJJOQ7WWatdQR49Ky++NdriC3A8jYyAhJaB/QBLVxDFXNK84tgioxyokKlhYDo/MHnpSrfA7FDzO
pu/OqxOTn5w23UjjZLapeaNAmHIQTuxNdRJXOoDRjo69JSPGCiy8rHCXVd/+n+qjLy0n+ztIX1p6
bU+bqtCyuf51FruM6cF24HZeNBpPs+UfvbtDpQzpF63r73xOUhqXtYp/CW+Hpo12HjxedfhE1EEG
+3m85HmFaRgy9FrXBB4gDhkNMmO/bBvtP4Jwpifk6IMwMOVPy279gE2IQdMk62DeO7JDO1YVzx7p
6e6bqcnZr5GbM156ze0qlDsQAJWz7GLN6BM5i3ga+/JYpvBT1BP9JzjgMuDWq1dtWkyWRe34uCkD
ukG+kmiB7cLpfvarob8dM5QEisa9771Feq3s3sg3qMzWlAsbAF6V7MUE5RoyXERIv8TTev2GiG2S
+zTeUy5jIfs3tdIsmGkrhxzeftzpLJgqqbdTk90JTUHpaR0SILiofxakYDh1IcX9AxmzQdjPHQB5
yViOqjOVm9/GdadW/26pbryJ2lzIARq2x/6zcXUV307AS4bd9TVxs4tdmgolPUZ+iEffbTSpBy2C
9Lf59asiw3oUn4u/I/98OS2gSYhIUYoY48fMRQJ9pwte6rvDP+1NkvFCGzHi/toIHYsbOP3Z0fyh
XR23kHAGsv/mwsu41fO6kmYA28lmXRc5SZmtWIzTJmmD7OEfnJ0RdZKnqbKDQyBVwDKJX/PABfCv
f46QF++9tb/pNjlWLHBhJY1VhwzrxtJfYgT//Hihax/qEcuW4jf59KLKU3GSBslnxH+kBYkioiz6
a8mfVRoaNfWd45vwG2WQvuyOKartURlghjEFXgahl8SXdD+b4vZBaH3kUYjN5bxwy1I4Vr+mT+F2
kUQU5MgUgTccMikqU6gXB6ZNeHE7R+5/d3HfkOU8mIZifFDTQGWLn1z29tPqmURPZwTMGwELbEpl
dZdv3MHHhzAUK3lGKLf7pnDUzom6EnVpCLOZ0QaW5modp5YgtAH4Qs8cig0Vk9gOZfGB3f4wPTvP
WrgwSUL6byxaNsBv8c3a+YWIfycTSxob07TOzCwri7Q1iEBa6HOGM7AFghz8reHNAjdBmYVFJZeU
JcF/n//kfXHgagYfICzi5Kjemnp1wt5Umi+ohu4y4Kp6iDplLXrCitu6i7EqJCmuVDTh3d6Cz4bE
a3MusQBjNt6XmgFdeanT2E8JVf1sJgtVni40zmUOGUfdjxXA6iLhJ8w0SdBubyjGPfFl1vOEOAPc
yoqliB/I/qy8CE6r3FRswg5oN1fxji2OfMGTjxFSVVl8MVX/vsdi61IcAm09mmcObgDpPM+z0dK+
CD2S00a3qLx/BTfKmaXXQLobvt0S4ShV++05epIQfNnSEyzIvldvSXX45G0oa5Vp/9nwCDn5E03n
ZamLqcbvm4mK7fydqZeQoiGm9D6HnLmRqNJuETieudndBpdNQ8RrYd3GRFWsZbQP0nVO2Dz5BkaN
LoKQbISeqicvIFDJMrG+BOfIQheax9mPTyGHqxFIJhPmSCm09vNwrHus5UN865Lq+9CjrxenWVoK
4W7m93d3ylz8Vh7bfhLYkIl9rbrI+gQd3EnmK3zVatfyS5ia8Z7ImHLVp3fnRpESsbLBCLAoRJ9f
3q/Tgz3Xoc6v7q4NNxS4tP2FQK8kq4t2DByZDoSmAHTeBmqm9lKK2uEq0mWeayTrkxQF6suwTZiM
mOOm3ytkejl2JL2gQrwiqCnevUSRy6xOlOR3KsFv1nf/0vFnjg4WVKz3v1qIY0X1aReTRuEd1jUx
Jl9fGHdC2BSC6nZ6jJyuBdb4RL9dNgIR+JS234LLHWGOQZwnetqdcejsJwFLl1I28VZHui0XsdFR
6/tl8nCo79ELW9fikQfR2opQwMsoo8qJ7i2O/mHGwwiss5gBiricpNTeTtQEUj/YlJipv8YbHdy8
L8yNAOAUPT7PruX2N/nIl9siY1hRUlEUtNfCMg7uqgRh6VQ91IuKPruO+Bo4DQlPbsIiVGYQ0uMF
or/Tmi4qHeE23Er0g/KJMVfDLaS6m1ia+igH+tJ0xfxnHgoiI6Vx9jk8AHPiJqUfA50+bm39PNeb
Zq5SjOhnWsCGWZKKE8jn5m6WLIfEjGXwjYenUqV92b8Dql6GiLK/b/NwcFU6o/dbnj+HKUYyf26M
71/xmtRqmjyJNY6O06/9IFaoX8Ja5dunuE/yMBob/OqobxkcsfrQLuj+x2b9PBqRXvWLd2TFhV0Z
yvf8pQTBKWqUFGqE6CNFOnvbopsVV2GgX0HbWZqwFrUO3YO/9oi4P5iO1VkCMsCnfpJAVuvC5Vmq
owUsKnVgfspmfQwCkAlD5KPd5Wg/P7iS9Je7EKMyX3Y5nJ7y+KMjOJa3u1DQzTYTjbwboQ9Ak3Th
Ie5SS+WFj3uZ+2ueVBeYnoyhSXdxVItLs3Srs9BZSqJzhd+UWCxJMPGy87MHev1bO0djWqoA4Vdu
U9b0s2DIc6ul8unrlRmH0Lkdh0zqlip24Fh5XDWvoVkM6l6Xk4Vm06SuBr0S57j9sjn6lVK0QLl8
3DinODCFTsWTCaD/qhu/+KtCCS+u6fD8YrPQWMXlPyaiUYbQSmgvvCcjyyf0nAjDLdIN9C+O9W8g
AtlNqYA+jmMTmZTgSLW4MGFJsdQjkTT5Y7RPC3Rjqe7AS/FECBnxnSDhxOqWMJZcnswvlU+vKUdA
u079xXdtn+SSvPkxf2//pCnmiaW4o4pkHPqucdHkebh5sjEIdkQtjG8z2Ti6gHgoqE0WwSeY1XDK
A6kr4KyYnyTZCz4rbHjjsEzesX4PHWTmDTzKcPahdlPP6Ai73kx7BWiH1o89lPqtNxMzxEQ7oTDr
HGo5fKUTKXeHfkk9TbkTSSfzEHIBaz3/IHqE0DnFAylfjyuH1D/+j85uzw9boD0dnyik087ba7E0
eXHNz0tX48DA4UWOj8NhHE5+Wytc8og5+5UBqDMaq6FMH/GREP5YvroHCPhjNP5zGxW68ePFTuYi
FyD813bDSmNidlG3jQuKMHSYAYaroYPIcvp9zWhGKOfaiiBGo5Xpmir7vRCZVMY5bHUAdaOSydTI
op5db90ojfArsIzPRqBGiWdXlF66WGd0f0lQTGt/6cV8miY/dFLK7OBdEVB/1U0Srg2WsbWFLZRa
f4lsiYLRZLIHELv7GzOKSLuKQ52oPWF/RtP5UitbZOU7iJU+R19yo8h6uMGou3855MLLsHzIJ+Zo
W9BFKbCwaH9ZGQjgIhc6Yt4Si4KPfE5OekZuNNyS0ejBATcjQ9GzL5RwFIeAQmkJTESvcZ3qSnvq
mVBHJrByYs7DgaL6nWpP98aUHUTWkBp6z3Vb7o+ieFIhXcyV4aEj56Zzf8AaWCiXO4vPtAFEWYSQ
l/lGPPtINs14Vl6Xg1AOaReNJp4phG9hRXg+pOs+vZcFu8XgFZ8ep3FmgsdxRDVuT3B/lccBW1E4
5EFCztq+4CxKM4nirGoxKjQTWNVLOCbu+ZjaJeboarkZ3KczgSZPaoJB1F1VPm8uvjKHVMETc0sM
R6KnL2yEYYJIx6q5OlGkkInZ1TNtR7UAQubCUdqS86RSrpmIPeqP19MnOwj9Eb6hOHGyk0YSGbHm
gh8RRdRl1WSA6kHZbRRGxZyag+JwUrWpvj2GTWD+FCYPl9LGbCgfVGREHPFREPEwpAgB4M/jg79B
Pmp0KwlHKxx8Xo0w2XhgYFuHYaTC+bN7tz1sbftyVAGxON14MVojECwO37sD8HYQamKHzRhwpvIj
DXaNZZEJHa3g4+cTzAXhiv4f1DYwYscu9v0HvTRC8dNV4ekTIhBm/R8KiYddx19f5FKl9dK7kL0I
obtVm8DVVWlKkMeQ7p4v0SLvw28WvdTEgmiQRm672JSOOzwSL+aPA6iM0DmMhpqKDRs+CRVeWdYQ
hahWN/857d1LZY5lBBq7QADBuqomUYvKUZUiyjaI2Q2RpBh105mWa2Stb6TgyM/r0AYZl135pj9x
THdhkZ9xHl51LgDbyqIl5UTOMKOCw+emkaFCBNncPRl7Fd6EvaP0ItxE4dVONn3zM51rRaRZgHlu
RRcyKGZ6qVxyRMMnvMwIn8mQ5hAdjhZajpCBXGVQZ4dkcTY3ZwPaVWdJIPrqa/uZuICZOvUni6IB
ZzxYM52V6SoLI6FFENcHilMFDNHpQoTUIrh8vXdQTEini4rGBSLQ/kPA+zONqh2xVilB2dUrM0uH
COCGONotLbB0i7MP0sLM69zXFNAU62O8d9pvFIZJLmuJ5eKdEep1phGjWpYUqYy3OxS6OrlGZqer
4u1RSMujeaJY8uWReYc/o5y5ZPuHCIGlyAfhZK3w+ACrpZvWN6zSmkoEojPicFYNlm2Ua0xCG5Al
cAQ9dKlxjkXkoECfatbsE7dC5D/F8RiXKgDpXxFOpyBPS7aVqDhS/CaftcTJL6HzpEZFdRogW+Uh
pHyf7ln5wo1JsVhapJ8UPdMTy4qhew6e9XkorfDN64gbD50Nth2CWLnvRyHPiL4mFQVjMdNBMvc8
A3Sea8MUawpBotvkePD3Trd8tmlM/lxFXBnZYrfzyYlX84CT8Auxe/rcuKwphrQxE5W4iV2rfo6s
3ZWvnQ9vs8M0tznpti8eWHCmd2ZDO39CBfCiZxwTk+byoG+OSwj5ypZ+P5VqNrPx0mmLy1aQuQAg
a4MgM6BYQUv4YijW5uaZ66i1WR1ccxkrW0g8dRjSFbermCO4cJsZNhGOhqKBBuOs6XI2E8pDkJNo
W3YajFf9vzLgnEwqA1ozG0ZrfmeNmfLz9+FzkImX8dQLpyLNoFhHCkDPzZImNxb02ZN/tL7IkDKr
mp2GyKe9PudsX/F1/zWx8ZWCn0QqyPubr8MWYC7uE1Uj/0+FpOa/XfxiCHwRpx9cUo21IweYoELh
n9sjB/jdLudkGuCqs2LSxMLGGqkJ3sYFO4uekpbT0KVMJAiUH3auUYqePkHt1EQm0kRck4RG83tB
et0+SRJsQ1A4YWKgsyEZD9C0uJ9DROA6SAf+a6rYjrbtNsuXUfjk386W9PgscfCzzrmPpNHSP9Qf
tP3kZVIrjnzhSK5iCLlvHIZ95sw/MiQ1aGJOyA2VkeXsfsFguIKBT2ko1Sn7CTsSwTruZnt9YdxR
y4lhzajL/5ylvBOcjuylla7JMqXgrZ43wrRO6PKsSEPFdhDL1pqYQEVC7xc/6YI2s80kA/NObdl/
dj7MLNnjeiUhLAcMKXw5YEVklm76lCbSdJytf8OtLD2wdRv1IbtL1mz1BZt7x5cGf298AJb0zqsv
wmI8LS85djJarW6XZdOP4H21kdCOsUE+VI+4yqFERFqeSULLeNE8Y18xejPpfJKipYwLeeB7+Ckp
WPV2OSH3/ePYKHEZ4Axp4MBYY/6Ld04NRxq0i6rNbbuz+nl+pzFNyH2++rFuL5FyFppt1x47rhI3
pIxA12lIx57Nx6F1UlbJeTspBZMVo0eOM2GqlHJwA1H6E5tlAlRBBK8jVxGIypX4jv90AYE/3hws
QszrdIP5I7mLmTAvoICHXcD9HxtOD2Tcf0FXFipZLQjOn194V1kUs1WkTuwCCmbLuZjhmhFc676Y
yqGJ90Tb40D8hGlpN2/tuUAsngEtBFDOI3AWT72eACAcfH1MMxbgHBaC+1eXlFFlQkfGEeIyi4pM
RjOLFfhkyHUEkZb1Xn1y3RX78s0TXd/wmCjrlQiTQbPL6fYE2/g2h1WiH1oaWKAI1Lxo/T4tSkkG
+R69em/NaB+Z5WPNMHaUQc+AvsmfQEjzDLthY+XGhsGJ1RiUBSuixoZ7tRrH0UHihcOyBnumihsZ
x55e0fySUSiu4h6hA6Yv9JUTAOmVBJpnjd+DN8ACdiD++ziVBXczmzPFC9Snz2k0BPIwR3jXr3TV
TwEWkX/TyEk1dmmu9YHciOFQ9Sp1fufEXJ5zk8f3m5/qKUk8sdfhoC8EaBUhAaBfj39a1+2R1Vdy
xZTRFllPtmyu5m7pp9eZTk4Q/4o3u24iQJfwYSTUVmUA9c4t/SEiCp/6MoxJlzyTbPO/INDEnMhT
dJ2PbjK2Qz7fBmevPPZ8AD31oYtmljFskohufHH8Mg5Zt/BTks2VhLY9AhSDtO3JNIAsOwxap3cs
ZMOZMh0RJjIJzCsiCJ7ePiY2jqbLJP5hBZiCSjm6yhb+w7lyKIULf6X3D4D2UCB4ALR6dOUJesr7
M7Yb57z5ZS1SdYotwRJMrN6l2KMLXcxqIVMpvjUZ7Lu4suQ8R0hEOMaLFSDnWuQq4AQ+8k+7+tbW
+JSFLxtKnqB1aGGfqp+FGCY4y7jlZhu8XKlsRV0TSFL01LMHDw4MbyqEBnQ3nPtSakVWeCpatJu8
MW7dMQvKNaViEEAmSdIe1F3R7T8cPiVwPVYuzXPT0+uuDouap8rZWIzUcpW4A1jJN3cvzrCLPl5D
n+6I3re4s64FKw15kqwsefCoVZ6yXkMLViDcxqPWT7+HePQ54GX9Nw/fI7Wi8pxjagDW4UVsCOTO
+FjcsbYP6eHI0cj4KXeKXAVXWac1ck0ZE6mubnTCA/Ni8RLbiu13FxbdimvtUa7+a8tCSvC8sYEB
QQFPzE+DIIUhqwwCCGHDpns2vCbWuPo099cyIFJ6hWoprf5OnZQv2NFwuPV3JB1UsNL1R2/4TQsx
lXR3jurYstus3rqFv8GvcBC7hkDYwzgXOJ8nuLK6J5CvARUky4E6WH80yiThXEWUuKwNLoTwkL29
0NTyx7NV0EnVEfaajk1ldbwla2+HWXegqIFkDBTpFP7mL9caF/lzvYPx86tLTYOQDaafnh4JA6wn
geI0LjUVkdO3CehK1bTmJtBY6uJO5KqEnZFB/gpiB0oT2rh+ul4iFgSbbM3lWQeX6ZPVZRTgL/0U
SyeQFPTheHfeffoTQBGcvvMzQ/9chRIbV221Zd7ygLgRDbaqLgoHd8cDkSPJz5hZ3H6bPNXsG5X0
YAvZ/hi0tQyIxn/2790FbYCd4qCba/eHgiE9jUYs8zimomrZiy8vHXr49hBAq2RdqCExPjiySMnG
zhfz2lxEiOhTeGeaZxgefyVMkDuW+q6uZxrq2TvDUxthAmUK47XQB0l40T/HSsiLLzKUZRMEPW8P
9BzItWr/j7bjZ6P0ywwjn5v9OAryF3anyEg5ZXPNW0tSpPKu4cli2qd0m6M7WbdOv/+05WXL+GOK
8SKtotpI5mkBaaJPHyop1ZgrfufJXBnFdSGaHIHODL6RdI7rdEGoW72DMqg3yUh3IpOQGU5Udg4e
tF4LtO36/QxiK+pj1tt5ZVMdqudXHPLhU5JAEaIftYFXgoEsIl3WJ3e2Kv7Aeaftf6PFD2h8F9KR
7HHmrJ7laL1i6Afw3OXYu5yDGx0SjuqxTShNmR5h3ta9RopbfXu3+1pqd99GjNsKWpYABcVRWRBN
/y/7YHjdXPPAeCxV3bJq6nfZy+/k+KdrE5MIl/RiKAMXUmKyah0O3E0A68LyKDU+OfIyK+YkNA==
`pragma protect end_protected
