`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
GtonvLyRIHa0BG5ascvXN09MZ3qOiFCm0qhQWasCekdFVRCizFoeirO1cOSD3S/L7XBtqzCllo4q
Q7pZwE0bdQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NcAWItlcyJiW5iNdkc1sQhABTpjXqZkOrg1X+Tcfgn7grREOKMnmze0hKfPSK2fx03p+1DXa9nI9
aDMO4y3pcvrSQRCRWXgMFS2qba1ARCCZEOEfr1i6f6+Nx8FGN5X5I1YnoGroW/YZxqunrLG+EqYi
XcxUyjBIkX9CxLSivhQ=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LPH3S1XGG8M+74c5vorJTX4Jd0Q7p5hXR2nHLPyVATbLKyNyCj3u2979H/5+r0KMFY+Eci03CiNr
huLATC3oqO+Ri3s+z9ShUHH0kb+eyBSFWWv4Vz/y3dKeMo7xd/qiF6cFD/jwZmVC699OpPLFZ+//
+v9QSba8dbzt+SXEN/jt0+eliBPMdqYocom4RnNiRzWVLRpczdP8jPK0iZ0dswvulkciexDQ2OOo
AH7xVOxZOGncQh6Vnj6rFermvVKMjP+f3wo5tFO3kt6qIlYJvlMl4+beZEF1FvA7E6pKL2F1zinI
FTyZEqwMwZWW/ux/d9gBr39V6BUQmOQXaUku1w==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XhsVvFI9R4kEmwKEMm1/ve3kzL6X2enhhJxnoXVsTfGBwYA297bpytmIip5AhwFQisRjBoqJ0K8l
8Pn3j20/SKo4hFrQQGF0dNNW6natF+zLk6mmfJ9vN5kjz0dnY6GDFbN+3VxaI7EfmTameGip8Srg
gxxI126PbwVBsgU+CTpGeuVit895aMS8BmBuDurrl1wtMGtV+dEhJIRJc0Aq1Wrns6Y56i0yfgPm
51nrGVg0WniIJHCwCd1amAGBP8K+XEMqgFg7Ax6FDLMI9fkEMpr36t/NLdEvEWInQ+uThyiFxWQr
JKb25unvEuv/D0FeWrozh8XdjpoKLAw1GPNMVg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
W3obImnatzWtWQxjvGXfWFuKaXr5FfPdOSZAbNOW8Mwmo4wQnwYiA7HkLDXfdrmslndHMaUxH/ah
zQFKiuR+SbrPT7aIULBLqqh72i8AksoYWph5t+HS6djOrRH3vsKtdR3ywmgroEjQ2QUcAo6U9K34
zqxoj8P9N8GP6+jAQYo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
p5NJqyb9TdyH8yE0AGM2W7x67vL0sjxs/jTTPTMrKPRWFxxZNuqsL6RAPf/W7gzVERxAO3iFqJD+
UoyFnOxci4budxkwr1k61TSgdoxD0V3HQjFvRukqTPnveyj/ep+eTC4LGfMpV/TPdXASgmKbIegz
1MyLz2/mIQLVdf6YMINHpls+EKIpYMQZpwK/hPkYr3E3OOOvzvQxNC9VDhaDMvYytD0fGysZMNYl
wnQ2rJfehLe6ywYzM95pSaORaRL+1Yx2J5fIpMdmGCqTlIRPg/vBGdEvfU7LTH681IczR8haG53W
YAR00ATaZUq26o3QwofFA/jZlZZYcN6rMAOtfQ==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OsRx87MiUvQMyOGPSETijoG08vE4+CeK9YRUiBEhaa6o5uSa2mSyUldHexlwxMR1rBWiQ6uyqUCt
nOrLjKhAiPGydi/JTIixYfKsNMv/tZTwiL+UoHRiZBVFKKOx3LAC8mgFXdUdYGwZnPhPVBIrRJxE
Rc1n40BeUgXQa/BvVgZFq1WN5zlUWx0e+VzL4EHCQl8ppq0b9oCO2dY5tSR8oDlWW/ZOlS5/u72T
OBDaxVQ+J7PWFUnUbY29E2dI2dNIjwjCjYqO+AssBOBH6HZcymhsJOjXSsS6xO1jpNeJMejZ9zqd
GqVBeDYMHSNvyuKhK1iLew/SAb/tdD8vIj8Gsg==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AYMh8vGmPAmkV/4T9vXCAbcwNUQ/U5Uw5Swerl5fs3AFaCZc0Qd8qyJ+58+zr5M2R7LYmJxqm46e
wTkAaUYx5X+VmZ+SG/c+BTOKZ03KypVWl/ISK1LXC/o7S+auCccud+8zMCxRUsKHuKYyIw/9r4Xo
hq9KP5hjv/dyE2FloIaus9WXSRmy3BsOrnOz34Y21Q3ThEHJzIUzPC9BzWKJqAiXhmZqFyQNpIPt
k/qfbsSvBqSTLaJSexAjyCb6KJ+cjdu04kb0KxNQHwNLCdnF8ejcSevf63EwGkmE+UzodGVDp+ZB
5rDYdmQGjq0EQCsB9QHiQJ9xNvYS9co+5Ki68Q==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ft/0b3HbGm8+/u8rq/UN1q9QtlQ7ydmhNvkUH1HFaaEw8IoZqW/LGV+djzXBf+a0L7Lslm4B8/ds
ZIPflSuox2viiVlo6Gu/oLKkTEg1tP9VJQ0SBlLuKdd+1Wtm5pN17pffr2TMr03eYDI2Wj8CqIF+
sz9vF9ralD5iy24MBrbk7D1MMaUjK1iYLEbGPul5XaMw+wCbhmYkQz1aq+m95hJ31EOKL5VFcBvw
0G1ICvealfGN8TBm1MOsgcXCDnEIfZlhrRoDLXx1+eTwJ9G46IioWqKUIgceTRCiJ0HPDdCrElbb
sSVKrR1ThH2yUQnQwI9fGdD6wpMKCSYrtlh7xw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3328)
`pragma protect data_block
ewowGykr0Xg9OiH+t3U9UlOPgMElQRW0LA6J5LYPrNqPLV0wA5QzeAl7lYortahRDwNCwnmRGJn3
d/GMWAW9/F3YuUgL37MHO+9Pa4ySSy4+zm59roD4KlFT8mq/d3msCWC4JSTC0FzADBnYtPgCXaRO
U0y91cmi7WPPjpe9CAp6HaIFzF913mnoxUS7vmm0t3nB6rp9vNGI9iAwSYKlQ+uFM+Ugjz7d0T09
48/5TNIVMwYDktCEArec6K/CqOlmxgaecDsgO3eIGRfmbql2uktOzDaZ9f8sY5/P2B3KcvUEkZoU
bYtrnMfFLvsEiBwlXBV2uCbFGd2Hf7rvCcmK4gfmsh9XfyDfJjNBoUDOIdggY5oj1lZjssYkCDkU
qo2Otq4KAyA/8GQlsR5ZTmn+s7dY0eFjzGWYUw7t+f9vM4DKkg63LthH8byZ4FPNGiuZd+UY+upQ
ceffWAEWgVshLZlHVpqfFZvCQhevUFKZmbKbXW9Q7fr/K8zqAYULPrjh3x6jZCrDDKHZbhG+5tVK
XDTtbu/ad52mCXXavBAO22CrtDmMdgWqXg4ZWVV7Y/hTcc+y43UFRmujEtFR92BMDHDxLAYbdg4N
ROqoi4jyaPBTrwcDr+BUDTulhUKLlPrxpNynTlxOxr2BgmooRdKD6NyM6F0ja9xJb5Lf9S4Awsad
3KVEqj3tWBc+DbfvmUsBQQh6DtXNljFi/8GkYeeHzKewmYDanG5pyOiVUeekHZlw5Rkj6psM/rEo
OChP1w8oWxOPN6kpdRctFK2RiA44BxpqHEQFomaYhMa8xiFDJ7K/6RFZafG77OoffpLpS5dF8/Tu
K+Dw0JkT/6lNyWKLAaszM4cA+eQfVsBPZdmlu3Vk9onREu7GB63OBm+cFiwvCegHHEgvbf0Qn9YP
ojK1VohnyeWbvJIqZH/b9CLAxQePkwtqTibz90z7LDTc26a5cibOGhwvnkAux4ewVIn39pFHloTY
qaG7+9hBxgs32u+/d74+x61McL88Pg8APvkEAWyNhZMgjXTijwz0fHeBn1xxHGJzAZyZ8Ek25caI
SbFlZ7MMYdQZP/D9aLsIcFHAyaYvCkjDFml3y/QrpGtTT7nqsfdRZwzrTDayPebhOTcT+v80AiiG
wLyDVLTzSjHfntgQzKMfszKv9o/9M6K5lHJdCCBjtZiohPiFdKydAo8IkUz7T/OTikRjUkLlFi2B
krexmaz5es1FbbijP30TbhWkboLIBcAIAGpIu06WNFhiECQQNQ4e/s8a7ZyD7IjiMrvwj04YQ7/9
sfD+BFmsTeaD6fc7JaV46/FNo1n9CJKmhNQ0+XzW7+mjfnR3oXWwR6uI7v3OBMmGsi/Mh2pBu237
IYgRu70teEuGx8etmgx8yiwoxgKRCg5GbYGF0IGycRumiCGJZiKog8ozNC9akk0CpowEK5KdKIY6
XR5Hb2gj8W2SAjwyUsx63cCCazCDKKt1z7MBGwrd0Phr+YzjMKa6b0nqt189gT/CQPDDrjUrCfHk
GCjhwOZljpxmkSeX2GYj7Ty34/0XQU9gi1tpT3oRuew5W+rIRe7sYI+SqYJVL3G2vlWwwneLDNkP
ks3kyppxbrFGB/tSg5WIwdW98eV9oJwzNLX2r1aUSHhLveniCHqHbHy/J/hcw2zR4q0P9vc8/zbe
qqXSG65hZAJjNGpOvudzbhntM8ckhYPKP9NKA852esrp9ESiZJELlBM+nTz7TSW+6qtffT8hmTuc
/SJZ6Mq5myO8YZK3JLky/26xqeu6V1tO30KbSgvxCLIerqIbBT3PuBpRxmkrFrpYI9eM0A7D8TCM
XZkNi7hl/QIDodasrpNyUagh8ecZR/0H3lzihFDEOQ0jgqCJ+re0z3a3CW1jQoPagT9oYPAyUZi7
Q23xglDbtbeCfcnw2m25ftoGlfp8E+vGKWEvWzJzO2DMs7Gjks4YjFixjqNxYxUfQL/qb+3iy9Fk
FeX/cwSEDmgbigoK82TvM89akFSsfXwNVsihTKU8/trjz0Lv7TZy30rCSPsa8L0Nfy7/KLCFPP32
NfW1gs6xLJUIsrfCCmtXj1+26OLMSobvj6h2qB+j/nzQc8ExW4mzJHX4PLj4ivB9K6zpfNM4cVqO
I4F65Tw09f3ZTb4sRfBiHz61H1b9DwZ06jKNt8JmgD8FY8eavliPmGBBZYQsu8GbF5d4arEdn8Uj
nGXciCyeF9Gtkk01YFZeEtWJdaCPtLsjliOYtJkW5ajV7uJK+15jSP7zWEjihjyeRL9meSVLeVJy
aUSTJKK1X+mh2bg9IePE+xJIS/IBQ+mhnXdAvouvLgbS1Ai7y1AGH/WK7Eohk+oJnss2mR4i7r5e
TuttvccPnNKmZoM3t52fOX6XTwT8Qj5wdpfPYu486vtFEZj+laaNkUwTRKI8LhAAxIjUitVrGgvM
ZYoWjr1JX7oSPFb8/vjMXkUUZEWKiUL9qShCo3Ll9FSWfJAWk/mBE9LyIQYvSgqNM6nSMn4zUruG
jI4ASsuVI5Xt94y1HOBl7pUQzJyXYS6NPTb7QKPrrL3B5QxoZy5hOWlMb8NihOsX/RoWM0h0nXOp
n+JmZgI6mjnYkQA9rJU7T8Sj+tj+VQTaE4C/5mn6Ykum8lyqzte5awyFuVooBdX0jqTpe9fuv6k5
S4HZZlyqq1Xlcs+LZrh197QcolkkTgjrY2cYbCACUeDIkPmY0JEa7cyvXk0rRCYWzsp0W9GiV6mO
pZbv72KfLMSuMjWcUp6Zcs6VUGAa+hczqBT6Qc36ohYvqgAtWxRQDCmAn2xSmCQIzwSmgmLEI1Nh
EQTSWUrd1jvoe9IjcX49yOV+IsNKGqDBj7tNOrRnBliD9ELOlTVQXYltB4+TwN4fblB5YmaXWWkg
n08teLhTKeIm0YCTUGl8np91/lYu81ycx2trg60DopGoyXcD/tt+oJvDWXNUN/KucSH/Sn+pUZDa
ekKgiNIkZ23mprt1SuC97gbZxqh3UOTYWeBb+fTe4qr+ktFAnVn3mwUgwfgCEYRIVBAGv9YouoK8
VhnC0DRrKD1/InLOJf2uG966kxoqHPGZur/ldrt9EdmSW09k5eqm6Hkg8cdXzZZMHeg9udV4M9LJ
pplAEJ6IqFpXTIz8RbZRqZ1FyBtJbEad3L54XIsPcEmkq6Xbj+LwLtRF9xl7BBFVtzfXDpNK+dbj
OXbEDzghEwG8/m2p46o20D0mQGjkIGzyKl0r+UhlG1U7k8RdCGzRWD3W6/9kvQLkR/56zoeQIWsg
7i/3WtvHRyfJIU1+2zsjwW1AFAnjAxiP2n3OJc+7JeqG92acwuvViM+00h04Ikd0nBG5xBrLTL0M
EvyOwQW15NsXsWRd6EsDsYHInMu2Um7V9HzKQiP1ElJCju5Fpr+N8bT2NWmdrXDkEVnJ9V4hqXFm
mp+67PZ0qRnv+WqZdf5y1G/tHCnVIWbO65X38fM1wG6yXjNL7eM6OFRbAqdp4GXpEwReXQUZqLRG
cQAqdZkNRcp+eIy+AXM/7Xa025bitaesfD/MSAZ/Dqfl8jIfLAUlwCtW/hP2akDSzA2k6G0Vpg+3
F4dEBsKoPdtjdcfKw5B8inGXLDDGkT3xbDmHDcwGz0cJsq9Vigp3ZbpaJAlCkpv1BYBHTDc15yZo
Fljcn+pdmFb1V4Dsj3dthHtDcJId1BuwhN92TTrh5AKrb+WH+NRhWqbw80waUOl36Z8D5k7D0KOy
rH9ZV/ssz+/9aPOCeG8hrpHn7R8/RMm3I277l1nBf+Nc+AQeo4L7AY9FbptHlJGRt9vkrWm8qCnz
ltgVGKnJbCbn/0Un3zh6W7b1w/TzkL2FzD0yomo0hHs4LwNP5/TmQLDB/7t/aOZrSg7MyZpGj00Z
LyfB+OeOPhkrOXDhc4esoOBGfdqRcVzYbCocMTrtduREDK2PEUMaoDD5ACmpaMlAKTgFhKCF/2mN
XyTz3GT1tCTKXG6jLQFmol/J2MFaMfjc8seFTujufTOQJnO6uKNdMoF/qJy18i3FWxksjhIc31Mm
fUctcN/zyHZt+skBi61wGLkk/9z8eIBmtff4+lAypwKQkxvVQzZUBYCjoCn2AT8mLCSUeNVZPq17
tvwnplh40ErBj23cuY6TKyk6v7pSmJSMEFnaNZBHueh7ZH2dlvMuEFJESt9ESqIbC5I9nK+oNd9Q
UDnAdrd68roPFQGfzowbbufm1uRwuaog/AZbJZapGEg3x5QwY0XWx4M0bjXpcZATbyP17d/FZb9I
320ntyJbNEOV74dZceXJX2Tz5V0quviCVy8FvGuhItRoo4MPcoUTGqTtTm1hushXtoNYDuNPl1iw
8vF36jg7e7Etwi46o0JMrA4ML6Kw/MNazs+3fa/IvQB7/XIwSG5+h8W5bndeHaGiCCDz8g45Ap7C
Vc30BlO0oQLWeIky/O6xXcSW67TSIQ==
`pragma protect end_protected
